module test_circuit (
	input in0,
	input in1,
	input in2,
	input in3,
	input in4,
	input in5,
	input in6,
	input in7,
	input in8,
	input in9,
	input in10,
	input in11,
	input in12,
	input in13,
	input in14,
	input in15,
	input in16,
	input in17,
	input in18,
	input in19,
	input in20,
	input in21,
	input in22,
	input in23,
	input in24,
	input in25,
	input clk,
	input rst,
	output out0,
	output out1,
	output out2,
	output out3,
	output out4,
	output out5,
	output out6,
	output out7,
	output out8,
	output out9,
	output out10,
	output out11,
	output out12,
	output out13,
	output out14,
	output out15,
	output out16,
	output out17,
	output out18,
	output out19,
	output out20,
	output out21,
	output out22,
	output out23,
	output out24,
	output out25
);


wire net11589;
wire net11583;
wire net11582;
wire net11579;
wire net11578;
wire net11572;
wire net11571;
wire net11570;
wire net11569;
wire net11566;
wire net11565;
wire net11560;
wire net11559;
wire net11557;
wire net11556;
wire net11554;
wire net11553;
wire net11552;
wire net11550;
wire net11549;
wire net11548;
wire net11545;
wire net11544;
wire net11541;
wire net11537;
wire net11536;
wire net11534;
wire net11533;
wire net11530;
wire net11528;
wire net11527;
wire net11523;
wire net11522;
wire net11521;
wire net11520;
wire net11518;
wire net11513;
wire net11512;
wire net11510;
wire net11505;
wire net11504;
wire net11503;
wire net11502;
wire net11501;
wire net11500;
wire net11499;
wire net11498;
wire net11495;
wire net11494;
wire net11491;
wire net11488;
wire net11484;
wire net11477;
wire net11476;
wire net11475;
wire net11474;
wire net11473;
wire net11472;
wire out0;
wire net11468;
wire net11467;
wire net11466;
wire net11464;
wire net11463;
wire net11460;
wire net11459;
wire net11458;
wire net11457;
wire net11456;
wire net11455;
wire net11454;
wire net11451;
wire net11445;
wire net11444;
wire net11443;
wire net11441;
wire net11440;
wire net11438;
wire net11437;
wire net11434;
wire net11433;
wire net11432;
wire net11429;
wire net11428;
wire net11427;
wire net11425;
wire net11422;
wire net11420;
wire net11418;
wire net11417;
wire net11415;
wire net11413;
wire net11411;
wire net11408;
wire net11406;
wire net11403;
wire net11401;
wire net11399;
wire net11398;
wire net11395;
wire net11393;
wire net11392;
wire net11391;
wire net11390;
wire net11376;
wire net11375;
wire net11373;
wire net11378;
wire net11368;
wire net11367;
wire net11363;
wire net11359;
wire net11358;
wire net11356;
wire net11355;
wire net11353;
wire net11348;
wire net11347;
wire net11343;
wire net11342;
wire net11340;
wire net11338;
wire net11335;
wire net11328;
wire out7;
wire net11326;
wire net11325;
wire net11321;
wire out10;
wire net11319;
wire net11318;
wire net11317;
wire net11315;
wire net11314;
wire net11312;
wire net11310;
wire net11309;
wire net11308;
wire net11307;
wire net11306;
wire net11302;
wire net11300;
wire net11299;
wire net11295;
wire net11294;
wire net11293;
wire net11292;
wire net11291;
wire net11285;
wire net11377;
wire net11284;
wire net11282;
wire net11281;
wire net11277;
wire net11270;
wire net11267;
wire net11266;
wire net11265;
wire net11333;
wire net11264;
wire net11263;
wire out2;
wire net11260;
wire net11259;
wire net11257;
wire net11254;
wire net11252;
wire net11251;
wire net11286;
wire net11250;
wire net11249;
wire net11248;
wire net11247;
wire net11245;
wire net11241;
wire net11239;
wire net11238;
wire net11237;
wire net11236;
wire net11235;
wire net11234;
wire net11233;
wire net11231;
wire net11230;
wire net11228;
wire net11227;
wire net11221;
wire net11220;
wire net11216;
wire net11215;
wire net11346;
wire net11212;
wire net11462;
wire net11210;
wire net11209;
wire net11208;
wire net11206;
wire net11205;
wire net11204;
wire net11203;
wire net11202;
wire net11201;
wire net11198;
wire net11197;
wire net11195;
wire net11194;
wire net11379;
wire net11192;
wire net11191;
wire net11190;
wire net11188;
wire net11186;
wire net11185;
wire net11177;
wire net11174;
wire net11170;
wire net11168;
wire net11165;
wire net11163;
wire net11161;
wire net11160;
wire net11159;
wire net11158;
wire net11157;
wire net11156;
wire net11151;
wire net11150;
wire net11148;
wire net11144;
wire net11142;
wire net11137;
wire out5;
wire net11133;
wire net11132;
wire net11127;
wire net11126;
wire net11452;
wire net11124;
wire net11123;
wire net11120;
wire net11116;
wire net11115;
wire net11112;
wire net11108;
wire net11107;
wire net11106;
wire net11102;
wire net11100;
wire net11099;
wire net11091;
wire net11090;
wire net11088;
wire net11086;
wire net11083;
wire net11082;
wire net11080;
wire net11078;
wire net11077;
wire net11073;
wire net11072;
wire net11069;
wire net11067;
wire net11065;
wire net11064;
wire net11063;
wire net11059;
wire net11058;
wire net11057;
wire net11056;
wire net11555;
wire net11054;
wire net11062;
wire net11051;
wire net11515;
wire net11049;
wire net11048;
wire net11540;
wire net11046;
wire net11044;
wire net11042;
wire net11041;
wire net11040;
wire net11039;
wire net11036;
wire net11519;
wire net11035;
wire net11034;
wire net11027;
wire net11026;
wire net11025;
wire net11023;
wire net11255;
wire net11021;
wire net11394;
wire net11016;
wire net11015;
wire net11010;
wire net11008;
wire net11007;
wire net11003;
wire net11189;
wire net11001;
wire net10997;
wire net10996;
wire net10992;
wire net10988;
wire net10981;
wire net10980;
wire net10979;
wire net10976;
wire net10968;
wire net10967;
wire net10965;
wire net10962;
wire net10961;
wire net10959;
wire net10957;
wire net10955;
wire net10954;
wire net10953;
wire net10945;
wire net10944;
wire net10943;
wire net10942;
wire net10938;
wire net10937;
wire net10936;
wire net10935;
wire net10934;
wire net10933;
wire net10932;
wire net10930;
wire net10928;
wire net10927;
wire net10924;
wire net10922;
wire net10921;
wire net10913;
wire net10912;
wire net10910;
wire net10908;
wire net10906;
wire net10905;
wire net10903;
wire net10902;
wire net10900;
wire net10899;
wire net10898;
wire net10896;
wire net10894;
wire net10893;
wire net10889;
wire net10887;
wire net10886;
wire net10885;
wire net10883;
wire net10874;
wire net10873;
wire net10871;
wire net10869;
wire net10866;
wire net10865;
wire net10864;
wire net10862;
wire net10861;
wire net10859;
wire net10858;
wire net10857;
wire net10855;
wire net10850;
wire net10848;
wire net10847;
wire net10843;
wire net10842;
wire net10841;
wire net10840;
wire net10839;
wire net11588;
wire net10836;
wire net10835;
wire net10831;
wire net10830;
wire net10828;
wire net10827;
wire net10825;
wire net10824;
wire net10823;
wire net10821;
wire net10837;
wire net10820;
wire net10818;
wire net10817;
wire net10816;
wire net10815;
wire net10814;
wire net10812;
wire net10811;
wire net10808;
wire net10806;
wire net10804;
wire net10802;
wire net10801;
wire net10800;
wire net10798;
wire net10797;
wire net10796;
wire net10795;
wire net10793;
wire net10791;
wire net11274;
wire net10789;
wire net10787;
wire net10786;
wire net10785;
wire net10782;
wire net10780;
wire net10779;
wire net10771;
wire net10767;
wire net10764;
wire net10762;
wire net10759;
wire net10758;
wire net10757;
wire net10755;
wire net10750;
wire net10749;
wire net10748;
wire net10747;
wire net10746;
wire net10745;
wire net10743;
wire net10742;
wire net10735;
wire net10734;
wire net10733;
wire net10730;
wire net10729;
wire net10727;
wire net10725;
wire net10724;
wire net11508;
wire net10719;
wire net10718;
wire net10717;
wire net10715;
wire net10711;
wire net10710;
wire net10709;
wire net10705;
wire net10704;
wire net10703;
wire net10700;
wire net10699;
wire net10693;
wire net10692;
wire net10691;
wire net10690;
wire net10689;
wire net10687;
wire net10685;
wire net10683;
wire net10681;
wire net10679;
wire net10677;
wire net10675;
wire net11339;
wire net10673;
wire net10672;
wire net10670;
wire net10669;
wire net10667;
wire net10666;
wire net10665;
wire net10664;
wire net10662;
wire net10658;
wire net10656;
wire net10652;
wire net10650;
wire net10648;
wire net10647;
wire net10646;
wire net10645;
wire net10640;
wire net10638;
wire net11581;
wire net10637;
wire net10634;
wire net10631;
wire net10625;
wire net11416;
wire net10623;
wire net10622;
wire net10621;
wire net10620;
wire net10619;
wire net10613;
wire net10610;
wire net10609;
wire net10607;
wire net10604;
wire net10602;
wire net10601;
wire net10600;
wire net10597;
wire net10595;
wire net10594;
wire net10592;
wire net10591;
wire net10585;
wire net10583;
wire net10580;
wire net10579;
wire net10578;
wire net10576;
wire net10575;
wire net10574;
wire net10572;
wire net10571;
wire net10567;
wire net10565;
wire net10564;
wire net10563;
wire net11404;
wire net10736;
wire net10561;
wire net10559;
wire net10558;
wire net10553;
wire net11152;
wire net10552;
wire net10551;
wire net10549;
wire net10548;
wire net10546;
wire net10545;
wire net10544;
wire net10538;
wire net10535;
wire net10533;
wire net10532;
wire net10526;
wire net10524;
wire net10523;
wire net10522;
wire net10520;
wire net10519;
wire net10518;
wire net10517;
wire net10515;
wire net10511;
wire net10510;
wire net10509;
wire net10503;
wire net10498;
wire net10497;
wire net10494;
wire net10493;
wire net10492;
wire net10490;
wire net10487;
wire net10485;
wire net10482;
wire net10778;
wire net10479;
wire net10475;
wire net10474;
wire net10473;
wire net10472;
wire net10505;
wire net10469;
wire net10468;
wire net10461;
wire net10456;
wire net10455;
wire net10453;
wire net10451;
wire net10448;
wire net10446;
wire net10445;
wire net10440;
wire net10439;
wire net10438;
wire net10436;
wire net10435;
wire net10433;
wire net10431;
wire net10430;
wire net10428;
wire net10425;
wire net10424;
wire net10423;
wire net10422;
wire net10419;
wire net10416;
wire net10414;
wire net10413;
wire net10412;
wire net10411;
wire net10409;
wire net10408;
wire net10404;
wire net10403;
wire net10401;
wire net10400;
wire net10398;
wire net10395;
wire net10394;
wire net10385;
wire net10384;
wire net10382;
wire net10381;
wire net10379;
wire net10378;
wire net10377;
wire net10376;
wire net10375;
wire net10969;
wire net10368;
wire net10367;
wire net10364;
wire net10363;
wire net10358;
wire net10353;
wire net10348;
wire net10343;
wire net10341;
wire net10340;
wire net10339;
wire net10911;
wire net10335;
wire net10334;
wire net10333;
wire net10332;
wire net10330;
wire net10329;
wire net10328;
wire net10326;
wire net10323;
wire net10322;
wire net10321;
wire net10320;
wire net10318;
wire net11446;
wire net10317;
wire net10311;
wire net10310;
wire net10307;
wire net10306;
wire net10305;
wire net10303;
wire net10301;
wire net10300;
wire net10299;
wire net10297;
wire net11386;
wire net10295;
wire net10293;
wire net10292;
wire net10291;
wire net10290;
wire net10288;
wire net10286;
wire net10285;
wire net10283;
wire net11172;
wire net10280;
wire net10277;
wire net10276;
wire net10275;
wire net10274;
wire net10272;
wire net10271;
wire net10269;
wire net10268;
wire net10267;
wire net10266;
wire net10265;
wire net10260;
wire net10259;
wire net10257;
wire net11061;
wire net10256;
wire net10255;
wire net10253;
wire net10252;
wire net10249;
wire net11131;
wire net10248;
wire net10244;
wire net10242;
wire net10240;
wire net10239;
wire net10287;
wire net10238;
wire net10236;
wire net10235;
wire net10234;
wire net10232;
wire net10231;
wire net10229;
wire net10226;
wire net10225;
wire net10224;
wire net10222;
wire net10221;
wire net10219;
wire net10218;
wire net10216;
wire net10215;
wire net10214;
wire net10211;
wire net10210;
wire net10209;
wire net10204;
wire net10202;
wire net11374;
wire net10201;
wire net10193;
wire net10190;
wire net10186;
wire net10185;
wire net10184;
wire net10183;
wire net10182;
wire net10181;
wire net10180;
wire net10179;
wire net10175;
wire net10174;
wire net10173;
wire net10169;
wire net10168;
wire net10167;
wire net10784;
wire net10164;
wire net10160;
wire net10155;
wire net10154;
wire net10152;
wire net10151;
wire net10149;
wire net10146;
wire net10145;
wire net10228;
wire net10144;
wire net10141;
wire net10138;
wire net10136;
wire net10135;
wire net10132;
wire net10131;
wire net10129;
wire net10127;
wire net10126;
wire net10125;
wire net10124;
wire net10118;
wire net10117;
wire net10116;
wire net10114;
wire net10109;
wire net10108;
wire net10107;
wire net10105;
wire net10104;
wire net10102;
wire net10099;
wire net10098;
wire net10096;
wire net10095;
wire net10092;
wire net10091;
wire net10089;
wire net10088;
wire net10582;
wire net10087;
wire net10086;
wire net10085;
wire net10082;
wire net10080;
wire net10075;
wire net10073;
wire net10324;
wire net10072;
wire net10071;
wire net10070;
wire net10067;
wire net10066;
wire net10064;
wire net10061;
wire net10053;
wire net10051;
wire net10048;
wire net10047;
wire net10046;
wire net10044;
wire net10043;
wire net10042;
wire net10041;
wire net10039;
wire net10033;
wire net10031;
wire net10030;
wire net10028;
wire net10027;
wire net10024;
wire net10022;
wire net10020;
wire net10017;
wire net10016;
wire net10015;
wire net10011;
wire net10009;
wire net10153;
wire net10008;
wire net10005;
wire net10001;
wire net10000;
wire net9997;
wire net9992;
wire net9991;
wire net9988;
wire net9987;
wire net9985;
wire net9983;
wire net9982;
wire net9980;
wire net9979;
wire net9978;
wire net9976;
wire net9975;
wire net9974;
wire net9973;
wire net9970;
wire net9968;
wire net10465;
wire net9966;
wire net9961;
wire net9960;
wire net9959;
wire net9958;
wire net9957;
wire net9953;
wire net10566;
wire net9951;
wire net11287;
wire net9948;
wire net11146;
wire net9947;
wire net10845;
wire net9938;
wire net9937;
wire net9935;
wire net9934;
wire net9931;
wire net9927;
wire net9925;
wire net9924;
wire net9923;
wire net9922;
wire net9918;
wire net9917;
wire net9916;
wire net9912;
wire net9911;
wire net9995;
wire net9909;
wire net9908;
wire net10270;
wire net9907;
wire net9906;
wire net9905;
wire net9901;
wire net9900;
wire net9899;
wire net9898;
wire net9896;
wire net10464;
wire net9894;
wire net9893;
wire net9891;
wire net9887;
wire net9884;
wire net9883;
wire net9881;
wire net9879;
wire net9878;
wire net11141;
wire net9877;
wire net9876;
wire net9871;
wire net9870;
wire net10337;
wire net9869;
wire net9868;
wire net9865;
wire net9863;
wire net9862;
wire net11478;
wire net10060;
wire net9861;
wire net9860;
wire net9859;
wire net9858;
wire net9857;
wire net10246;
wire net9856;
wire net9855;
wire net9852;
wire net9850;
wire net11585;
wire net9847;
wire net9845;
wire net9843;
wire net10189;
wire net9932;
wire net9841;
wire net9839;
wire net9836;
wire net9833;
wire net9831;
wire net10489;
wire net9830;
wire net9826;
wire net9825;
wire net9823;
wire net9822;
wire net9821;
wire net9820;
wire net9816;
wire net9812;
wire net9809;
wire net9807;
wire net9805;
wire net10313;
wire net9803;
wire net10856;
wire net9802;
wire net9801;
wire net9798;
wire net9797;
wire net9796;
wire net9795;
wire net9791;
wire net9790;
wire net9789;
wire net10296;
wire net9788;
wire net9786;
wire net9785;
wire net9783;
wire net9781;
wire net9780;
wire net9778;
wire net9774;
wire net9773;
wire net9772;
wire net9769;
wire net9768;
wire net9766;
wire net10629;
wire net9765;
wire net9764;
wire net9761;
wire net9760;
wire net9759;
wire net9758;
wire net9757;
wire net9756;
wire net9755;
wire net9751;
wire net9750;
wire net9749;
wire net9748;
wire net9747;
wire net9746;
wire net9743;
wire net11176;
wire net9742;
wire net9741;
wire net9739;
wire net9738;
wire net9737;
wire net9735;
wire net9777;
wire net9734;
wire net9732;
wire net9731;
wire net9729;
wire net9727;
wire net9726;
wire net9724;
wire net11298;
wire net9723;
wire net9721;
wire net9720;
wire net9715;
wire net9711;
wire net9709;
wire net9708;
wire net9704;
wire net9703;
wire net9700;
wire net9699;
wire net9696;
wire net9695;
wire net9694;
wire net9693;
wire net9692;
wire net9691;
wire net9690;
wire net9689;
wire net9688;
wire net9685;
wire net9683;
wire net9682;
wire net9680;
wire net9678;
wire net9677;
wire net9675;
wire net9673;
wire net9672;
wire net9671;
wire net10369;
wire net9668;
wire net11580;
wire net9667;
wire net9665;
wire net10187;
wire net9663;
wire net9661;
wire net9660;
wire net9659;
wire net9657;
wire net9653;
wire net9651;
wire net9679;
wire net9650;
wire net9649;
wire net9648;
wire net9647;
wire net9645;
wire net9641;
wire net9640;
wire net9638;
wire net10282;
wire net9634;
wire net9631;
wire net9629;
wire net9628;
wire net9625;
wire net9623;
wire net9622;
wire net9621;
wire net9753;
wire net9618;
wire net10018;
wire net9617;
wire net9616;
wire net9613;
wire net9612;
wire net9610;
wire net9607;
wire net9606;
wire net9604;
wire net10162;
wire net9603;
wire net9602;
wire net9601;
wire net9600;
wire net9598;
wire net9597;
wire net9596;
wire net9594;
wire net9592;
wire net9591;
wire net9589;
wire net9588;
wire net9587;
wire net9585;
wire net10651;
wire net9583;
wire net9581;
wire net11011;
wire net10279;
wire net9580;
wire net9579;
wire net9578;
wire net9576;
wire net9575;
wire net9574;
wire net10142;
wire net9573;
wire net9571;
wire net9570;
wire net9568;
wire net9565;
wire net9561;
wire net9555;
wire net9548;
wire net9547;
wire net9545;
wire net9544;
wire net9538;
wire net9537;
wire net9535;
wire net9534;
wire net9533;
wire net9529;
wire net9528;
wire net9525;
wire net9524;
wire net9519;
wire net9518;
wire net9516;
wire net9515;
wire net9514;
wire net9513;
wire net9512;
wire net9511;
wire net9508;
wire net9507;
wire net10918;
wire net9506;
wire net10999;
wire net9505;
wire net9504;
wire net9503;
wire net9502;
wire net9500;
wire net9499;
wire net9496;
wire net9492;
wire net9484;
wire net10365;
wire net9483;
wire net9479;
wire net9474;
wire net9473;
wire net9470;
wire net9469;
wire net9467;
wire net9464;
wire net9462;
wire net10254;
wire net9459;
wire net9457;
wire net9455;
wire net11125;
wire net9454;
wire net9452;
wire net9449;
wire net10829;
wire net9448;
wire net11187;
wire net9444;
wire net9443;
wire net9439;
wire net9438;
wire net9437;
wire net9436;
wire net9434;
wire net10853;
wire net9432;
wire net9431;
wire net9430;
wire net9429;
wire net9427;
wire net9424;
wire net9423;
wire net9422;
wire net9421;
wire net9419;
wire net9418;
wire net9416;
wire net9415;
wire net9412;
wire net9411;
wire net9632;
wire net9407;
wire net9406;
wire net9405;
wire net9404;
wire net9399;
wire net9398;
wire net9394;
wire net10587;
wire net9393;
wire net9392;
wire net9390;
wire net9389;
wire net9387;
wire net9386;
wire net9385;
wire net11311;
wire net9384;
wire net9383;
wire net9381;
wire net9378;
wire net9377;
wire net9376;
wire net9375;
wire net9373;
wire net9369;
wire net9364;
wire net9363;
wire net9362;
wire net9361;
wire net9360;
wire net9358;
wire net9357;
wire net11279;
wire net9356;
wire net9352;
wire net9351;
wire net9350;
wire net10396;
wire net9349;
wire net10611;
wire net9347;
wire net9346;
wire net9344;
wire net9343;
wire net9342;
wire net9341;
wire net9338;
wire net9337;
wire net9336;
wire net9333;
wire net9332;
wire net9331;
wire net9330;
wire net9326;
wire net9325;
wire net9324;
wire net9323;
wire net9320;
wire net9316;
wire net10161;
wire net9315;
wire net9314;
wire net9313;
wire net9311;
wire net10712;
wire net9310;
wire net9309;
wire net9306;
wire net9305;
wire net9304;
wire net10525;
wire net9303;
wire net10094;
wire net9300;
wire net9299;
wire net9298;
wire net9294;
wire net9293;
wire net10663;
wire net9291;
wire net9290;
wire net9295;
wire net9289;
wire net9288;
wire net9283;
wire net9282;
wire net9281;
wire net9280;
wire net9278;
wire net9276;
wire net10956;
wire net9275;
wire net9269;
wire net9268;
wire net9266;
wire net9265;
wire net9263;
wire net9261;
wire net9256;
wire net9253;
wire net9252;
wire net9251;
wire net9250;
wire net9248;
wire net9244;
wire net9240;
wire net9239;
wire net9237;
wire net9236;
wire net9234;
wire net9231;
wire net9228;
wire net9227;
wire net9226;
wire net9339;
wire net9224;
wire net9222;
wire net9221;
wire net9220;
wire net9215;
wire net9213;
wire net9212;
wire net9211;
wire net9210;
wire net9209;
wire net9208;
wire net9207;
wire net9205;
wire net10176;
wire net9204;
wire net9200;
wire net9199;
wire net9197;
wire net9195;
wire net9194;
wire net9193;
wire net9190;
wire net9188;
wire net11323;
wire net9185;
wire net9183;
wire net10506;
wire net9182;
wire net9536;
wire net9181;
wire net9180;
wire net9178;
wire net9176;
wire net9175;
wire net9171;
wire net9167;
wire net9166;
wire net9165;
wire net9164;
wire net9161;
wire net9160;
wire net9159;
wire net9158;
wire net9258;
wire net9157;
wire net9156;
wire net11103;
wire net9154;
wire net9153;
wire net9152;
wire net9151;
wire net11435;
wire net9147;
wire net9146;
wire net9145;
wire net9144;
wire net10447;
wire net9142;
wire net9141;
wire net9139;
wire net9136;
wire net9133;
wire net9132;
wire net9131;
wire net9130;
wire net9967;
wire net9126;
wire net9116;
wire net9174;
wire net9114;
wire net9112;
wire net9108;
wire net9107;
wire net9106;
wire net9105;
wire net9103;
wire net9100;
wire net9099;
wire net9095;
wire net9091;
wire net9090;
wire net9089;
wire net9088;
wire net9087;
wire net9674;
wire net9086;
wire net9084;
wire net9083;
wire net9081;
wire net9080;
wire net9076;
wire net9075;
wire net9488;
wire net9074;
wire net9073;
wire net9071;
wire net9069;
wire net9068;
wire net9063;
wire net9061;
wire net9059;
wire net9058;
wire net9057;
wire net9056;
wire net9710;
wire net9054;
wire net9053;
wire net9052;
wire net9051;
wire net9050;
wire net9046;
wire net9989;
wire net9045;
wire net9040;
wire net9039;
wire net9038;
wire net11542;
wire net9035;
wire net9032;
wire net9029;
wire net9027;
wire net9026;
wire net9020;
wire net9019;
wire net9018;
wire net9016;
wire net9015;
wire net10504;
wire net9014;
wire net9013;
wire net9011;
wire net9010;
wire net9007;
wire net9005;
wire net9463;
wire net9004;
wire net9003;
wire net9002;
wire net9001;
wire net9000;
wire net8998;
wire net10359;
wire net8997;
wire net8996;
wire net8995;
wire net8993;
wire net8992;
wire net8991;
wire net8989;
wire net8986;
wire net8984;
wire net8983;
wire net8982;
wire net8980;
wire net9475;
wire net8978;
wire net8976;
wire net8975;
wire net8974;
wire net8973;
wire net8972;
wire net10543;
wire net8970;
wire net11334;
wire net8969;
wire net11278;
wire net8968;
wire net8966;
wire net8965;
wire net8961;
wire net8959;
wire net8958;
wire net8956;
wire net8954;
wire net8953;
wire net11574;
wire net8946;
wire net8945;
wire net8941;
wire net8940;
wire net8939;
wire net8937;
wire net10312;
wire net8934;
wire net8927;
wire net9630;
wire net8924;
wire net8921;
wire net9155;
wire net8920;
wire net8919;
wire net8917;
wire net8915;
wire net8913;
wire net8905;
wire net8903;
wire net8902;
wire net8901;
wire net8900;
wire net8899;
wire net8897;
wire net8895;
wire net8893;
wire net11038;
wire net8890;
wire net8889;
wire net8887;
wire net8885;
wire net8884;
wire net8882;
wire net9238;
wire net8880;
wire net8877;
wire net8876;
wire net8875;
wire net8873;
wire net8871;
wire net8870;
wire net8869;
wire net11573;
wire net8868;
wire net8867;
wire net8865;
wire net8863;
wire net8862;
wire net8861;
wire net10958;
wire net8860;
wire net8858;
wire net10593;
wire net8857;
wire net8856;
wire net8864;
wire net8855;
wire net8854;
wire net8853;
wire net8852;
wire net8851;
wire net8850;
wire net8849;
wire net8845;
wire net8844;
wire net8838;
wire net8837;
wire net8836;
wire net9055;
wire net8831;
wire net9806;
wire net8827;
wire net8826;
wire net8822;
wire net8821;
wire net8820;
wire net8819;
wire net8816;
wire net10442;
wire net10241;
wire net8814;
wire net8812;
wire net8811;
wire net8810;
wire net8809;
wire net8808;
wire net8806;
wire net8803;
wire net11092;
wire net8802;
wire net8799;
wire net8798;
wire net8796;
wire net8795;
wire net10388;
wire net9043;
wire net8791;
wire net8787;
wire net8786;
wire net8785;
wire net8784;
wire net11085;
wire net8782;
wire net8780;
wire net8779;
wire net8777;
wire net10081;
wire net8776;
wire net8769;
wire net8768;
wire net8766;
wire net8764;
wire net8763;
wire net9752;
wire net8762;
wire net8761;
wire net8760;
wire net8758;
wire net8753;
wire net8751;
wire net8750;
wire net8749;
wire net8747;
wire net8746;
wire net8745;
wire net8744;
wire net8741;
wire out12;
wire net8740;
wire net8739;
wire net8738;
wire net8737;
wire net8736;
wire net8735;
wire out14;
wire net8733;
wire net8732;
wire net8731;
wire out22;
wire net8728;
wire net10140;
wire net8727;
wire net8726;
wire net10530;
wire net8725;
wire net10178;
wire net8724;
wire net8723;
wire net9828;
wire net8722;
wire net8721;
wire net8720;
wire net8719;
wire net8717;
wire net9784;
wire out18;
wire net8715;
wire net8714;
wire net8713;
wire net8712;
wire net8805;
wire net8710;
wire out11;
wire net8708;
wire net8707;
wire net8705;
wire net8704;
wire net8702;
wire net8701;
wire net8699;
wire net8696;
wire net10963;
wire net8695;
wire net8693;
wire out6;
wire net8692;
wire net8691;
wire net8689;
wire net8918;
wire net8688;
wire net8686;
wire net8683;
wire net8682;
wire net9490;
wire net8681;
wire net8680;
wire net8678;
wire net8677;
wire net8675;
wire net8673;
wire net8672;
wire net8671;
wire net8669;
wire net8668;
wire net8667;
wire net8666;
wire net8665;
wire net8661;
wire net8660;
wire net10716;
wire net10084;
wire net8658;
wire net8653;
wire net8652;
wire net8651;
wire net8648;
wire net8646;
wire net9170;
wire net8644;
wire net8643;
wire net8642;
wire net8641;
wire net8639;
wire net10529;
wire net8638;
wire net8718;
wire net8637;
wire net8636;
wire net8635;
wire net8634;
wire net9192;
wire net8633;
wire net8632;
wire net8631;
wire net11028;
wire net8628;
wire net10660;
wire net8626;
wire net8625;
wire net10741;
wire net8624;
wire net8623;
wire net8621;
wire net8619;
wire net8615;
wire net11183;
wire net8874;
wire net8613;
wire net8611;
wire net8981;
wire net8607;
wire net8606;
wire net8605;
wire net8600;
wire net8598;
wire net8597;
wire net8589;
wire net8588;
wire net10882;
wire net8587;
wire net10148;
wire net8585;
wire net8584;
wire net8971;
wire net8580;
wire net8579;
wire net8577;
wire net9875;
wire net8576;
wire net8574;
wire net8572;
wire net8571;
wire net8570;
wire net8569;
wire net8568;
wire net11098;
wire net8567;
wire net8564;
wire net8560;
wire net8558;
wire net8556;
wire net8555;
wire net8554;
wire net8553;
wire net8552;
wire net9892;
wire net8551;
wire net11145;
wire net8911;
wire net8549;
wire net8547;
wire net8546;
wire net11229;
wire net8545;
wire net8544;
wire net8929;
wire net8541;
wire net8539;
wire net8538;
wire net8534;
wire net8530;
wire net9371;
wire net8529;
wire net8528;
wire net8527;
wire net10012;
wire net8526;
wire net8525;
wire net8524;
wire net8815;
wire net8521;
wire net10437;
wire net8520;
wire net8519;
wire net8518;
wire net8513;
wire net8512;
wire net10345;
wire net9225;
wire net8510;
wire net8509;
wire net8507;
wire net8498;
wire net8497;
wire net9840;
wire net8495;
wire net8493;
wire net8492;
wire net11093;
wire net8489;
wire net8488;
wire net8486;
wire net8480;
wire net8479;
wire net10247;
wire net8478;
wire net11272;
wire net8477;
wire net8475;
wire net11214;
wire net8474;
wire net8471;
wire net8469;
wire net8468;
wire net8466;
wire net8462;
wire net8460;
wire net11012;
wire net8459;
wire net8458;
wire net8456;
wire net8523;
wire net8455;
wire net8454;
wire net8453;
wire net8452;
wire net8450;
wire net8449;
wire net8444;
wire net8442;
wire net8438;
wire net8437;
wire net8434;
wire net8433;
wire net8432;
wire net8429;
wire net8842;
wire net8428;
wire net10586;
wire net8427;
wire net8426;
wire net8425;
wire net8423;
wire net8421;
wire net8418;
wire net8417;
wire net8414;
wire net8413;
wire net8412;
wire net8411;
wire net8410;
wire net8409;
wire net8781;
wire net8408;
wire net8407;
wire net8406;
wire net8405;
wire net8404;
wire net8400;
wire net8397;
wire net8396;
wire net8395;
wire net8394;
wire net8391;
wire net8390;
wire net8389;
wire net8388;
wire net11327;
wire net8387;
wire net8382;
wire net8381;
wire net8378;
wire net9955;
wire net8377;
wire net8374;
wire net8372;
wire net8371;
wire net8369;
wire net8368;
wire net8367;
wire net8366;
wire net8365;
wire net8363;
wire net8362;
wire net8360;
wire net8358;
wire net8355;
wire net8353;
wire net10237;
wire net8350;
wire net8348;
wire net9522;
wire net8347;
wire net8685;
wire net8345;
wire net9374;
wire net8344;
wire net8343;
wire net8342;
wire net8341;
wire net8339;
wire net9111;
wire net8337;
wire net8335;
wire net10596;
wire net8332;
wire net9654;
wire net8331;
wire net8330;
wire net8329;
wire net8328;
wire net8326;
wire net8323;
wire net11410;
wire net8322;
wire net8321;
wire out20;
wire net8319;
wire net8318;
wire net8317;
wire net8316;
wire net8314;
wire net9030;
wire net8312;
wire net8306;
wire net8304;
wire net11360;
wire net8301;
wire net8300;
wire net8297;
wire net8296;
wire net8295;
wire net8292;
wire net8288;
wire net11389;
wire net8286;
wire net8284;
wire net8283;
wire net8281;
wire net8280;
wire net8279;
wire net8276;
wire net8273;
wire net8272;
wire net8271;
wire net10230;
wire net8269;
wire net8266;
wire net8265;
wire net8264;
wire net8263;
wire net8261;
wire net9233;
wire net8260;
wire net8357;
wire net8257;
wire net8254;
wire net8253;
wire net8252;
wire net8249;
wire net10036;
wire net8247;
wire net8245;
wire net8244;
wire net8242;
wire net8241;
wire net8240;
wire net8239;
wire net8238;
wire net8236;
wire net8235;
wire net8234;
wire net8232;
wire net8231;
wire net10177;
wire net8227;
wire net8226;
wire net8225;
wire net8223;
wire net8222;
wire net8220;
wire net8219;
wire net8218;
wire net8217;
wire net8216;
wire net8213;
wire net8212;
wire net8210;
wire net9279;
wire net8209;
wire net8208;
wire net10386;
wire net8207;
wire net8206;
wire net8205;
wire net8203;
wire net8202;
wire net11128;
wire net8201;
wire net11424;
wire net8199;
wire net8198;
wire net8754;
wire net8197;
wire net8196;
wire net8195;
wire net11169;
wire net8193;
wire net8191;
wire net8190;
wire net11366;
wire net8188;
wire net8187;
wire net8186;
wire net10916;
wire net8185;
wire net8183;
wire net8179;
wire net8178;
wire net8175;
wire net9187;
wire net8172;
wire net8823;
wire net8168;
wire net8166;
wire net8165;
wire net8164;
wire net8161;
wire net8159;
wire net8158;
wire net9605;
wire net8157;
wire net8156;
wire net8155;
wire net8153;
wire net11269;
wire net8516;
wire net8152;
wire net10338;
wire net8150;
wire net8149;
wire net8148;
wire net9713;
wire net8146;
wire net8145;
wire net8144;
wire net8143;
wire net8142;
wire net8140;
wire net8139;
wire net8138;
wire net9493;
wire net8136;
wire net8129;
wire net8128;
wire net8127;
wire net8125;
wire net8124;
wire net8123;
wire net8119;
wire net8118;
wire net8117;
wire net8114;
wire net10194;
wire net8113;
wire net8112;
wire net8448;
wire net8110;
wire net10618;
wire net8109;
wire net8106;
wire net8105;
wire net8101;
wire net8100;
wire net8097;
wire net8096;
wire net8095;
wire net8093;
wire net10486;
wire net8092;
wire net9366;
wire net8087;
wire net8084;
wire net9286;
wire net8083;
wire net8082;
wire net10844;
wire net9885;
wire net8081;
wire net10200;
wire net8080;
wire net8077;
wire net8076;
wire net9701;
wire net8075;
wire net8074;
wire net8073;
wire net8069;
wire net8068;
wire net8066;
wire net8063;
wire net8062;
wire net8060;
wire net8058;
wire net8057;
wire net8055;
wire net8051;
wire net8050;
wire net8049;
wire net8048;
wire net8047;
wire net8046;
wire net8044;
wire net8043;
wire net8042;
wire net8040;
wire net8039;
wire net8035;
wire net11301;
wire net8034;
wire net8032;
wire net10415;
wire net8788;
wire net8030;
wire net8029;
wire net8028;
wire net8027;
wire net8026;
wire net9963;
wire net8025;
wire net8024;
wire net8023;
wire net8021;
wire net8018;
wire net8017;
wire net8016;
wire net8015;
wire net8012;
wire net8011;
wire net8009;
wire net8007;
wire net11094;
wire net10355;
wire net8006;
wire net8005;
wire net11110;
wire net8004;
wire net8003;
wire net8002;
wire net8001;
wire net7999;
wire net7997;
wire net7996;
wire net11407;
wire net10123;
wire net8496;
wire net7994;
wire net7993;
wire net7991;
wire net10387;
wire net7990;
wire net7989;
wire net7988;
wire net7986;
wire net7985;
wire net7983;
wire net7980;
wire net7977;
wire net7974;
wire net7973;
wire net7970;
wire net7960;
wire net7958;
wire net7954;
wire net7953;
wire net7950;
wire net7949;
wire net9322;
wire net7948;
wire net11050;
wire net7944;
wire net8305;
wire net7943;
wire net7939;
wire net7937;
wire net7935;
wire net8354;
wire net7934;
wire net7933;
wire net7932;
wire net7930;
wire net7929;
wire net7928;
wire net7926;
wire net7925;
wire net7924;
wire net7923;
wire net7921;
wire net7920;
wire net7919;
wire net7917;
wire net7915;
wire net7914;
wire net7913;
wire net11217;
wire net9287;
wire net7912;
wire net7911;
wire net7910;
wire net9666;
wire net7909;
wire net10630;
wire net7908;
wire net7906;
wire net7905;
wire net11014;
wire net7902;
wire net7892;
wire net7891;
wire net7890;
wire net7889;
wire net7887;
wire net7884;
wire net7881;
wire net7879;
wire net8938;
wire net7878;
wire net7876;
wire net7874;
wire net7873;
wire net7871;
wire net9191;
wire net7870;
wire net7869;
wire out17;
wire net7865;
wire net7864;
wire net7863;
wire net7862;
wire net7861;
wire net8684;
wire net7860;
wire net7857;
wire net8091;
wire net7855;
wire net7852;
wire net7850;
wire net7849;
wire net7848;
wire net7847;
wire net7845;
wire net7843;
wire net7841;
wire net7840;
wire net7836;
wire net7833;
wire net7832;
wire net7824;
wire net7823;
wire net7822;
wire net7816;
wire net7814;
wire net11256;
wire net7813;
wire net7812;
wire net7811;
wire net7810;
wire net7809;
wire net7806;
wire net7803;
wire net7802;
wire net7797;
wire net7796;
wire net7795;
wire net7794;
wire net10418;
wire net7791;
wire net7790;
wire net7789;
wire net7787;
wire net7786;
wire net7785;
wire net7781;
wire net7779;
wire net7777;
wire net7776;
wire net7772;
wire net7771;
wire net7770;
wire net7769;
wire net7767;
wire net7765;
wire net9633;
wire net7763;
wire net7762;
wire net7761;
wire net8916;
wire net7760;
wire net7759;
wire net9644;
wire net7758;
wire net7756;
wire net11551;
wire net7755;
wire net7754;
wire net7753;
wire net10120;
wire net7752;
wire net7984;
wire net7751;
wire net7749;
wire net7748;
wire net7746;
wire net7745;
wire net7743;
wire net7742;
wire net7740;
wire net7737;
wire net7733;
wire net7732;
wire net7731;
wire net10458;
wire net7730;
wire net10951;
wire net7729;
wire net7726;
wire net7725;
wire net7724;
wire net7723;
wire net7721;
wire net7719;
wire net7715;
wire net7714;
wire net7712;
wire net7711;
wire net7710;
wire net7708;
wire net7707;
wire net7706;
wire net7704;
wire net7703;
wire net7699;
wire net9851;
wire net7696;
wire out19;
wire net7694;
wire net7693;
wire net11535;
wire net7691;
wire net7688;
wire net7687;
wire net7686;
wire net7679;
wire net7678;
wire net7784;
wire net7675;
wire net7674;
wire net7671;
wire net7670;
wire net7669;
wire net7668;
wire net7666;
wire net7665;
wire net7663;
wire net7662;
wire net7660;
wire net7659;
wire net10470;
wire net7656;
wire net7655;
wire net7654;
wire net7653;
wire net7652;
wire net7651;
wire net8988;
wire net7648;
wire net9260;
wire net7647;
wire net7645;
wire net7644;
wire net7643;
wire net7642;
wire net10929;
wire net8550;
wire net7641;
wire net7640;
wire net7636;
wire net7634;
wire net7633;
wire net7632;
wire net7631;
wire net7629;
wire net10480;
wire net7628;
wire net7627;
wire net7626;
wire net7625;
wire net7624;
wire net10143;
wire net7621;
wire net7619;
wire net7617;
wire net7615;
wire net7614;
wire net9025;
wire net7609;
wire net7607;
wire net7605;
wire net8752;
wire net7603;
wire net7601;
wire net11109;
wire net7600;
wire net7598;
wire net7595;
wire net7594;
wire net7593;
wire net11587;
wire net7592;
wire net7591;
wire net9771;
wire net7590;
wire net8385;
wire net7588;
wire net7587;
wire net7586;
wire net7585;
wire net7584;
wire net7582;
wire net7581;
wire net7579;
wire net9335;
wire net7577;
wire net7572;
wire net9113;
wire net7571;
wire net7570;
wire net7569;
wire net7568;
wire net7566;
wire net7565;
wire net7564;
wire net7562;
wire net7561;
wire net7560;
wire net7559;
wire net8131;
wire net7558;
wire net11181;
wire net7556;
wire net9705;
wire net7554;
wire net7553;
wire net7549;
wire net9717;
wire net7547;
wire net10639;
wire net7546;
wire net7545;
wire net7543;
wire net7541;
wire net7540;
wire net7539;
wire net9586;
wire net7538;
wire net7537;
wire net7956;
wire net7536;
wire net7535;
wire net7533;
wire net7531;
wire net10720;
wire net7530;
wire net7529;
wire net7527;
wire net9611;
wire net7526;
wire net7525;
wire net7523;
wire net7522;
wire net7521;
wire net11289;
wire net7520;
wire net7519;
wire net9669;
wire net7518;
wire net7517;
wire net7516;
wire net7514;
wire net7510;
wire net7509;
wire net8102;
wire net7508;
wire net7507;
wire net7505;
wire net7503;
wire net7502;
wire net7501;
wire net7500;
wire net10147;
wire net8979;
wire net7499;
wire net7498;
wire net7657;
wire net7497;
wire net7493;
wire net11045;
wire net10488;
wire net7489;
wire net10678;
wire net7488;
wire net3712;
wire net10603;
wire net3650;
wire net5066;
wire net5427;
wire net3699;
wire net4859;
wire net3697;
wire net7427;
wire net10644;
wire net3692;
wire net3687;
wire net11095;
wire net3684;
wire net4757;
wire net3678;
wire net3673;
wire net2661;
wire net3672;
wire net4673;
wire net8338;
wire net5036;
wire net11362;
wire net1050;
wire net3670;
wire net9022;
wire net3669;
wire net6666;
wire net3662;
wire net3657;
wire net10570;
wire net4219;
wire net8888;
wire net5980;
wire net7194;
wire net6390;
wire net3648;
wire net3641;
wire net1859;
wire net3637;
wire net4378;
wire net3635;
wire net8103;
wire net3622;
wire net324;
wire net3615;
wire net3609;
wire net649;
wire net6312;
wire net9079;
wire net3601;
wire net3597;
wire net3596;
wire net3590;
wire net3695;
wire net7859;
wire net4122;
wire net3588;
wire net3390;
wire net2119;
wire net3584;
wire net60;
wire net3582;
wire net3578;
wire net3575;
wire net3574;
wire net3570;
wire net4709;
wire net3567;
wire net3559;
wire net2665;
wire net3557;
wire net3556;
wire net1002;
wire net4495;
wire net3129;
wire net377;
wire net3548;
wire net8832;
wire net3660;
wire net5247;
wire net3546;
wire net2380;
wire net3545;
wire net9569;
wire net8104;
wire net3544;
wire net8593;
wire net6638;
wire net3543;
wire net7268;
wire net9933;
wire net3539;
wire net3538;
wire net3536;
wire net4159;
wire net8346;
wire net3535;
wire net3529;
wire net2047;
wire net3525;
wire net7410;
wire net3523;
wire net3521;
wire net10833;
wire net5119;
wire net3517;
wire net7271;
wire net7931;
wire net3512;
wire net3175;
wire net9138;
wire net3511;
wire net3509;
wire net4564;
wire net11053;
wire net6676;
wire net3508;
wire net3507;
wire net9740;
wire net3502;
wire net3500;
wire net3494;
wire net919;
wire net7196;
wire net8470;
wire net3493;
wire net5719;
wire net3491;
wire net3489;
wire net10007;
wire net329;
wire net3488;
wire net8908;
wire net7311;
wire net3487;
wire net3532;
wire net3486;
wire net3485;
wire net3484;
wire net3480;
wire net4321;
wire net3478;
wire net3476;
wire net10826;
wire net2043;
wire net9033;
wire net3473;
wire net571;
wire net3469;
wire net3466;
wire net3455;
wire net3451;
wire net8303;
wire net3260;
wire net3649;
wire net3449;
wire net5042;
wire net8022;
wire net5709;
wire net3444;
wire net2461;
wire net3442;
wire net3440;
wire net3439;
wire net144;
wire net3519;
wire net872;
wire net5099;
wire net6791;
wire net3426;
wire net8603;
wire net2003;
wire net6715;
wire net3427;
wire net3542;
wire net9328;
wire net3423;
wire net3419;
wire net4987;
wire net3688;
wire net171;
wire net4354;
wire net3638;
wire net11079;
wire net8536;
wire net3411;
wire net2884;
wire net3410;
wire net3408;
wire net1343;
wire net10555;
wire net10350;
wire net6850;
wire net11490;
wire net3547;
wire net3406;
wire net8189;
wire net135;
wire net3401;
wire net7616;
wire net3396;
wire net3210;
wire net3394;
wire net3387;
wire net5745;
wire net3384;
wire net3382;
wire net3380;
wire net3377;
wire net7513;
wire net6701;
wire net9292;
wire net3376;
wire net3366;
wire net3370;
wire net7428;
wire net3369;
wire net10854;
wire net9124;
wire net3367;
wire net3363;
wire net1951;
wire net7285;
wire net9115;
wire net3360;
wire net621;
wire net5422;
wire net3354;
wire net1870;
wire net3350;
wire net3345;
wire net5930;
wire net9854;
wire net4533;
wire net3634;
wire net3341;
wire net7183;
wire net3339;
wire net5845;
wire net3336;
wire net10914;
wire net354;
wire net3330;
wire net3327;
wire net10636;
wire net1054;
wire net10212;
wire net6551;
wire net3326;
wire net3325;
wire net9148;
wire net3323;
wire net5533;
wire net11496;
wire net3318;
wire net7804;
wire net4881;
wire net3316;
wire net1321;
wire net3314;
wire net1702;
wire net3302;
wire net3294;
wire net9273;
wire net3288;
wire net3286;
wire net3284;
wire net581;
wire net11439;
wire net7415;
wire net3921;
wire net3280;
wire net2894;
wire net3589;
wire net3691;
wire net5590;
wire net8038;
wire net3278;
wire net2687;
wire net10738;
wire net3277;
wire net3275;
wire net4097;
wire net11577;
wire net9541;
wire net3658;
wire net10499;
wire net3257;
wire net2284;
wire net7220;
wire net11213;
wire net3252;
wire net3246;
wire net3234;
wire net3240;
wire net3239;
wire net5808;
wire net7269;
wire in24;
wire net4645;
wire net7416;
wire net3235;
wire net6464;
wire net3232;
wire net3230;
wire net532;
wire net5925;
wire net3228;
wire net3149;
wire net3227;
wire net5044;
wire net3225;
wire net11068;
wire net3224;
wire net3438;
wire net10769;
wire net7695;
wire net1451;
wire net8793;
wire net3219;
wire net3218;
wire net5214;
wire net5183;
wire net3211;
wire net3352;
wire net8336;
wire net5697;
wire net7075;
wire net3207;
wire net2852;
wire net9919;
wire net7286;
wire net11196;
wire net3198;
wire net3193;
wire net11118;
wire net6500;
wire net3191;
wire net10635;
wire net3186;
wire net3184;
wire net4949;
wire net3180;
wire net7267;
wire net3647;
wire net3177;
wire net3173;
wire net7727;
wire net3169;
wire net9972;
wire net9810;
wire net1060;
wire net3165;
wire net3498;
wire net3157;
wire net8833;
wire net3375;
wire net8472;
wire net147;
wire net3145;
wire net3143;
wire net3141;
wire net3140;
wire net3137;
wire net3134;
wire net3130;
wire net3126;
wire net8771;
wire net2091;
wire net533;
wire net10615;
wire net5789;
wire net6923;
wire net7018;
wire net3160;
wire net6275;
wire net3121;
wire net1918;
wire net10756;
wire net3112;
wire net126;
wire net3111;
wire net8663;
wire net7511;
wire net3067;
wire net2981;
wire net8839;
wire net3110;
wire net5123;
wire net3109;
wire net3102;
wire net224;
wire net836;
wire net5999;
wire net5375;
wire net3097;
wire net9684;
wire net3321;
wire net3096;
wire net8542;
wire net8464;
wire net749;
wire net2783;
wire net7998;
wire net3459;
wire net5815;
wire net7006;
wire net3088;
wire net7242;
wire net10895;
wire net7567;
wire net3125;
wire net3526;
wire net7927;
wire net5683;
wire net3085;
wire net1175;
wire net2560;
wire net3083;
wire net8215;
wire net2435;
wire net10641;
wire net3808;
wire net3698;
wire net3082;
wire net3081;
wire net2565;
wire net11341;
wire net3076;
wire net3215;
wire net7151;
wire net3071;
wire net9382;
wire net3949;
wire net3070;
wire net11397;
wire net3068;
wire net4842;
wire net6767;
wire net3600;
wire net7306;
wire net3058;
wire net2138;
wire net3057;
wire net2211;
wire net9129;
wire net574;
wire net3431;
wire net3055;
wire net3492;
wire net3053;
wire net5876;
wire net3049;
wire net3047;
wire net8532;
wire net7244;
wire net9217;
wire net3042;
wire net11105;
wire net3039;
wire net6528;
wire net11402;
wire net9214;
wire net3036;
wire net3035;
wire net3099;
wire net1258;
wire net3034;
wire net3032;
wire net3030;
wire net10023;
wire net7524;
wire net1080;
wire net3029;
wire net10308;
wire net3028;
wire net3023;
wire net2962;
wire net3021;
wire net3017;
wire net1663;
wire net3016;
wire net9355;
wire net5554;
wire net8932;
wire net3015;
wire net847;
wire net11087;
wire net3014;
wire net4414;
wire net9450;
wire net3011;
wire net3077;
wire net10904;
wire net3010;
wire net5794;
wire net8649;
wire net3006;
wire net411;
wire net10372;
wire net6852;
wire net11405;
wire net3005;
wire net3004;
wire net3003;
wire net1704;
wire net11143;
wire net9064;
wire net3002;
wire net3000;
wire net2996;
wire net3158;
wire net7131;
wire net1525;
wire net916;
wire net2989;
wire net11361;
wire net9767;
wire net3187;
wire net2022;
wire net5200;
wire net6740;
wire out8;
wire net2987;
wire net1830;
wire net6770;
wire net6251;
wire net2979;
wire net2978;
wire net159;
wire net2975;
wire net10984;
wire net10728;
wire net2972;
wire net2730;
wire net326;
wire net10263;
wire net6700;
wire net7684;
wire net2971;
wire net4955;
wire net3562;
wire net4191;
wire net2969;
wire net3481;
wire net2968;
wire net2967;
wire net1022;
wire net287;
wire net3059;
wire net3118;
wire net10994;
wire net7176;
wire net2954;
wire net2863;
wire net10360;
wire net9247;
wire net2509;
wire net6044;
wire net2950;
wire net2058;
wire net5520;
wire net3458;
wire net2949;
wire net792;
wire net2946;
wire net2714;
wire net2681;
wire net6721;
wire net2941;
wire net2940;
wire net8251;
wire net2939;
wire net11006;
wire net2938;
wire net11135;
wire net2936;
wire net7894;
wire net753;
wire net2932;
wire net2930;
wire net6782;
wire net11232;
wire net6858;
wire net11350;
wire net2928;
wire net9245;
wire net5767;
wire net2923;
wire net2921;
wire net2918;
wire net2917;
wire net2915;
wire net1442;
wire net3679;
wire net6584;
wire net2913;
wire net3859;
wire net7155;
wire net5225;
wire net8964;
wire net4032;
wire net2908;
wire net4094;
wire net2903;
wire net4135;
wire net2902;
wire net9122;
wire net2436;
wire net5492;
wire net7918;
wire net4096;
wire net5265;
wire net534;
wire net10421;
wire net3616;
wire net3533;
wire net2891;
wire net11154;
wire net6354;
wire net2886;
wire net5222;
wire net1664;
wire net2878;
wire net2195;
wire net1705;
wire net2877;
wire net8923;
wire net8514;
wire net6667;
wire net10941;
wire net6895;
wire net2875;
wire net1256;
wire net3074;
wire net2872;
wire net7250;
wire net10032;
wire net2870;
wire net4238;
wire net2869;
wire net4437;
wire net4475;
wire net4560;
wire net2595;
wire net8610;
wire net2516;
wire net1992;
wire net9085;
wire net6657;
wire net2847;
wire net461;
wire net6897;
wire net2836;
wire net35;
wire net5199;
wire net4652;
wire net5548;
wire net2988;
wire net2871;
wire net2834;
wire net10753;
wire net8262;
wire net2832;
wire net2831;
wire net4978;
wire net7309;
wire net2829;
wire net3447;
wire net2752;
wire net9097;
wire net5368;
wire net2826;
wire net2818;
wire net3714;
wire net6357;
wire net2817;
wire net4128;
wire net7971;
wire net2811;
wire net3116;
wire net2807;
wire net5561;
wire net7900;
wire net5735;
wire net2806;
wire net6496;
wire net3467;
wire net8494;
wire net2705;
wire net2801;
wire net2800;
wire net5443;
wire net9203;
wire net2798;
wire net2796;
wire net9813;
wire net3655;
wire net2793;
wire net9567;
wire net3342;
wire net7107;
wire net2790;
wire net8379;
wire net1631;
wire net3710;
wire net1568;
wire net4512;
wire net3995;
wire net3133;
wire net7310;
wire net2784;
wire net2781;
wire net8907;
wire net3831;
wire net4138;
wire net2402;
wire net2777;
wire net3162;
wire net2145;
wire net9270;
wire net146;
wire net11563;
wire net2952;
wire net11211;
wire net11104;
wire net802;
wire net2767;
wire net2766;
wire net5588;
wire net3306;
wire net9639;
wire net6689;
wire net9577;
wire net6806;
wire net2763;
wire net945;
wire net4085;
wire net5372;
wire net5432;
wire net11273;
wire net2758;
wire net2756;
wire net2749;
wire net923;
wire net3961;
wire net11409;
wire net2747;
wire net9465;
wire net9267;
wire net690;
wire net3203;
wire net9249;
wire net1601;
wire net2743;
wire net10761;
wire net3950;
wire net6240;
wire net5193;
wire net6601;
wire net2742;
wire net4666;
wire net8620;
wire net5801;
wire net6272;
wire net3388;
wire net2368;
wire net3528;
wire net585;
wire net3212;
wire net5397;
wire net2738;
wire net2495;
wire net1173;
wire net4323;
wire net10606;
wire net7324;
wire net2733;
wire net6028;
wire net7701;
wire net2000;
wire net3276;
wire net7372;
wire net2723;
wire net8912;
wire net2722;
wire net2720;
wire net10573;
wire net1215;
wire net5480;
wire net11222;
wire net2707;
wire net5675;
wire net6569;
wire net2700;
wire net777;
wire net3980;
wire net2694;
wire net3516;
wire net1508;
wire net9965;
wire net2622;
wire net7354;
wire net1197;
wire net2691;
wire net2689;
wire out4;
wire net795;
wire net2684;
wire net10196;
wire net8508;
wire net2680;
wire net3348;
wire net2497;
wire net2679;
wire net2674;
wire net1459;
wire net2873;
wire net2760;
wire net2666;
wire net10034;
wire net3612;
wire net3221;
wire net11303;
wire net5313;
wire net2663;
wire net3811;
wire net9426;
wire net105;
wire net2659;
wire net10731;
wire net2658;
wire net10026;
wire net407;
wire net3268;
wire net4808;
wire net2657;
wire net2653;
wire net2381;
wire net2652;
wire net2650;
wire net1934;
wire net2649;
wire net9023;
wire net2648;
wire net1786;
wire net1037;
wire net2791;
wire net2642;
wire net454;
wire net4528;
wire net2634;
wire net4608;
wire net2631;
wire net2626;
wire net2772;
wire net2625;
wire net6280;
wire net10920;
wire net6302;
wire net3202;
wire net4113;
wire net10351;
wire net6979;
wire net4964;
wire net9620;
wire net2620;
wire net9745;
wire net3199;
wire net2618;
wire net626;
wire net6673;
wire net1800;
wire net3346;
wire net231;
wire net3251;
wire net3964;
wire net7034;
wire net9446;
wire net6600;
wire net9137;
wire net2782;
wire net2610;
wire net2603;
wire net11164;
wire net361;
wire net4086;
wire net2601;
wire net2600;
wire net662;
wire net8778;
wire net2596;
wire net3802;
wire net2591;
wire net9530;
wire net276;
wire net8828;
wire net2588;
wire net4819;
wire net2586;
wire net2014;
wire net9451;
wire net2232;
wire net2375;
wire net6123;
wire net2583;
wire net2581;
wire net3775;
wire in17;
wire net9990;
wire net4650;
wire net2579;
wire net2695;
wire net5839;
wire net7961;
wire net3579;
wire net2960;
wire net2576;
wire net2574;
wire net9799;
wire net6922;
wire net2571;
wire net2569;
wire net10851;
wire net9491;
wire net3031;
wire net2568;
wire net1575;
wire net7799;
wire net3153;
wire net10775;
wire net10540;
wire net2655;
wire net4907;
wire net8765;
wire net7623;
wire net6843;
wire net2566;
wire net2563;
wire net10810;
wire net5332;
wire net2561;
wire net6644;
wire net7476;
wire net2557;
wire net2555;
wire net1597;
wire net6793;
wire net2543;
wire net2672;
wire net2542;
wire net2541;
wire net1241;
wire net7612;
wire net5883;
wire net2538;
wire net1544;
wire net5457;
wire net8325;
wire net2536;
wire net7801;
wire net5933;
wire net11384;
wire net2535;
wire net1563;
wire net5098;
wire net10405;
wire net2534;
wire net2532;
wire net2208;
wire net2527;
wire net9904;
wire net1688;
wire net10783;
wire net7965;
wire net3624;
wire net10752;
wire net7898;
wire net2524;
wire net8891;
wire net4747;
wire net6618;
wire net6545;
wire net2521;
wire net2520;
wire net4532;
wire net2519;
wire net2518;
wire net2241;
wire net2517;
wire net3586;
wire net2504;
wire net3247;
wire net1203;
wire net2502;
wire net2500;
wire net2499;
wire net3581;
wire net8543;
wire net3392;
wire net5312;
wire net2491;
wire net2487;
wire net2482;
wire net2956;
wire net5093;
wire net9733;
wire net3560;
wire net6660;
wire net5692;
wire net6542;
wire net2480;
wire net2479;
wire net2478;
wire net7750;
wire net2476;
wire net1592;
wire net8987;
wire net65;
wire net2645;
wire net5245;
wire net1613;
wire net5690;
wire net6619;
wire net5238;
wire net9687;
wire net8485;
wire net2469;
wire net2115;
wire net2896;
wire net734;
wire net2460;
wire net2459;
wire net7302;
wire net2453;
wire net2452;
wire net5022;
wire net2448;
wire net1460;
wire net2660;
wire net8711;
wire net2444;
wire net11337;
wire net7938;
wire net2442;
wire net2233;
wire net2440;
wire net2439;
wire net8935;
wire net2438;
wire net3470;
wire net2842;
wire net2951;
wire net2498;
wire net2033;
wire net2431;
wire net8457;
wire net1888;
wire net8948;
wire net870;
wire net2429;
wire net6532;
wire net2810;
wire net4108;
wire net2425;
wire net2424;
wire net2422;
wire net8825;
wire net4444;
wire net10998;
wire net3155;
wire net208;
wire net4180;
wire net8614;
wire net2421;
wire net604;
wire net10632;
wire net3300;
wire net178;
wire net6745;
wire net2416;
wire net2525;
wire net5067;
wire net2413;
wire net1446;
wire net2412;
wire net2411;
wire net7182;
wire net2408;
wire net7972;
wire net2407;
wire net1914;
wire net912;
wire net2404;
wire net2401;
wire net2400;
wire net4607;
wire net6249;
wire net2399;
wire net2397;
wire net2391;
wire net1477;
wire net2390;
wire net10055;
wire net2389;
wire net2388;
wire net6522;
wire net2386;
wire net2385;
wire net10294;
wire net5806;
wire net1181;
wire net2379;
wire net10872;
wire net2378;
wire net1848;
wire net2377;
wire net3619;
wire net2840;
wire net2271;
wire net1611;
wire net7895;
wire net6720;
wire net2370;
wire net2364;
wire net8578;
wire net1520;
wire net10417;
wire net2362;
wire net4204;
wire net2361;
wire net3850;
wire net7431;
wire net2356;
wire net2353;
wire net2724;
wire net10508;
wire net3803;
wire net2352;
wire net3148;
wire net1139;
wire net10990;
wire net10223;
wire net2351;
wire net9104;
wire net6705;
wire net9714;
wire net2349;
wire net7085;
wire net8293;
wire net2718;
wire net8501;
wire net2347;
wire net2383;
wire net2345;
wire net2858;
wire net2344;
wire net2343;
wire net4250;
wire net8756;
wire net7387;
wire net2338;
wire net5430;
wire net2335;
wire net2334;
wire net9368;
wire net3163;
wire net9425;
wire net2006;
wire net1463;
wire net8465;
wire net3541;
wire net8033;
wire net7738;
wire net7281;
wire net9782;
wire net2326;
wire net9041;
wire net2325;
wire net2317;
wire net5091;
wire net1747;
wire net10289;
wire net8990;
wire net8169;
wire net138;
wire net365;
wire net2312;
wire net9060;
wire net2309;
wire net3413;
wire net7009;
wire net1640;
wire net11344;
wire net3668;
wire net4457;
wire net2302;
wire net1118;
wire net390;
wire net2528;
wire net2296;
wire net10302;
wire net1738;
wire net1030;
wire net10925;
wire net10507;
wire net2292;
wire net10261;
wire net3124;
wire net2291;
wire net6097;
wire net11031;
wire net2290;
wire net762;
wire net5890;
wire net6968;
wire net2307;
wire net6281;
wire net2287;
wire net8361;
wire net5202;
wire net9096;
wire net1909;
wire net3885;
wire net133;
wire net216;
wire net1261;
wire net7417;
wire net2716;
wire net2280;
wire net2846;
wire net2279;
wire net2426;
wire net164;
wire net8067;
wire net2830;
wire net2275;
wire net4011;
wire net2274;
wire net2719;
wire net3269;
wire net5030;
wire net11382;
wire net3623;
wire net2276;
wire net2272;
wire net3305;
wire net6714;
wire net2269;
wire net1596;
wire net2735;
wire net3307;
wire net2263;
wire net5075;
wire net10770;
wire net5670;
wire net2904;
wire net4118;
wire net2262;
wire net2259;
wire net7193;
wire net2252;
wire net2251;
wire net2249;
wire net5984;
wire net2248;
wire net11461;
wire net4790;
wire net2247;
wire net1116;
wire net11199;
wire net11147;
wire net2245;
wire net10880;
wire net2765;
wire net2244;
wire net2243;
wire net6625;
wire net2242;
wire net2240;
wire net3295;
wire net1713;
wire net2238;
wire net2237;
wire net7221;
wire net8789;
wire net179;
wire net1571;
wire net2230;
wire net2229;
wire net8930;
wire net4272;
wire net2277;
wire net7690;
wire net5572;
wire net3066;
wire net5626;
wire net3554;
wire net2226;
wire net4116;
wire net5499;
wire net3310;
wire net2224;
wire net10476;
wire net2222;
wire net11002;
wire net1865;
wire net6178;
wire net2219;
wire net10483;
wire net8504;
wire net2313;
wire net4206;
wire net1822;
wire net6485;
wire net1975;
wire net2204;
wire net10714;
wire net3527;
wire net4196;
wire net5105;
wire net2192;
wire net2191;
wire net2187;
wire net4006;
wire net2184;
wire net5908;
wire net7483;
wire net2182;
wire net2741;
wire net7975;
wire net327;
wire net9065;
wire net3103;
wire net3291;
wire net4844;
wire net2174;
wire net2172;
wire net3836;
wire net7300;
wire net10198;
wire net3522;
wire net2171;
wire net2165;
wire net2164;
wire net2163;
wire net11421;
wire net4775;
wire net2162;
wire net5017;
wire net2161;
wire net1340;
wire net9274;
wire net5607;
wire net6579;
wire net11354;
wire net2160;
wire net1208;
wire net9312;
wire net2157;
wire in5;
wire net396;
wire net2154;
wire net7899;
wire net7231;
wire net7184;
wire net2152;
wire net2151;
wire net3890;
wire net2149;
wire net2144;
wire net10357;
wire net7358;
wire net9482;
wire net2493;
wire net6435;
wire net2142;
wire net9554;
wire net8370;
wire net6595;
wire net2135;
wire net10684;
wire net2134;
wire net9017;
wire net7551;
wire net853;
wire net8461;
wire net3250;
wire net5382;
wire net8645;
wire net8467;
wire net2354;
wire net2822;
wire net2693;
wire net11516;
wire net8403;
wire net5638;
wire net2137;
wire net3643;
wire net2129;
wire net4315;
wire net10158;
wire net9890;
wire net3120;
wire net2126;
wire net5891;
wire net2125;
wire net3436;
wire net1876;
wire net1741;
wire net2123;
wire net219;
wire net2120;
wire net3752;
wire net794;
wire net4363;
wire net1069;
wire net8957;
wire net1365;
wire net6606;
wire net10970;
wire net10614;
wire net7866;
wire net2114;
wire net2113;
wire net2111;
wire net10696;
wire net2108;
wire net2106;
wire net2710;
wire net343;
wire net2105;
wire net8120;
wire net2270;
wire net1809;
wire net10556;
wire net2102;
wire net292;
wire net2881;
wire net11450;
wire net3496;
wire net9994;
wire net2101;
wire net2959;
wire net2097;
wire net2708;
wire net2096;
wire net330;
wire net1219;
wire net5507;
wire net2474;
wire net2094;
wire net9557;
wire net6868;
wire net9956;
wire net2088;
wire net2086;
wire net8380;
wire net3267;
wire net8960;
wire net2508;
wire net10500;
wire net2085;
wire net2215;
wire net6537;
wire net2570;
wire net655;
wire net2084;
wire net2041;
wire net503;
wire net2078;
wire net6248;
wire net2180;
wire net3989;
wire net9523;
wire net8730;
wire net6946;
wire net3237;
wire net2073;
wire net2393;
wire net2072;
wire net2970;
wire net2068;
wire net2064;
wire net5702;
wire net9929;
wire net212;
wire net2061;
wire net9034;
wire net7853;
wire net2060;
wire net4319;
wire net9520;
wire net3308;
wire net2057;
wire net3626;
wire net8627;
wire net2054;
wire net425;
wire net3381;
wire net2769;
wire net1796;
wire net2010;
wire net4329;
wire net2859;
wire net2048;
wire net515;
wire net2045;
wire net2265;
wire net6350;
wire net6908;
wire net2042;
wire net7969;
wire net2039;
wire net2037;
wire net1958;
wire net2032;
wire net2246;
wire net1155;
wire net1429;
wire net7716;
wire net2026;
wire net1170;
wire net4754;
wire net2023;
wire net2725;
wire net177;
wire net2021;
wire net10100;
wire net2210;
wire net1368;
wire net7968;
wire net4415;
wire net6395;
wire net10076;
wire net7867;
wire net2019;
wire net6594;
wire net2018;
wire net2016;
wire net2332;
wire net211;
wire net11070;
wire net6226;
wire net2015;
wire net2776;
wire net8445;
wire net7359;
wire net2007;
wire net9162;
wire net2005;
wire net3248;
wire net2001;
wire net11365;
wire net430;
wire net2098;
wire net1998;
wire net1997;
wire net1853;
wire net750;
wire net5278;
wire net2948;
wire net11481;
wire net6708;
wire net1994;
wire net3762;
wire net6194;
wire net2040;
wire net1993;
wire net2009;
wire net310;
wire net10150;
wire net8311;
wire net6727;
wire net2506;
wire net1991;
wire net6892;
wire net10983;
wire net2104;
wire net763;
wire net3738;
wire net1190;
wire net1989;
wire net6776;
wire net4922;
wire net3080;
wire net1985;
wire net8392;
wire net744;
wire net9941;
wire net1984;
wire net350;
wire net3726;
wire net8951;
wire net4254;
wire net1983;
wire net1291;
wire net3955;
wire net1977;
wire net1308;
wire net11276;
wire net1974;
wire net1754;
wire net4034;
wire net11122;
wire net8174;
wire net255;
wire net11114;
wire net2792;
wire net5576;
wire net2255;
wire net2572;
wire net1466;
wire net2890;
wire net3967;
wire net2505;
wire net5367;
wire net5369;
wire net1967;
wire net1964;
wire net2985;
wire net1961;
wire net2845;
wire net1960;
wire net9481;
wire net6332;
wire net1959;
wire net1956;
wire net2197;
wire net2471;
wire net3416;
wire net6025;
wire net10278;
wire net9173;
wire net2974;
wire net4137;
wire net1948;
wire net1946;
wire net10950;
wire net2510;
wire net1945;
wire net2567;
wire net1943;
wire net1942;
wire net1940;
wire net1939;
wire net10909;
wire net6218;
wire net9624;
wire net8447;
wire net2841;
wire net10768;
wire net1937;
wire net4937;
wire net861;
wire net11532;
wire net9036;
wire net3338;
wire net2823;
wire net2545;
wire net1931;
wire net5031;
wire net9417;
wire net6115;
wire net8134;
wire net5493;
wire net6598;
wire net1923;
wire net1922;
wire net970;
wire net1921;
wire net9485;
wire net5558;
wire net6316;
wire net2214;
wire net1913;
wire net1912;
wire net7378;
wire net4812;
wire net1767;
wire net2933;
wire net8654;
wire net2888;
wire net1903;
wire net8925;
wire net1899;
wire net1897;
wire net8327;
wire net999;
wire net10931;
wire net6429;
wire net1896;
wire net3705;
wire net1555;
wire net4107;
wire net1895;
wire net3090;
wire net1894;
wire net10052;
wire net1889;
wire net6166;
wire net2257;
wire net7606;
wire net7259;
wire net3337;
wire net2585;
wire net1293;
wire net8608;
wire net3279;
wire net2036;
wire net1887;
wire net10617;
wire net10399;
wire net4647;
wire net2398;
wire net1884;
wire net1883;
wire net294;
wire net5749;
wire net1864;
wire net1861;
wire net500;
wire net1857;
wire net1856;
wire net1855;
wire net172;
wire net9028;
wire net4174;
wire net3681;
wire net1854;
wire net10599;
wire net2599;
wire net10868;
wire net1850;
wire net4570;
wire net4948;
wire net2337;
wire net1849;
wire net10393;
wire net10206;
wire net686;
wire net7290;
wire net3371;
wire net1846;
wire net904;
wire net442;
wire net10319;
wire net5192;
wire net1842;
wire net1841;
wire net3209;
wire net4044;
wire net1908;
wire net11111;
wire net1840;
wire net6462;
wire net11140;
wire net1838;
wire net10926;
wire net7573;
wire net1851;
wire net1837;
wire net2503;
wire net5678;
wire net6907;
wire net8994;
wire net1835;
wire net8773;
wire net4422;
wire net1826;
wire net6058;
wire net1556;
wire net5253;
wire net5612;
wire net10281;
wire net1819;
wire net10792;
wire net1817;
wire net3530;
wire net340;
wire net3194;
wire net1813;
wire net3652;
wire net3378;
wire net3084;
wire net1501;
wire net5756;
wire net2261;
wire net3242;
wire net10986;
wire net4839;
wire net2110;
wire net1029;
wire net4802;
wire net3884;
wire net4846;
wire net1811;
wire net313;
wire net4172;
wire net3317;
wire net11387;
wire net10661;
wire net2076;
wire net1806;
wire net5508;
wire net2628;
wire net776;
wire net10491;
wire net2740;
wire net2575;
wire net1802;
wire net5989;
wire net10197;
wire net6467;
wire net3349;
wire net9497;
wire net2494;
wire net11331;
wire net1795;
wire net1318;
wire net6297;
wire net2305;
wire net1792;
wire net9409;
wire net8430;
wire net977;
wire net1791;
wire net2761;
wire net4700;
wire net335;
wire net9367;
wire net6934;
wire net4229;
wire net5823;
wire net5924;
wire net3105;
wire net5556;
wire net7922;
wire net4684;
wire net4863;
wire net7955;
wire net6555;
wire net2704;
wire net9787;
wire net6159;
wire net8151;
wire net1780;
wire net1775;
wire net6976;
wire net3593;
wire net3195;
wire net1654;
wire net1774;
wire net9636;
wire net3503;
wire net2754;
wire net1987;
wire net5674;
wire net10901;
wire net1771;
wire net7335;
wire net1770;
wire net11113;
wire net3362;
wire net1769;
wire net5172;
wire net1768;
wire net8830;
wire net6197;
wire net6960;
wire net8356;
wire net1766;
wire net9800;
wire net1763;
wire net10452;
wire net2816;
wire net2329;
wire net1759;
wire net9143;
wire net4236;
wire net1757;
wire net2481;
wire net2874;
wire net2753;
wire net3233;
wire net1749;
wire net7374;
wire net5621;
wire net11296;
wire net4618;
wire net6531;
wire net2295;
wire net1372;
wire net8170;
wire net114;
wire net8111;
wire net5914;
wire net1742;
wire net5768;
wire net1739;
wire net6451;
wire net4815;
wire net9517;
wire net6574;
wire net3462;
wire net1734;
wire net1733;
wire net2640;
wire net1732;
wire net483;
wire net7916;
wire net1731;
wire net6664;
wire net5288;
wire net1730;
wire net8840;
wire net4280;
wire net4813;
wire net1729;
wire net2731;
wire net1726;
wire net5147;
wire net1725;
wire net4803;
wire net1724;
wire net9942;
wire net5446;
wire net9494;
wire net1723;
wire net116;
wire net28;
wire net1722;
wire net22;
wire net10588;
wire net6838;
wire net7744;
wire net1721;
wire net9272;
wire net8602;
wire net8086;
wire net2892;
wire net1720;
wire net11032;
wire net1716;
wire net578;
wire net11178;
wire net1179;
wire net8070;
wire net5858;
wire net5816;
wire net1040;
wire net3220;
wire net246;
wire net783;
wire net1828;
wire net43;
wire net541;
wire net6604;
wire net4828;
wire net3693;
wire net3037;
wire net8107;
wire net2253;
wire net1941;
wire net6651;
wire net772;
wire net7059;
wire net10751;
wire net2643;
wire net761;
wire net8952;
wire net478;
wire net15;
wire net8383;
wire net4301;
wire net9397;
wire net5025;
wire net746;
wire net168;
wire net2827;
wire net6160;
wire net11514;
wire net738;
wire net10713;
wire net1938;
wire net5560;
wire net3204;
wire net9435;
wire net9285;
wire net1638;
wire net737;
wire net1125;
wire net10819;
wire net2879;
wire net3293;
wire net10972;
wire net5458;
wire net4904;
wire net7327;
wire net9993;
wire net736;
wire net11076;
wire net1785;
wire net414;
wire net5344;
wire net1122;
wire net2696;
wire net7078;
wire net2559;
wire net7462;
wire net730;
wire net4917;
wire net3146;
wire out9;
wire net2617;
wire net728;
wire net3599;
wire net406;
wire net9396;
wire net5624;
wire net1999;
wire net4156;
wire net725;
wire net4517;
wire net808;
wire net2732;
wire net2392;
wire net724;
wire net6546;
wire net1526;
wire net2787;
wire net2220;
wire net721;
wire net10946;
wire net9889;
wire net7315;
wire net3632;
wire net7661;
wire net1315;
wire net1814;
wire net797;
wire net7548;
wire net1502;
wire net4756;
wire net1475;
wire net715;
wire net1100;
wire net1689;
wire net4316;
wire net9461;
wire net1178;
wire net11524;
wire net4708;
wire net3046;
wire net703;
wire net1519;
wire net679;
wire net9550;
wire net1265;
wire net9928;
wire net3552;
wire net700;
wire net11412;
wire net4170;
wire net3666;
wire net699;
wire net1075;
wire net706;
wire net4789;
wire net596;
wire net25;
wire net691;
wire net1488;
wire net5351;
wire net2906;
wire net10037;
wire net676;
wire net3078;
wire net7683;
wire net2258;
wire net6107;
wire net1051;
wire net960;
wire net8894;
wire net8274;
wire net2887;
wire net6641;
wire net693;
wire net2515;
wire net914;
wire net1264;
wire net7379;
wire net2446;
wire net670;
wire net7672;
wire net397;
wire net5387;
wire net7054;
wire net6940;
wire net2668;
wire net1218;
wire net6954;
wire net1656;
wire net4962;
wire net1660;
wire net1773;
wire net648;
wire net842;
wire net153;
wire net644;
wire net1418;
wire net5248;
wire net3008;
wire net1373;
wire net640;
wire net4841;
wire net1827;
wire net5348;
wire net5070;
wire net3389;
wire net1797;
wire net282;
wire net6311;
wire net10541;
wire net7166;
wire net637;
wire net2692;
wire net3977;
wire net2038;
wire net1947;
wire net7261;
wire net238;
wire net1383;
wire net7349;
wire net3024;
wire net579;
wire net2604;
wire net713;
wire net4766;
wire net2083;
wire net707;
wire net559;
wire net5884;
wire net632;
wire net8299;
wire net770;
wire net8949;
wire net2188;
wire net3409;
wire net1331;
wire net4499;
wire net2578;
wire net2651;
wire net631;
wire net611;
wire net9793;
wire net4899;
wire net1146;
wire net617;
wire net986;
wire net1615;
wire net6368;
wire net6816;
wire net7109;
wire net817;
wire net4176;
wire net3504;
wire net3355;
wire net2409;
wire net2544;
wire net603;
wire net9202;
wire net4290;
wire net3063;
wire net1153;
wire net599;
wire net8439;
wire net328;
wire net766;
wire net6707;
wire net3454;
wire net11538;
wire net7026;
wire net1573;
wire net2608;
wire net591;
wire net11479;
wire net996;
wire net6373;
wire net2260;
wire net2973;
wire net4591;
wire net1113;
wire net2475;
wire net587;
wire net934;
wire net1863;
wire net3920;
wire net9401;
wire net1415;
wire net10701;
wire net7698;
wire net6205;
wire net8419;
wire net3608;
wire net5881;
wire net7868;
wire net1560;
wire net650;
wire net7877;
wire net6824;
wire net58;
wire net8484;
wire net3217;
wire net9241;
wire net8843;
wire net5268;
wire net85;
wire net3027;
wire net4266;
wire net9615;
wire net4927;
wire net4347;
wire net7363;
wire net4143;
wire net186;
wire net8259;
wire net3073;
wire net1882;
wire net1393;
wire net9853;
wire net4348;
wire net710;
wire net3249;
wire net4529;
wire net1976;
wire net612;
wire net1010;
wire net957;
wire net5236;
wire net573;
wire net864;
wire net4998;
wire net3060;
wire net4745;
wire net3056;
wire net357;
wire net1965;
wire net768;
wire net1014;
wire net1681;
wire net8977;
wire net247;
wire net1687;
wire net5889;
wire net4282;
wire net564;
wire net3914;
wire net4577;
wire net6879;
wire net2020;
wire net1772;
wire net4498;
wire net189;
wire net5191;
wire net383;
wire net2788;
wire net1673;
wire net3782;
wire net555;
wire net1379;
wire net3737;
wire net553;
wire net2205;
wire net6826;
wire net9044;
wire net2636;
wire net7294;
wire net551;
wire net10407;
wire net8130;
wire net4390;
wire net1063;
wire net549;
wire net10258;
wire net3595;
wire net1428;
wire net6792;
wire net6363;
wire net546;
wire net2580;
wire net6680;
wire net5961;
wire net544;
wire net6353;
wire net3262;
wire net11184;
wire net9410;
wire net4896;
wire net3661;
wire net1;
wire net7385;
wire net10923;
wire net2602;
wire in3;
wire net1270;
wire net4584;
wire net10879;
wire net2584;
wire net896;
wire net11371;
wire net7402;
wire net2029;
wire net535;
wire net3168;
wire net1552;
wire net9453;
wire net2729;
wire net2726;
wire net642;
wire net2159;
wire net659;
wire net830;
wire net3610;
wire net4431;
wire net729;
wire net3379;
wire net823;
wire net1250;
wire net2117;
wire net10726;
wire net1695;
wire net3860;
wire net1886;
wire net1468;
wire net7830;
wire net3445;
wire net98;
wire net524;
wire net4001;
wire net876;
wire net1052;
wire net3587;
wire net3333;
wire net5180;
wire net2079;
wire net9509;
wire net2953;
wire net297;
wire net10006;
wire net8729;
wire net5055;
wire net516;
wire net2779;
wire net1472;
wire net1793;
wire net6982;
wire net8290;
wire net7552;
wire net514;
wire net10732;
wire net8942;
wire net511;
wire net4685;
wire net3618;
wire net1335;
wire net5148;
wire net4151;
wire net685;
wire net107;
wire net2539;
wire net3881;
wire net269;
wire net9652;
wire net346;
wire net8575;
wire net510;
wire net7122;
wire net1233;
wire net1025;
wire net506;
wire net927;
wire net3100;
wire net333;
wire net9466;
wire net3062;
wire net3214;
wire net1927;
wire net975;
wire net1952;
wire net505;
wire net2864;
wire net9804;
wire net8629;
wire net8256;
wire net3550;
wire net6150;
wire net1376;
wire net2630;
wire net1409;
wire net3696;
wire net1437;
wire net1829;
wire net1032;
wire net9595;
wire net8255;
wire net3086;
wire net501;
wire net2931;
wire net3407;
wire net1481;
wire net652;
wire net495;
wire net7364;
wire net494;
wire net988;
wire net11509;
wire net492;
wire net2143;
wire net489;
wire net485;
wire net2745;
wire net985;
wire net488;
wire net10878;
wire net646;
wire net838;
wire net5396;
wire net2170;
wire net475;
wire net6502;
wire net8275;
wire net2209;
wire net639;
wire net674;
wire net525;
wire net3400;
wire net7875;
wire net474;
wire net3094;
wire net4975;
wire net1867;
wire net8834;
wire net473;
wire net10822;
wire net6157;
wire net2955;
wire net1145;
wire net4658;
wire net472;
wire net3331;
wire net3340;
wire net1347;
wire net3101;
wire net3958;
wire net3707;
wire net2616;
wire net3061;
wire net2331;
wire net967;
wire net5346;
wire net6035;
wire net3646;
wire net7051;
wire net1057;
wire net2675;
wire net1567;
wire net1272;
wire net2176;
wire net11469;
wire net10410;
wire net4372;
wire net8014;
wire net780;
wire net7202;
wire net364;
wire net3395;
wire net1266;
wire net8121;
wire net7904;
wire net5097;
wire net6057;
wire net4099;
wire net5582;
wire net283;
wire net6856;
wire net9353;
wire net3289;
wire net10208;
wire net6002;
wire net2737;
wire net3127;
wire net1114;
wire net9066;
wire net3972;
wire net1295;
wire net10444;
wire net2056;
wire net3832;
wire net9408;
wire net3965;
wire net3159;
wire net459;
wire net545;
wire net6003;
wire net4225;
wire net453;
wire net624;
wire net629;
wire net731;
wire net450;
wire net7946;
wire net448;
wire net5559;
wire net1196;
wire net2122;
wire net5363;
wire net5;
wire net10649;
wire net8898;
wire net1012;
wire net4443;
wire net10884;
wire net3285;
wire net3944;
wire net9006;
wire net1074;
wire net2216;
wire net3704;
wire net561;
wire net7484;
wire net444;
wire net8656;
wire net2638;
wire net2071;
wire net1374;
wire net3621;
wire net10389;
wire net8950;
wire net8904;
wire net504;
wire net2997;
wire net336;
wire net280;
wire net8881;
wire net969;
wire net437;
wire net4483;
wire net7764;
wire net3064;
wire net3631;
wire net8926;
wire net162;
wire net11547;
wire net1017;
wire net4787;
wire net10315;
wire net718;
wire net10772;
wire net6725;
wire net2430;
wire net4893;
wire net3095;
wire net5764;
wire net3900;
wire net10383;
wire net8612;
wire net432;
wire net1761;
wire net5294;
wire net8706;
wire net2118;
wire net1645;
wire net428;
wire net774;
wire net556;
wire net3312;
wire net2706;
wire net7487;
wire net771;
wire net5184;
wire net5648;
wire net928;
wire net1336;
wire net1220;
wire net5235;
wire net11483;
wire net3033;
wire net293;
wire net2324;
wire net2107;
wire net11246;
wire net5829;
wire net689;
wire net7218;
wire net422;
wire net1743;
wire clk;
wire net5308;
wire net2637;
wire net3122;
wire net6691;
wire net3576;
wire net4327;
wire net382;
wire net563;
wire net5841;
wire net1188;
wire net3663;
wire net5465;
wire net758;
wire net8650;
wire net2746;
wire net1625;
wire net417;
wire net901;
wire net10547;
wire net2030;
wire net3791;
wire net415;
wire net4389;
wire net5217;
wire net3142;
wire net4781;
wire net412;
wire net748;
wire net1224;
wire net2299;
wire net9118;
wire net702;
wire net5077;
wire net7425;
wire net634;
wire net1981;
wire net3838;
wire net7610;
wire net5879;
wire net554;
wire net4216;
wire net9725;
wire net1192;
wire net6786;
wire net7583;
wire net2597;
wire net3939;
wire net10846;
wire net8071;
wire net3026;
wire net3721;
wire net4454;
wire net11351;
wire net680;
wire net2677;
wire net6442;
wire net6797;
wire net403;
wire net4296;
wire net2066;
wire net2943;
wire net4852;
wire net8878;
wire net7053;
wire net1330;
wire net3216;
wire net3274;
wire net9128;
wire net5131;
wire net854;
wire net10722;
wire net8922;
wire net2656;
wire net4833;
wire net5512;
wire net8320;
wire net1678;
wire net1236;
wire net3397;
wire net166;
wire net1621;
wire net6466;
wire net388;
wire net402;
wire net387;
wire net2924;
wire net1097;
wire net3565;
wire net4489;
wire net4243;
wire net1874;
wire net385;
wire in21;
wire net10671;
wire net10304;
wire net9818;
wire net5303;
wire net2825;
wire net384;
wire net2050;
wire net2456;
wire net885;
wire net2234;
wire net3639;
wire net2156;
wire net8655;
wire net207;
wire net317;
wire net7528;
wire net3273;
wire net1089;
wire net4610;
wire net5482;
wire net6548;
wire net10078;
wire net1666;
wire net4400;
wire net1277;
wire net2298;
wire net155;
wire net1087;
wire net2070;
wire net3858;
wire net3344;
wire net3568;
wire net5048;
wire net2934;
wire net1034;
wire in8;
wire net4370;
wire net4449;
wire net10361;
wire net4818;
wire net6296;
wire net759;
wire net10892;
wire net1518;
wire net2089;
wire net3399;
wire net5358;
wire net152;
wire net139;
wire net5987;
wire net895;
wire net1249;
wire net3651;
wire net742;
wire net8947;
wire net2759;
wire net2893;
wire net4689;
wire net9642;
wire net5682;
wire net2533;
wire net3680;
wire net2025;
wire net10834;
wire net132;
wire net7713;
wire net1221;
wire net862;
wire net131;
wire net6498;
wire net733;
wire net2673;
wire net129;
wire net2529;
wire net4453;
wire net5780;
wire net10513;
wire net7044;
wire net3418;
wire net633;
wire net318;
wire net2304;
wire net9486;
wire net8772;
wire net7029;
wire net810;
wire net6735;
wire net6853;
wire net6986;
wire net258;
wire net10207;
wire net2789;
wire net3115;
wire net5563;
wire net123;
wire net592;
wire net11352;
wire net7466;
wire net117;
wire net3973;
wire net9553;
wire net121;
wire net10721;
wire net5976;
wire net1297;
wire net0;
wire net3167;
wire net11262;
wire net4303;
wire net8985;
wire net1982;
wire net10130;
wire net3403;
wire net462;
wire net653;
wire net3682;
wire net5759;
wire net1617;
wire net4306;
wire net285;
wire net600;
wire net5877;
wire net1234;
wire net7821;
wire net2236;
wire net1043;
wire net8020;
wire net4579;
wire net2995;
wire net11004;
wire net9936;
wire net73;
wire net10947;
wire net4401;
wire net11329;
wire net825;
wire net4402;
wire net10019;
wire net1765;
wire net113;
wire net2550;
wire net6089;
wire net752;
wire net3290;
wire net1332;
wire net309;
wire net791;
wire net4218;
wire net7370;
wire net538;
wire net833;
wire net8592;
wire in13;
wire net10065;
wire net4239;
wire net311;
wire net362;
wire net1226;
wire net978;
wire net2712;
wire net110;
wire net949;
wire net886;
wire net8618;
wire net2374;
wire net890;
wire net4075;
wire net2709;
wire net6153;
wire net69;
wire net8502;
wire net793;
wire net2167;
wire net9779;
wire net846;
wire net1569;
wire net4041;
wire net10374;
wire net627;
wire net59;
wire net717;
wire net3443;
wire net874;
wire net11388;
wire net7622;
wire net695;
wire net7467;
wire net1658;
wire net5258;
wire net513;
wire net9946;
wire net6147;
wire net3372;
wire net3113;
wire net6652;
wire net463;
wire net751;
wire net1551;
wire net915;
wire net7145;
wire net103;
wire net5609;
wire net2848;
wire net44;
wire net11166;
wire net849;
wire net100;
wire net97;
wire net2964;
wire net4411;
wire net6095;
wire net1878;
wire net394;
wire net4866;
wire net4993;
wire net3311;
wire net8537;
wire net787;
wire net2819;
wire net239;
wire net10002;
wire net27;
wire net195;
wire net1929;
wire net657;
wire net3945;
wire net94;
wire net1185;
wire net8487;
wire net2067;
wire net6663;
wire in12;
wire net9402;
wire net409;
wire net482;
wire net264;
wire net209;
wire net4683;
wire net582;
wire net3332;
wire net2646;
wire net8694;
wire net6530;
wire net5379;
wire net971;
wire net6921;
wire net88;
wire net1900;
wire net4553;
wire net9403;
wire net3164;
wire net5893;
wire net5243;
wire net735;
wire net99;
wire net3505;
wire net925;
wire net9984;
wire net7880;
wire net5406;
wire net2485;
wire net826;
wire net3179;
wire net199;
wire net2318;
wire net458;
wire net6760;
wire net678;
wire net262;
wire net1287;
wire net4759;
wire net3633;
wire net3571;
wire net1789;
wire net5407;
wire net10852;
wire net87;
wire net11033;
wire net7177;
wire net5568;
wire net290;
wire net66;
wire net8963;
wire net5473;
wire net6737;
wire net5112;
wire net1710;
wire net486;
wire net9969;
wire net9012;
wire net7278;
wire net2357;
wire net1046;
wire net10550;
wire net6360;
wire net857;
wire net81;
wire net3298;
wire net9420;
wire net3420;
wire net2264;
wire net2514;
wire net7216;
wire net6596;
wire net9962;
wire net202;
wire net5040;
wire net2339;
wire net572;
wire net3795;
wire net7728;
wire net1212;
wire net1545;
wire net2428;
wire net11;
wire net3322;
wire net11330;
wire net1448;
wire in7;
wire net374;
wire net9296;
wire net4447;
wire net799;
wire net1486;
wire net1707;
wire net4162;
wire net11313;
wire net7982;
wire net6356;
wire net2074;
wire net2100;
wire net889;
wire net8835;
wire net877;
wire net490;
wire net1064;
wire net2647;
wire net8640;
wire net298;
wire net467;
wire net241;
wire net851;
wire net9;
wire net1028;
wire net6017;
wire net998;
wire net9943;
wire net3166;
wire net11223;
wire net4373;
wire net160;
wire net1223;
wire net765;
wire net2853;
wire net252;
wire net10101;
wire net8287;
wire net7470;
wire net1603;
wire net31;
wire net288;
wire net2200;
wire net441;
wire net673;
wire net1314;
wire net3402;
wire net2155;
wire net6957;
wire net3236;
wire net2283;
wire net3686;
wire net773;
wire net3391;
wire net4653;
wire net7092;
wire net3303;
wire in6;
wire net4619;
wire net167;
wire net1414;
wire net9712;
wire net2876;
wire net2750;
wire net2189;
wire net9255;
wire net7320;
wire net2330;
wire net891;
wire net5617;
wire net11562;
wire net11324;
wire net8221;
wire net3304;
wire net8422;
wire net6381;
wire net75;
wire net2053;
wire net2513;
wire net8308;
wire net523;
wire net9082;
wire net2983;
wire net45;
wire net5488;
wire net3171;
wire net4979;
wire net935;
wire net3468;
wire net5603;
wire net4;
wire net9110;
wire net334;
wire net2268;
wire net477;
wire net9844;
wire net1489;
wire net2522;
wire net481;
wire net11175;
wire net3299;
wire net6;
wire net8531;
wire net5913;
wire net665;
wire net2371;
wire net10863;
wire net9609;
wire net1788;
wire net9093;
wire net4362;
wire net5602;
wire net379;
wire net197;
wire net6612;
wire net11543;
wire net1387;
wire net10380;
wire net779;
wire net10467;
wire net3414;
wire net106;
wire net8896;
wire net6509;
wire net5350;
wire net995;
wire net7575;
wire net3876;
wire net2451;
wire net566;
wire net1210;
wire net1172;
wire net1498;
wire net7788;
wire net2621;
wire net1419;
wire net2670;
wire net68;
wire net6400;
wire net1405;
wire net7406;
wire net723;
wire net1177;
wire net6344;
wire net1110;
wire net696;
wire net4074;
wire net2008;
wire net8511;
wire net1632;
wire net7069;
wire net8177;
wire net7825;
wire net245;
wire net3192;
wire net1834;
wire net2839;
wire net2396;
wire net6079;
wire net3592;
wire net667;
wire net3452;
wire net18;
wire net1214;
wire net11568;
wire net7061;
wire net90;
wire net10165;
wire net5947;
wire net1425;
wire net8;
wire net8609;
wire net1677;
wire net1727;
wire net3460;
wire net2849;
wire net10867;
wire net2688;
wire net2804;
wire net2082;
wire net1443;
wire in23;
wire net3558;
wire net5866;
wire net7907;
wire net7630;
wire net4017;
wire net9646;
wire net9608;
wire net163;
wire net3170;
wire net7414;
wire net51;
wire net5680;
wire net10371;
wire net2034;
wire net5800;
wire net2285;
wire net726;
wire net1165;
wire net11009;
wire net5577;
wire net5748;
wire net7132;
wire net10496;
wire net7800;
wire net347;
wire net5090;
wire net1007;
wire net1408;
wire net6909;
wire net2526;
wire net9637;
wire net4910;
wire net84;
wire net2577;
wire net2667;
wire net6122;
wire net398;
wire net1610;
wire net2363;
wire net7966;
wire net6188;
wire net3128;
wire in4;
wire net3309;
wire net1971;
wire net9526;
wire net240;
wire net9379;
wire net4799;
wire net1885;
wire net175;
wire net682;
wire net570;
wire net1777;
wire net7805;
wire net274;
wire in16;
wire net1549;
wire net4497;
wire net5886;
wire net2308;
wire net1252;
wire net1503;
wire net1676;
wire net5216;
wire net2633;
wire net496;
wire net1055;
wire net426;
wire net8441;
wire net348;
wire net1668;
wire net962;
wire net10420;
wire net36;
wire net4441;
wire net507;
wire net5673;
wire net1338;
wire net2201;
wire net671;
wire net7381;
wire net7491;
wire net3383;
wire net8595;
wire net21;
wire net143;
wire net609;
wire net1421;
wire net920;
wire net6911;
wire net3450;
wire net625;
wire net393;
wire net522;
wire net2463;
wire net1745;
wire in20;
wire net491;
wire net10838;
wire net818;
wire net4988;
wire net300;
wire net157;
wire net2081;
wire net10336;
wire net1935;
wire net95;
wire net7596;
wire net79;
wire net835;
wire net20;
wire net4002;
wire net10079;
wire net86;
wire net601;
wire net2256;
wire net3361;
wire net1530;
wire net3983;
wire net154;
wire net1006;
wire net9930;
wire net4260;
wire net11492;
wire net6706;
wire net7658;
wire net1893;
wire net10991;
wire net251;
wire net1420;
wire net5449;
wire in18;
wire net6484;
wire net775;
wire net10989;
wire net10527;
wire net3364;
wire net254;
wire net7646;
wire net64;
wire net8013;
wire net408;
wire net4063;
wire net2530;
wire net2049;
wire net951;
wire net11507;
wire net12;
wire net11470;
wire net536;
wire net7897;
wire net83;
wire net33;
wire net11449;
wire net4167;
wire net11304;
wire net1011;
wire net9873;
wire net2150;
wire net185;
wire net5637;
wire net10347;
wire net4738;
wire net5792;
wire net3200;
wire net1820;
wire net10763;
wire net5699;
wire net638;
wire net10698;
wire net8755;
wire net128;
wire net5392;
wire net3176;
wire net2866;
wire net7818;
wire net2980;
wire net4326;
wire net1205;
wire net37;
wire net2384;
wire net7124;
wire net4184;
wire net530;
wire net9391;
wire net5117;
wire net6156;
wire net1511;
wire net38;
wire net3569;
wire net11119;
wire net3630;
wire net127;
wire net7257;
wire net1346;
wire net11283;
wire net2814;
wire net569;
wire net10707;
wire net502;
wire net158;
wire net6458;
wire net6724;
wire net3428;
wire net145;
wire net8194;
wire net213;
wire net5936;
wire net11584;
wire net7834;
wire net499;
wire net6278;
wire net50;
wire net2128;
wire net6069;
wire net2103;
wire net4945;
wire net7355;
wire net229;
wire net732;
wire net4869;
wire net457;
wire net645;
wire net4668;
wire net1636;
wire net11448;
wire net479;
wire net149;
wire net10316;
wire net57;
wire net6006;
wire net984;
wire net8126;
wire net3495;
wire net2838;
wire net3845;
wire net3172;
wire net9284;
wire net137;
wire net2203;
wire net3182;
wire net4960;
wire net7494;
wire net5024;
wire net5436;
wire net5481;
wire net11017;
wire net10809;
wire net9480;
wire net6303;
wire net1586;
wire net3843;
wire net1148;
wire net1168;
wire net10460;
wire net2346;
wire net380;
wire net11423;
wire net3197;
wire net359;
wire net993;
wire net191;
wire net755;
wire net47;
wire net5013;
wire net3625;
wire net10971;
wire net1104;
wire net5834;
wire net512;
wire net7282;
wire net3052;
wire net2415;
wire net8743;
wire net7074;
wire net1305;
wire net10760;
wire net13;
wire net3899;
wire net3001;
wire net3421;
wire net89;
wire net2942;
wire net741;
wire net3534;
wire net10063;
wire net3446;
wire net6818;
wire net944;
wire net11316;
wire net1714;
wire net5177;
wire net5267;
wire net9489;
wire net3465;
wire net6885;
wire net1213;
wire net1410;
wire net3188;
wire net395;
wire net6733;
wire net2992;
wire net2387;
wire net49;
wire net6702;
wire net7021;
wire net664;
wire net9866;
wire net7618;
wire net296;
wire net10171;
wire net855;
wire net55;
wire net134;
wire net3474;
wire net3585;
wire net1182;
wire net4054;
wire net5928;
wire net6941;
wire net6717;
wire net2212;
wire in1;
wire net74;
wire net4692;
wire net2077;
wire net11575;
wire net210;
wire net3254;
wire net4098;
wire net1954;
wire net4211;
wire net1237;
wire net10220;
wire net1317;
wire net9119;
wire net7331;
wire net5977;
wire net176;
wire net80;
wire net756;
wire net1970;
wire net10915;
wire net1858;
wire net9277;
wire net1243;
wire net1284;
wire net2857;
wire net5306;
wire net1639;
wire net852;
wire net3683;
wire net1465;
wire net6064;
wire net3642;
wire net445;
wire net7490;
wire net3785;
wire net5053;
wire net5661;
wire net9686;
wire net8617;
wire net70;
wire net2193;
wire net279;
wire net11173;
wire net3453;
wire net2;
wire net2468;
wire net192;
wire net594;
wire net174;
wire net6092;
wire net560;
wire net1755;
wire net225;
wire net1653;
wire net7705;
wire net265;
wire net6474;
wire net10948;
wire net9186;
wire net1804;
wire net2437;
wire net96;
wire net8230;
wire net3513;
wire net4939;
wire in2;
wire net610;
wire net180;
wire net4252;
wire net550;
wire net4520;
wire net3694;
wire net1542;
wire net3434;
wire net4153;
wire net5132;
wire net1447;
wire net9582;
wire net101;
wire net3784;
wire net3711;
wire net281;
wire net181;
wire net698;
wire net3510;
wire net1986;
wire net2278;
wire net182;
wire net3201;
wire net641;
wire net7604;
wire net6990;
wire net1033;
wire net10919;
wire net7613;
wire net785;
wire net701;
wire net286;
wire net5221;
wire net8742;
wire net2547;
wire net3139;
wire net476;
wire net3393;
wire net722;
wire net1095;
wire net4832;
wire net1803;
wire net301;
wire net1683;
wire net3315;
wire net8573;
wire net2427;
wire net345;
wire net3461;
wire net537;
wire net1881;
wire net10342;
wire net5373;
wire net8759;
wire net7429;
wire net2703;
wire net4460;
wire net966;
wire net4924;
wire net2333;
wire net1016;
wire net8099;
wire net193;
wire net1348;
wire net7042;
wire net48;
wire net8774;
wire net2627;
wire net194;
wire net3927;
wire net4337;
wire net5628;
wire net198;
wire net360;
wire net2833;
wire net2012;
wire net8841;
wire net6549;
wire net6881;
wire net236;
wire net9445;
wire net320;
wire net4304;
wire net295;
wire net204;
wire net3620;
wire net8824;
wire net3174;
wire net3613;
wire net7942;
wire net7692;
wire net3747;
wire net589;
wire net53;
wire net583;
wire net214;
wire net3665;
wire net9882;
wire net6994;
wire net7441;
wire net1262;
wire net10985;
wire net8010;
wire net767;
wire net3797;
wire net7147;
wire net237;
wire net4255;
wire net9848;
wire net480;
wire net5681;
wire net8282;
wire net1901;
wire net924;
wire net9127;
wire net2701;
wire net3898;
wire net3320;
wire net233;
wire net6744;
wire net8482;
wire net3718;
wire net220;
wire net6131;
wire net520;
wire net981;
wire net3892;
wire net7440;
wire net366;
wire net607;
wire net7080;
wire net651;
wire net7768;
wire net620;
wire net6997;
wire net939;
wire net3347;
wire net10454;
wire net4586;
wire net3773;
wire net5152;
wire net1614;
wire net2486;
wire net452;
wire net2372;
wire net2592;
wire net63;
wire net11305;
wire net2227;
wire net7139;
wire net10264;
wire net1371;
wire net613;
wire net6914;
wire net760;
wire net7303;
wire net223;
wire net5362;
wire net4996;
wire net897;
wire net908;
wire net438;
wire net10362;
wire net9134;
wire net2994;
wire net2678;
wire net10074;
wire net6517;
wire net8690;
wire net227;
wire net3611;
wire net9021;
wire net7346;
wire in9;
wire net660;
wire net6036;
wire net6414;
wire net542;
wire net2702;
wire net1326;
wire net628;
wire net2914;
wire net9184;
wire net5518;
wire net1748;
wire net526;
wire net1495;
wire net2573;
wire net4605;
wire net10309;
wire net230;
wire net10754;
wire net1492;
wire net3755;
wire net3297;
wire net5186;
wire net577;
wire net5095;
wire net661;
wire net1910;
wire net1467;
wire net10049;
wire net7469;
wire net10897;
wire net4773;
wire net3147;
wire net8167;
wire net2202;
wire net8398;
wire net5061;
wire net4774;
wire net418;
wire net323;
wire net11047;
wire net10245;
wire net552;
wire net2899;
wire net244;
wire net3701;
wire net7782;
wire net7219;
wire net2773;
wire net905;
wire net10686;
wire net338;
wire net672;
wire net3098;
wire net4273;
wire net2865;
wire net1790;
wire net24;
wire net1602;
wire net3640;
wire net801;
wire net2147;
wire net10773;
wire net5087;
wire net249;
wire net8436;
wire net7550;
wire net5218;
wire net8132;
wire net1593;
wire net9246;
wire net3417;
wire net5943;
wire net9619;
wire net6070;
wire net5696;
wire net2132;
wire net10134;
wire net9257;
wire net3915;
wire net5610;
wire net8859;
wire net3463;
wire net518;
wire net3848;
wire net10356;
wire net1499;
wire net2911;
wire net7792;
wire net3605;
wire net5952;
wire net6198;
wire net183;
wire net1434;
wire net272;
wire net1558;
wire net902;
wire net10612;
wire net200;
wire net635;
wire net8829;
wire net8243;
wire net5195;
wire net6256;
wire net3771;
wire net234;
wire net4545;
wire net598;
wire net1538;
wire net4130;
wire net4798;
wire net961;
wire net884;
wire net6277;
wire net487;
wire net6743;
wire net261;
wire net7515;
wire net1253;
wire net315;
wire net9775;
wire net1137;
wire net3441;
wire net1426;
wire net5586;
wire net7680;
wire net493;
wire net263;
wire net2221;
wire net4384;
wire net10059;
wire net8594;
wire net8359;
wire net112;
wire net3923;
wire net6094;
wire net1396;
wire net8906;
wire net2916;
wire net2477;
wire net4120;
wire net2654;
wire net2199;
wire net6423;
wire net5460;
wire net6647;
wire net8386;
wire net663;
wire net10598;
wire net1821;
wire net6421;
wire net11493;
wire net372;
wire net8277;
wire net2419;
wire net10156;
wire net7396;
wire net443;
wire net17;
wire net10590;
wire net270;
wire net8616;
wire net7820;
wire net3689;
wire net757;
wire net9635;
wire net1384;
wire net6951;
wire net997;
wire net7962;
wire net5309;
wire net3;
wire net2293;
wire net4636;
wire net727;
wire net10870;
wire net344;
wire net9259;
wire net6063;
wire net9380;
wire net3770;
wire net5906;
wire net9903;
wire net3475;
wire net4763;
wire net1643;
wire net2778;
wire net10973;
wire net5341;
wire net878;
wire net593;
wire net10907;
wire net278;
wire net7700;
wire net3685;
wire net1163;
wire in10;
wire net4961;
wire net436;
wire net10860;
wire net2140;
wire net3374;
wire net4930;
wire net11280;
wire net1001;
wire net4179;
wire net7084;
wire net2861;
wire net161;
wire net7544;
wire net5639;
wire net291;
wire net9098;
wire net5966;
wire net11162;
wire net9880;
wire net1595;
wire net1836;
wire net588;
wire net529;
wire net376;
wire net1359;
wire net10122;
wire net4317;
wire net370;
wire net3617;
wire net19;
wire net4884;
wire net5159;
wire net306;
wire net4944;
wire net1717;
wire net1778;
wire net8914;
wire net1026;
wire net10327;
wire net1009;
wire net446;
wire net141;
wire net9940;
wire net8909;
wire net7162;
wire net3009;
wire net1684;
wire net784;
wire net1696;
wire net7775;
wire net3245;
wire net10514;
wire net5108;
wire net1862;
wire net130;
wire net1204;
wire net4821;
wire net9658;
wire net932;
wire net7156;
wire net217;
wire net312;
wire net1018;
wire net332;
wire net1158;
wire net93;
wire net9949;
wire net5315;
wire net7;
wire net10;
wire net2327;
wire net9235;
wire net8734;
wire in22;
wire net11322;
wire net2935;
wire net7127;
wire net3007;
wire net2365;
wire net10891;
wire net4868;
wire net9317;
wire net3531;
wire net455;
wire net2855;
wire net423;
wire net958;
wire net3185;
wire net976;
wire net4633;
wire net8503;
wire net2289;
wire net72;
wire net3132;
wire net7858;
wire net221;
wire net11511;
wire net965;
wire net337;
wire net4568;
wire net968;
wire net7246;
wire net4507;
wire net7408;
wire net9318;
wire net3577;
wire net1452;
wire net5965;
wire net3676;
wire net2554;
wire net3667;
wire net3270;
wire net3573;
wire net1440;
wire net367;
wire net2821;
wire net597;
wire net3229;
wire net704;
wire net349;
wire net8399;
wire net2556;
wire net1200;
wire net2002;
wire net5497;
wire net9676;
wire net2552;
wire net2805;
wire net10624;
wire net4455;
wire net464;
wire net6712;
wire net1635;
wire net356;
wire net9177;
wire net2815;
wire net8463;
wire net2093;
wire net1823;
wire net9478;
wire net1693;
wire net8054;
wire net2764;
wire net4213;
wire net371;
wire net1756;
wire net11320;
wire net859;
wire net4750;
wire net6490;
wire net11130;
wire net4451;
wire net3969;
wire net373;
wire net7936;
wire net4202;
wire net800;
wire net9149;
wire net3628;
wire net2629;
wire net3913;
wire net807;
wire net811;
wire net8505;
wire net812;
wire net9722;
wire net5953;
wire net1059;
wire net813;
wire net5326;
wire net1588;
wire net275;
wire net6019;
wire net7361;
wire net5292;
wire net196;
wire net1925;
wire net3119;
wire net10121;
wire net4840;
wire net6580;
wire net816;
wire net6703;
wire net11546;
wire net8591;
wire net2473;
wire net1310;
wire net819;
wire net3745;
wire net822;
wire net1528;
wire net3238;
wire net824;
wire net3769;
wire net2639;
wire net1462;
wire net6441;
wire net2736;
wire net3435;
wire net6307;
wire net4696;
wire net831;
wire net3760;
wire net832;
wire net3856;
wire net7368;
wire net9926;
wire net7072;
wire net3702;
wire net2069;
wire in25;
wire net4542;
wire net102;
wire net5349;
wire net841;
wire net1369;
wire net843;
wire net844;
wire net10877;
wire net5536;
wire net2231;
wire net71;
wire net2235;
wire net11567;
wire net845;
wire net4330;
wire net7245;
wire net839;
wire net3356;
wire net894;
wire net1068;
wire net6237;
wire net1892;
wire net5882;
wire net1832;
wire net10995;
wire net368;
wire net1159;
wire net7031;
wire net1839;
wire net856;
wire net10097;
wire net3244;
wire net809;
wire net858;
wire net2728;
wire net1449;
wire net1021;
wire net4190;
wire net1736;
wire net860;
wire net972;
wire net10633;
wire net2813;
wire net863;
wire net5712;
wire net4737;
wire net3908;
wire net7967;
wire net2507;
wire net1482;
wire net3471;
wire net2062;
wire net866;
wire net868;
wire net10056;
wire net5279;
wire net2031;
wire net4500;
wire net1507;
wire net5525;
wire net869;
wire net5084;
wire net5399;
wire net6088;
wire net1450;
wire net6799;
wire net871;
wire net1968;
wire net1367;
wire net873;
wire net2698;
wire net5874;
wire net989;
wire net7260;
wire net2458;
wire net6832;
wire net3561;
wire net10119;
wire net4972;
wire net879;
wire net8770;
wire net3852;
wire net9327;
wire net5010;
wire net6861;
wire net3398;
wire net1401;
wire net1083;
wire net10739;
wire net259;
wire net1065;
wire net881;
wire net5335;
wire net2927;
wire net1930;
wire net1973;
wire net6948;
wire net887;
wire net656;
wire net5993;
wire net892;
wire net7872;
wire net4487;
wire net893;
wire net10344;
wire net7326;
wire net6149;
wire net898;
wire net6404;
wire net3266;
wire net6956;
wire net903;
wire net4521;
wire net2889;
wire net5283;
wire net1259;
wire net7798;
wire net3753;
wire net906;
wire net9824;
wire net378;
wire net4111;
wire net955;
wire net6170;
wire net910;
wire net8557;
wire net3432;
wire net1329;
wire net5019;
wire net911;
wire net2697;
wire net4309;
wire net11396;
wire net608;
wire net913;
wire net4855;
wire net2447;
wire net714;
wire net922;
wire net3873;
wire net2457;
wire net4973;
wire net2311;
wire net1207;
wire net10050;
wire net926;
wire net5864;
wire net7249;
wire net9365;
wire net616;
wire net1608;
wire net6566;
wire net584;
wire net7314;
wire net930;
wire net2131;
wire net5946;
wire net3089;
wire net5833;
wire net2323;
wire net933;
wire net2593;
wire net4933;
wire net10676;
wire net2294;
wire net4104;
wire net4124;
wire net5741;
wire net1509;
wire net4535;
wire net1298;
wire net936;
wire net788;
wire net3654;
wire net8416;
wire net1955;
wire net6145;
wire net8910;
wire net1339;
wire net4338;
wire net11240;
wire net938;
wire net940;
wire net3761;
wire net3813;
wire net7178;
wire net3405;
wire net3979;
wire net8790;
wire net1147;
wire net5633;
wire net9952;
wire net1093;
wire net941;
wire net1737;
wire net943;
wire net4220;
wire net1657;
wire net990;
wire net10765;
wire net7677;
wire net946;
wire net1980;
wire net3189;
wire net1907;
wire net6461;
wire net7896;
wire net1364;
wire net1191;
wire net1136;
wire net6214;
wire net8267;
wire net3093;
wire net948;
wire net614;
wire net5026;
wire net2414;
wire net6419;
wire net1969;
wire net8313;
wire net5403;
wire net1024;
wire net3226;
wire net4409;
wire net8041;
wire net953;
wire net3329;
wire net5784;
wire net954;
wire net2223;
wire net1183;
wire net959;
wire net248;
wire net6128;
wire net7901;
wire net4076;
wire net2609;
wire net5354;
wire net5814;
wire net170;
wire net1194;
wire net391;
wire net1407;
wire net11013;
wire net331;
wire net78;
wire net963;
wire net521;
wire net4931;
wire net5700;
wire net9913;
wire net1027;
wire net11155;
wire net8818;
wire net1816;
wire net1661;
wire net974;
wire net6288;
wire net5583;
wire net2004;
wire net979;
wire net980;
wire out16;
wire net1700;
wire net6723;
wire net4557;
wire net983;
wire net3282;
wire net8506;
wire net815;
wire net991;
wire net203;
wire net2267;
wire net1299;
wire net1928;
wire net6476;
wire net2856;
wire net1776;
wire net1000;
wire net3150;
wire net1003;
wire net466;
wire net2854;
wire net4139;
wire net789;
wire net1005;
wire net1008;
wire net3591;
wire net6654;
wire net2897;
wire net1427;
wire net8229;
wire net3604;
wire net8088;
wire net2662;
wire net1013;
wire net882;
wire net3343;
wire net11075;
wire net3208;
wire net10370;
wire net1629;
wire net416;
wire net4440;
wire net1023;
wire net2537;
wire net498;
wire net4856;
wire net1541;
wire net528;
wire net6203;
wire net1115;
wire net6766;
wire net10987;
wire net10205;
wire net2198;
wire net5411;
wire net1031;
wire net1694;
wire net2799;
wire net11024;
wire net4429;
wire net10982;
wire net1035;
wire net11243;
wire net7883;
wire net4482;
wire net5263;
wire net284;
wire net5660;
wire net1510;
wire net29;
wire net4527;
wire net606;
wire net4646;
wire net7957;
wire net1036;
wire net3263;
wire net4394;
wire net1871;
wire net9302;
wire net694;
wire net2770;
wire net1042;
wire net4513;
wire net9744;
wire net7345;
wire net9510;
wire net3703;
wire net567;
wire net1044;
wire net630;
wire net3048;
wire net7793;
wire net5668;
wire net1152;
wire net2895;
wire net5524;
wire net4010;
wire net2316;
wire net1045;
wire net2297;
wire net7637;
wire net1711;
wire net1400;
wire net5167;
wire net4267;
wire net1269;
wire net250;
wire net4990;
wire net2531;
wire net2613;
wire net5519;
wire net1048;
wire net6465;
wire net2755;
wire net1422;
wire net1879;
wire net10432;
wire net8420;
wire net1020;
wire net2492;
wire net1056;
wire net10314;
wire net2501;
wire net4425;
wire net5262;
wire net6697;
wire net6813;
wire net4601;
wire net5538;
wire net2454;
wire net5305;
wire net10434;
wire net602;
wire net1744;
wire net1062;
wire net9229;
wire net3751;
wire net10250;
wire net2614;
wire net1066;
wire net1067;
wire net6671;
wire net1071;
wire net42;
wire net5064;
wire net1072;
wire net4971;
wire net8967;
wire net8211;
wire net2780;
wire net1642;
wire net3231;
wire net9819;
wire net1622;
wire net2055;
wire net10626;
wire net1630;
wire net7563;
wire net1073;
wire net1227;
wire net1076;
wire net11385;
wire net1361;
wire net1150;
wire net9551;
wire net5038;
wire net2301;
wire net6455;
wire net11219;
wire net9730;
wire net6267;
wire net1868;
wire net1079;
wire net5272;
wire net2472;
wire net92;
wire net2809;
wire net3886;
wire net1500;
wire net3962;
wire net9643;
wire net6434;
wire net880;
wire net6764;
wire net5410;
wire net739;
wire net1081;
wire net386;
wire net5669;
wire net2757;
wire net1094;
wire net1323;
wire net7223;
wire net142;
wire net2011;
wire net5447;
wire net2612;
wire net389;
wire net7481;
wire net1098;
wire net9150;
wire net1406;
wire net273;
wire net1099;
wire net1493;
wire net1101;
wire net1103;
wire net10568;
wire net9814;
wire net7102;
wire net1105;
wire net3152;
wire net5284;
wire net2405;
wire net6684;
wire net8133;
wire net16;
wire net2206;
wire net2455;
wire net4515;
wire net1108;
wire net3835;
wire net9584;
wire net5229;
wire net1978;
wire net3768;
wire net3069;
wire net1634;
wire net1665;
wire net1039;
wire net9440;
wire net4026;
wire net3072;
wire net5963;
wire net1112;
wire net1119;
wire net314;
wire net1090;
wire net1120;
wire net1523;
wire net4023;
wire net1126;
wire net7192;
wire net3365;
wire net1818;
wire net1127;
wire net1712;
wire net10781;
wire net8440;
wire net1129;
wire net4336;
wire net5415;
wire net5455;
wire net1130;
wire net11138;
wire net1131;
wire net4742;
wire net5210;
wire net3065;
wire net684;
wire net1132;
wire out23;
wire net1589;
wire net7589;
wire net1133;
wire net8340;
wire net3292;
wire net7095;
wire net3054;
wire net2644;
wire net6872;
wire net6225;
wire net2564;
wire net5165;
wire net6980;
wire net619;
wire net1141;
wire net11381;
wire net2133;
wire net2594;
wire net4915;
wire net2488;
wire net5394;
wire out15;
wire net1144;
wire net4439;
wire net8767;
wire net1149;
wire net1077;
wire net456;
wire net7137;
wire net10917;
wire net392;
wire net6234;
wire net10560;
wire net1230;
wire net9121;
wire net1652;
wire net1411;
wire net3602;
wire net2121;
wire net8599;
wire net1160;
wire net4060;
wire net2795;
wire net2976;
wire net2937;
wire net9707;
wire net2320;
wire net1161;
wire net6677;
wire net11084;
wire net2715;
wire net2512;
wire net1164;
wire net1303;
wire net7239;
wire net2112;
wire net3499;
wire net1996;
wire net9101;
wire net6324;
wire net62;
wire net1171;
wire net2434;
wire net2540;
wire net5069;
wire net9521;
wire net3075;
wire net1174;
wire net6228;
wire net5421;
wire net201;
wire net9556;
wire net9092;
wire net1906;
wire net3566;
wire net2944;
wire net1180;
wire net5464;
wire net7319;
wire net2920;
wire net2139;
wire net2359;
wire net4908;
wire net3430;
wire net615;
wire net5820;
wire net10952;
wire net460;
wire net6877;
wire net1184;
wire net2867;
wire net2239;
wire net8590;
wire net1799;
wire net1186;
wire net9626;
wire net821;
wire net9792;
wire net2449;
wire net9388;
wire net34;
wire net5867;
wire net9442;
wire net358;
wire net1516;
wire net4110;
wire net6761;
wire net8817;
wire net1281;
wire net3603;
wire net9662;
wire net8310;
wire net76;
wire net3887;
wire net1199;
wire net1268;
wire net1311;
wire net1201;
wire net1202;
wire net10166;
wire net4551;
wire net7702;
wire net4609;
wire net9776;
wire net3424;
wire net8662;
wire net6876;
wire net1206;
wire net3044;
wire net2090;
wire net558;
wire net4671;
wire net668;
wire net3422;
wire net1578;
wire net11586;
wire net5838;
wire net1209;
wire net7328;
wire net9218;
wire net226;
wire net7638;
wire net1604;
wire net3138;
wire net1313;
wire net8698;
wire net1217;
wire net2403;
wire net4154;
wire net4313;
wire net120;
wire net2605;
wire net4493;
wire net1267;
wire net5645;
wire net2394;
wire net2099;
wire net1222;
wire net1491;
wire net1225;
wire net6591;
wire net1228;
wire net2369;
wire net2489;
wire net9921;
wire net2046;
wire net883;
wire net5483;
wire net964;
wire net5827;
wire net11101;
wire net1232;
wire net256;
wire net1238;
wire net6636;
wire net2803;
wire net3091;
wire net2376;
wire net8563;
wire net8056;
wire net1240;
wire net8228;
wire net888;
wire net747;
wire net3520;
wire net1244;
wire net9414;
wire net5271;
wire net1718;
wire net5166;
wire net5974;
wire net215;
wire net1245;
wire net3627;
wire net6431;
wire net7465;
wire net11019;
wire net3114;
wire net1248;
wire net2228;
wire net1251;
wire net4849;
wire net2794;
wire net3258;
wire net3104;
wire net1231;
wire net2868;
wire net140;
wire net1255;
wire net8674;
wire net2146;
wire net1162;
wire net3429;
wire net9049;
wire net1257;
wire net2991;
wire net4793;
wire net91;
wire net1990;
wire net67;
wire net11258;
wire net401;
wire net5257;
wire net3970;
wire net654;
wire net1276;
wire net1278;
wire net8943;
wire net909;
wire net3960;
wire out21;
wire net4231;
wire net9125;
wire net5037;
wire net6927;
wire net1279;
wire net1598;
wire net6526;
wire net5758;
wire net798;
wire net1280;
wire net5724;
wire net8298;
wire net1307;
wire net7681;
wire net5378;
wire net2885;
wire net468;
wire net6398;
wire net421;
wire net1480;
wire net636;
wire net10227;
wire net3092;
wire net1282;
wire net4068;
wire net11225;
wire net6221;
wire net6692;
wire net1283;
wire net5194;
wire net5400;
wire net9077;
wire net1357;
wire net1286;
wire net1288;
wire net7597;
wire net5774;
wire net11005;
wire net1289;
wire net3551;
wire net1292;
wire net6576;
wire net10627;
wire net2699;
wire net1296;
wire net1550;
wire net1911;
wire net10539;
wire net9062;
wire net4215;
wire net1301;
wire net1302;
wire net7353;
wire net688;
wire net1553;
wire net1471;
wire net4748;
wire net7158;
wire net1306;
wire net1585;
wire net8679;
wire net8184;
wire net4958;
wire net5277;
wire net10516;
wire net1316;
wire net2360;
wire net6774;
wire net440;
wire net7492;
wire net4133;
wire net1831;
wire net1522;
wire net1322;
wire net4230;
wire net2802;
wire net2558;
wire net5630;
wire net1327;
wire net5156;
wire net1398;
wire net3107;
wire net3790;
wire net1619;
wire net9117;
wire net1341;
wire net2406;
wire net1342;
wire net1350;
wire net1300;
wire net2464;
wire net5629;
wire net6148;
wire net1260;
wire net1351;
wire net10875;
wire net4470;
wire net1355;
wire net5887;
wire net1483;
wire net11497;
wire net8931;
wire net2958;
wire net4234;
wire net834;
wire net10262;
wire net5790;
wire net1360;
wire net3935;
wire net7463;
wire net2441;
wire net1627;
wire net1562;
wire net10040;
wire net3183;
wire net643;
wire net1319;
wire net7959;
wire net2169;
wire net1366;
wire net5057;
wire net2589;
wire net4462;
wire net952;
wire net3448;
wire net1580;
wire net6796;
wire net351;
wire net4452;
wire net8090;
wire net848;
wire net10723;
wire net7226;
wire net1375;
wire net9872;
wire net3464;
wire net3925;
wire net973;
wire net451;
wire net2734;
wire net7685;
wire net1378;
wire net1092;
wire net6882;
wire net8703;
wire net1380;
wire net7828;
wire net1381;
wire net4387;
wire net10426;
wire net6425;
wire net9614;
wire net1382;
wire net10025;
wire net1389;
wire net2880;
wire net1435;
wire net9829;
wire net2466;
wire net804;
wire net10680;
wire net3607;
wire net937;
wire net1385;
wire net1386;
wire net5539;
wire net1388;
wire net3045;
wire in15;
wire net711;
wire net1591;
wire net1784;
wire net7070;
wire net1391;
wire net2080;
wire net10203;
wire net2548;
wire net719;
wire net3572;
wire net1394;
wire net11426;
wire net1395;
wire net2721;
wire net6905;
wire net1962;
wire net1399;
wire net8928;
wire net931;
wire net381;
wire net429;
wire net1402;
wire net7015;
wire net1403;
wire net2213;
wire net2982;
wire net484;
wire net2075;
wire net4768;
wire net1085;
wire net1404;
wire net828;
wire net2450;
wire net1413;
wire net321;
wire net4081;
wire net2883;
wire net7450;
wire net2775;
wire net6337;
wire net8775;
wire net405;
wire net10391;
wire net10069;
wire net7504;
wire net1424;
wire net2423;
wire net1431;
wire net6565;
wire net6264;
wire net1944;
wire net1637;
wire net1432;
wire net2929;
wire net1600;
wire net3386;
wire net1433;
wire net1607;
wire net2250;
wire net1157;
wire net8801;
wire net1438;
wire net1441;
wire net5553;
wire net11134;
wire net9168;
wire net1344;
wire net1453;
wire net7101;
wire net7276;
wire net6472;
wire net697;
wire net4565;
wire net2999;
wire net433;
wire net6864;
wire net1333;
wire net1457;
wire net899;
wire net3537;
wire net1091;
wire net5837;
wire net1454;
wire net10577;
wire net7506;
wire net5360;
wire net1455;
wire net2254;
wire net2641;
wire net1844;
wire net2065;
wire net7475;
wire net3050;
wire net1456;
wire net1458;
wire net2844;
wire net7295;
wire net576;
wire net3043;
wire net10195;
wire net1626;
wire net6971;
wire net2683;
wire net1143;
wire net6038;
wire net6682;
wire net1461;
wire net1579;
wire net3563;
wire net1353;
wire net6229;
wire net1469;
wire net1169;
wire net1084;
wire net7262;
wire net4622;
wire net5027;
wire net5778;
wire net6068;
wire net1470;
wire net3518;
wire net6637;
wire net929;
wire net1473;
wire net447;
wire net1189;
wire net1478;
wire net5009;
wire net7022;
wire net2175;
wire net1271;
wire net5779;
wire net10390;
wire net3154;
wire net1484;
wire net6186;
wire net6975;
wire net7650;
wire net803;
wire net4015;
wire net3144;
wire net3644;
wire net3255;
wire net3019;
wire net1494;
wire net4079;
wire net5062;
wire net1496;
wire net5688;
wire net2966;
wire net9037;
wire net1497;
wire net6114;
wire net7204;
wire net3013;
wire net3181;
wire net1950;
wire net1504;
wire net10191;
wire net8596;
wire net3524;
wire net1670;
wire net4393;
wire net829;
wire net10192;
wire net1506;
wire net6573;
wire net8278;
wire net8268;
wire net14;
wire net8384;
wire net5695;
wire net1512;
wire net10688;
wire net5289;
wire net669;
wire net1513;
wire net10463;
wire net1514;
wire net10003;
wire net3549;
wire net1648;
wire net316;
wire net8481;
wire net1618;
wire net2562;
wire net7338;
wire net1916;
wire net1760;
wire net7418;
wire net8716;
wire net8200;
wire net1524;
wire net11018;
wire net1833;
wire net709;
wire in14;
wire net9981;
wire net3984;
wire net6730;
wire net8866;
wire net2671;
wire net375;
wire net5647;
wire net1485;
wire net1531;
wire net6607;
wire net1533;
wire net10014;
wire net1536;
wire net3490;
wire net10103;
wire net1584;
wire net5549;
wire net1735;
wire net5614;
wire net122;
wire net1547;
wire net9264;
wire net2178;
wire net1798;
wire net5058;
wire net1548;
wire net3954;
wire net7011;
wire net6924;
wire net115;
wire net7457;
wire net1554;
wire net8108;
wire net6645;
wire net778;
wire net557;
wire net190;
wire net5599;
wire net1557;
wire net3479;
wire net1559;
wire net677;
wire net1570;
wire net1746;
wire net837;
wire net3793;
wire net11482;
wire net11419;
wire net4847;
wire net5776;
wire net7016;
wire net77;
wire net1843;
wire net956;
wire net796;
wire net6973;
wire net7159;
wire net4035;
wire net4374;
wire net1564;
wire net11290;
wire net4072;
wire net2882;
wire net7635;
wire net2549;
wire net8748;
wire net1565;
wire net2116;
wire net3988;
wire net125;
wire net1926;
wire net1574;
wire net10774;
wire net1576;
wire net2919;
wire net8064;
wire net4413;
wire net1577;
wire net3283;
wire net1581;
wire net5264;
wire net4039;
wire net1587;
wire net8352;
wire net2087;
wire net1963;
wire net1920;
wire net6989;
wire net1594;
wire net3457;
wire net8204;
wire net7235;
wire net7241;
wire net1285;
wire net1078;
wire net242;
wire net2141;
wire net7082;
wire net9770;
wire net1606;
wire net1924;
wire net7046;
wire net1609;
wire net2523;
wire net308;
wire net2266;
wire net4901;
wire net1167;
wire net2669;
wire net7103;
wire net3805;
wire net2785;
wire net942;
wire net5727;
wire net1572;
wire net7555;
wire net1304;
wire net1620;
wire net257;
wire net1852;
wire net5555;
wire net3415;
wire net9986;
wire net1623;
wire net2355;
wire net1124;
wire net7185;
wire net1697;
wire net3108;
wire net1633;
wire net4148;
wire net8192;
wire net3106;
wire net5579;
wire net5371;
wire net11564;
wire net8582;
wire net618;
wire net2690;
wire net1641;
wire net527;
wire net1644;
wire net1646;
wire net1651;
wire net1650;
wire net4710;
wire net2909;
wire net2028;
wire net5440;
wire net4181;
wire net3117;
wire net4620;
wire net1490;
wire net4589;
wire net205;
wire net4058;
wire net4185;
wire net2774;
wire net1479;
wire net6351;
wire net867;
wire net1904;
wire net7945;
wire net1669;
wire net623;
wire net11271;
wire net4200;
wire net10653;
wire net10534;
wire net1671;
wire net8289;
wire net2686;
wire net2217;
wire net1672;
wire net3358;
wire net921;
wire net6483;
wire net712;
wire net1674;
wire net2824;
wire net3040;
wire net1682;
wire net108;
wire net3196;
wire net7296;
wire net7963;
wire net3241;
wire net9301;
wire net271;
wire net5242;
wire net5746;
wire net1685;
wire net3041;
wire net3933;
wire net1751;
wire net1703;
wire net1686;
wire net10429;
wire net10159;
wire net782;
wire net1690;
wire net52;
wire net1692;
wire net2092;
wire net6640;
wire net1698;
wire net439;
wire net5000;
wire net5950;
wire net605;
wire out3;
wire net2484;
wire net10331;
wire net3296;
wire net6965;
wire net1706;
wire net6039;
wire net7952;
wire net1709;
wire net692;
wire net6385;
wire net3713;
wire net7979;
wire net3716;
wire net4352;
wire net4398;
wire net1667;
wire net3717;
wire net3259;
wire net3719;
wire net1246;
wire net5799;
wire net3720;
wire net543;
wire net3722;
wire net1599;
wire net3772;
wire net9031;
wire net4657;
wire net1247;
wire net5494;
wire net982;
wire net7423;
wire net4796;
wire net3723;
wire net5843;
wire net3725;
wire net5002;
wire net3727;
wire net11400;
wire net3728;
wire net6862;
wire net3730;
wire net10054;
wire net9172;
wire net3731;
wire net5967;
wire net3732;
wire net3734;
wire net11447;
wire net10794;
wire net9042;
wire net3735;
wire net2432;
wire net4071;
wire net2127;
wire net3736;
wire net9254;
wire net3739;
wire net11486;
wire net8315;
wire net4087;
wire net8813;
wire net5849;
wire net8031;
wire net1866;
wire net5656;
wire net3740;
wire net3741;
wire net9864;
wire net9070;
wire net9009;
wire net1758;
wire net3743;
wire net9827;
wire net3744;
wire net3222;
wire net260;
wire net3748;
wire net7774;
wire net6023;
wire net3749;
wire net4163;
wire net1356;
wire net3754;
wire net3756;
wire net6639;
wire net1616;
wire net7130;
wire net3757;
wire net3758;
wire net3715;
wire net7458;
wire net1187;
wire net3759;
wire net3763;
wire net3764;
wire net8499;
wire net8446;
wire net3766;
wire net10466;
wire net6661;
wire net3767;
wire net3774;
wire net10694;
wire net4178;
wire net3776;
wire net5208;
wire net7120;
wire net5782;
wire net1444;
wire net6655;
wire net3779;
wire net3918;
wire net2336;
wire net3780;
wire net3783;
wire net3786;
wire net8483;
wire net1242;
wire net3787;
wire net3928;
wire net3788;
wire net3789;
wire net3265;
wire net1211;
wire net4874;
wire net6048;
wire net8214;
wire net4014;
wire net6449;
wire net4736;
wire net7576;
wire net3301;
wire net3796;
wire net5173;
wire net4735;
wire net2328;
wire net7142;
wire net3798;
wire net3799;
wire net3800;
wire net3801;
wire net3807;
wire net9977;
wire net6492;
wire net3809;
wire net4665;
wire net1086;
wire net3810;
wire net7347;
wire net3812;
wire net5376;
wire net3814;
wire net6329;
wire net10766;
wire net3433;
wire net3817;
wire net7000;
wire net3818;
wire net3819;
wire net6335;
wire net3820;
wire net3821;
wire net10531;
wire net3822;
wire net8233;
wire net3826;
wire net5092;
wire net3827;
wire net10111;
wire net9762;
wire net4103;
wire net3828;
wire net7766;
wire net3829;
wire net3846;
wire net3830;
wire net6473;
wire net3833;
wire net2907;
wire net6026;
wire net3834;
wire net10659;
wire net3837;
wire net2986;
wire net6387;
wire net3653;
wire net3839;
wire net3840;
wire net3841;
wire net4782;
wire net5613;
wire net3842;
wire net716;
wire net3844;
wire net7817;
wire net3847;
wire net3824;
wire net4951;
wire net2713;
wire net3849;
wire net40;
wire net6172;
wire net3851;
wire net11121;
wire net3853;
wire net3854;
wire net9441;
wire net4408;
wire net3855;
wire net3857;
wire net3861;
wire net3862;
wire net3864;
wire net9531;
wire net3866;
wire net7778;
wire net4510;
wire net3867;
wire net3868;
wire net3869;
wire net9433;
wire net3870;
wire net5140;
wire net3871;
wire net11431;
wire net4967;
wire net11489;
wire net1195;
wire net6142;
wire net3872;
wire net3874;
wire net5704;
wire net4161;
wire net3437;
wire net3875;
wire net8548;
wire net2922;
wire net1783;
wire net3877;
wire net7940;
wire net3878;
wire net10501;
wire net3879;
wire net3880;
wire net5158;
wire net10057;
wire net7808;
wire net3598;
wire net3882;
wire net1053;
wire net3888;
wire net10682;
wire net3629;
wire net3889;
wire net3891;
wire net3893;
wire net8098;
wire net465;
wire net1860;
wire net3894;
wire net3895;
wire net9297;
wire net8664;
wire net2418;
wire net3902;
wire net7444;
wire net3555;
wire net3903;
wire net3904;
wire net11020;
wire net7987;
wire net3905;
wire net5080;
wire net3906;
wire net9808;
wire net4016;
wire net3907;
wire net5530;
wire net3909;
wire net4811;
wire net8375;
wire net7773;
wire net3910;
wire net3911;
wire net5649;
wire net3912;
wire net3916;
wire net4733;
wire net6124;
wire net5456;
wire net5496;
wire net6298;
wire net6578;
wire net9219;
wire net3917;
wire net7071;
wire net3919;
wire net3272;
wire net3922;
wire net5664;
wire net6731;
wire net3924;
wire net11153;
wire net1354;
wire net3926;
wire net3929;
wire net8804;
wire net3931;
wire net1216;
wire net1750;
wire net1753;
wire net3932;
wire net1532;
wire net6073;
wire net3934;
wire net3936;
wire net5578;
wire net8604;
wire net3937;
wire net9447;
wire net3664;
wire net3938;
wire net3940;
wire net900;
wire net3941;
wire net10112;
wire net1193;
wire net4764;
wire net3943;
wire net3946;
wire net3947;
wire net3948;
wire net3951;
wire net3952;
wire net3953;
wire net3956;
wire net3957;
wire net9477;
wire net3959;
wire net3963;
wire net6043;
wire net3966;
wire net5412;
wire net6787;
wire net3968;
wire net5007;
wire net3971;
wire net419;
wire net3974;
wire net9196;
wire net3975;
wire net4235;
wire net6046;
wire net3978;
wire net1515;
wire net4186;
wire net9345;
wire net5622;
wire net3981;
wire net10536;
wire net3982;
wire net1936;
wire net3985;
wire net3986;
wire net3991;
wire net3992;
wire net7170;
wire net11081;
wire net2282;
wire net3993;
wire net3994;
wire net6120;
wire net3996;
wire net3997;
wire net6358;
wire net3998;
wire net7947;
wire net3706;
wire net4089;
wire net3999;
wire net8089;
wire net2828;
wire net4003;
wire net2490;
wire net6403;
wire net4109;
wire net5126;
wire net4005;
wire net6630;
wire net10695;
wire net4007;
wire net4008;
wire net9754;
wire net8376;
wire net4012;
wire net46;
wire net4018;
wire net6543;
wire net4020;
wire net7435;
wire net4021;
wire net4926;
wire net4022;
wire net5900;
wire net1135;
wire net4024;
wire net11200;
wire net4580;
wire net6072;
wire net11071;
wire net8061;
wire net4027;
wire net6510;
wire net539;
wire net5386;
wire net7047;
wire net4028;
wire net4030;
wire net4031;
wire net4033;
wire net4036;
wire net4037;
wire net4820;
wire net6998;
wire net4038;
wire net4040;
wire net4042;
wire net666;
wire net4043;
wire net4276;
wire net4045;
wire net1917;
wire net5743;
wire net9354;
wire net5164;
wire net994;
wire net4046;
wire net4049;
wire net9549;
wire net8630;
wire net7611;
wire net4051;
wire net4052;
wire net6427;
wire net4053;
wire net4055;
wire net8562;
wire net4057;
wire net4059;
wire net10807;
wire net10788;
wire net8687;
wire net6422;
wire net658;
wire net5503;
wire net4061;
wire net4062;
wire net10777;
wire net5685;
wire net7065;
wire net4064;
wire net4084;
wire net8872;
wire net790;
wire net4065;
wire net6176;
wire net7839;
wire net6634;
wire net4066;
wire net565;
wire net4067;
wire net4069;
wire net8334;
wire net2310;
wire net4070;
wire net6541;
wire net4073;
wire net4680;
wire net6322;
wire net4077;
wire net7664;
wire net907;
wire net150;
wire net4078;
wire net4080;
wire net4082;
wire net9566;
wire net4083;
wire net10581;
wire net8162;
wire net2623;
wire net4090;
wire net5299;
wire net4091;
wire net10106;
wire net9072;
wire net4719;
wire net4093;
wire net5948;
wire net4095;
wire out24;
wire net4728;
wire net4101;
wire net8008;
wire net4434;
wire net5227;
wire net6448;
wire net5991;
wire net6763;
wire net5088;
wire net10674;
wire net4105;
wire net1423;
wire net4106;
wire net10654;
wire net4112;
wire net4114;
wire net7230;
wire net4117;
wire net3724;
wire net4119;
wire net4123;
wire net3425;
wire net5469;
wire net5321;
wire net6866;
wire net2358;
wire net4125;
wire net4126;
wire net4127;
wire net10113;
wire net5769;
wire net4129;
wire net4131;
wire net9562;
wire net4132;
wire net4136;
wire net3038;
wire net4140;
wire net7838;
wire net2465;
wire net4141;
wire net4142;
wire net82;
wire net4144;
wire net11370;
wire net8533;
wire net1134;
wire net4145;
wire net4146;
wire net4147;
wire net1235;
wire net5116;
wire net2984;
wire net4150;
wire net8059;
wire net4152;
wire net7951;
wire net2786;
wire net5389;
wire net410;
wire net4155;
wire net11332;
wire net449;
wire net7344;
wire net4160;
wire net4164;
wire net3087;
wire net4165;
wire net1142;
wire net4168;
wire net3156;
wire net4169;
wire net1417;
wire net2185;
wire net4171;
wire net5230;
wire net4173;
wire net4177;
wire net2511;
wire net4182;
wire net7831;
wire net6506;
wire net10172;
wire net148;
wire net4183;
wire net4187;
wire net5074;
wire net4189;
wire net6649;
wire net9271;
wire net5071;
wire net4192;
wire net3901;
wire net6993;
wire net4193;
wire net497;
wire net4194;
wire net8116;
wire net6255;
wire net7270;
wire net4197;
wire net2027;
wire net4198;
wire net9998;
wire net4199;
wire net10137;
wire net4265;
wire net8424;
wire net6310;
wire net4203;
wire net4205;
wire net4207;
wire net4208;
wire net1701;
wire net4209;
wire net3564;
wire net5302;
wire net5423;
wire net2768;
wire net4212;
wire net4217;
wire net4221;
wire net3328;
wire net4222;
wire net4648;
wire net235;
wire net5990;
wire net4223;
wire net8094;
wire net4224;
wire net917;
wire net4226;
wire net4227;
wire net10813;
wire net4228;
wire net4232;
wire net11000;
wire net4233;
wire net5207;
wire net3729;
wire net4237;
wire net4240;
wire net4241;
wire net2218;
wire net7189;
wire net11129;
wire net4245;
wire net6204;
wire net9656;
wire net4246;
wire net2965;
wire net5198;
wire net4247;
wire net6125;
wire net4248;
wire net6416;
wire net4249;
wire net4251;
wire net6488;
wire net4253;
wire net8657;
wire net4256;
wire net1628;
wire net4258;
wire net6785;
wire net9950;
wire net4259;
wire net5345;
wire net7104;
wire net4262;
wire net8000;
wire net1439;
wire net4263;
wire net3178;
wire net4269;
wire net1566;
wire net4264;
wire net4268;
wire net5434;
wire net4274;
wire net5135;
wire net3243;
wire net342;
wire net4275;
wire net2624;
wire net4278;
wire net54;
wire net4279;
wire net4281;
wire net11179;
wire net4631;
wire net11487;
wire net4283;
wire net11414;
wire net9308;
wire net9262;
wire net4284;
wire net4285;
wire net4286;
wire net4588;
wire net4612;
wire net3319;
wire net4288;
wire net2177;
wire net4289;
wire net4291;
wire net4292;
wire net4294;
wire net4295;
wire net4297;
wire net8135;
wire net4298;
wire net11022;
wire net4299;
wire net7079;
wire net4300;
wire net8065;
wire net2587;
wire net4302;
wire net2632;
wire net4826;
wire net1416;
wire net4305;
wire net2024;
wire net5944;
wire net7115;
wire net4311;
wire net6991;
wire net10799;
wire net7608;
wire net4314;
wire net8933;
wire net8019;
wire net4491;
wire net4318;
wire net4325;
wire net4625;
wire net4328;
wire net6252;
wire net4331;
wire net7384;
wire net10960;
wire net10251;
wire net519;
wire net4157;
wire net4332;
wire net4836;
wire net7256;
wire net4333;
wire net4334;
wire net4335;
wire net6361;
wire net8393;
wire net4339;
wire net7390;
wire net10243;
wire net4340;
wire net3335;
wire net4341;
wire net8141;
wire net5502;
wire net4342;
wire net8797;
wire net4188;
wire net4343;
wire net4970;
wire net4344;
wire net4345;
wire net2322;
wire net5401;
wire net2321;
wire net5049;
wire net10478;
wire net9698;
wire net4349;
wire net4350;
wire net5060;
wire net10876;
wire net4351;
wire net7329;
wire net8085;
wire net6504;
wire net4356;
wire net4357;
wire net4358;
wire net2717;
wire net4359;
wire net6894;
wire net5086;
wire net4360;
wire net10554;
wire net7722;
wire net6151;
wire net10462;
wire net4361;
wire net118;
wire net4364;
wire net1121;
wire net4367;
wire net4368;
wire net4369;
wire net4371;
wire net8451;
wire net517;
wire net4375;
wire net7495;
wire net7126;
wire net4376;
wire net6380;
wire net6849;
wire net4377;
wire net1082;
wire net6376;
wire in19;
wire net4379;
wire net4380;
wire net7190;
wire net4381;
wire net7639;
wire net1845;
wire net5429;
wire net4382;
wire net4383;
wire net10881;
wire net302;
wire net1740;
wire net4385;
wire net10217;
wire net4000;
wire net4386;
wire net1762;
wire net1679;
wire net4261;
wire net4388;
wire net7815;
wire net5114;
wire net6629;
wire net4392;
wire net4395;
wire net4396;
wire net10512;
wire net4853;
wire net4397;
wire net11558;
wire net5100;
wire net5255;
wire net10562;
wire net8171;
wire net4399;
wire net4403;
wire net10628;
wire net3897;
wire net6299;
wire net2945;
wire in11;
wire net4405;
wire net4410;
wire net10966;
wire net4412;
wire net6539;
wire net4416;
wire net4417;
wire net4418;
wire net4419;
wire net9838;
wire net8285;
wire net6481;
wire net8846;
wire net4421;
wire net2314;
wire net6268;
wire net4423;
wire net4426;
wire net4427;
wire net6436;
wire net4428;
wire net7111;
wire net188;
wire net5529;
wire net4433;
wire net9370;
wire net4436;
wire net10199;
wire net4667;
wire net339;
wire net6821;
wire net4438;
wire net4957;
wire net4442;
wire net369;
wire net2445;
wire net4445;
wire net6758;
wire net4446;
wire net5597;
wire net434;
wire net4448;
wire net4450;
wire net7854;
wire net5388;
wire net6585;
wire net4458;
wire net3482;
wire net4461;
wire net2303;
wire net5589;
wire net1655;
wire net424;
wire net4463;
wire net4464;
wire net7837;
wire net4466;
wire net4467;
wire net4469;
wire net1801;
wire net4471;
wire net10642;
wire net10605;
wire net4293;
wire net2136;
wire net5912;
wire net1254;
wire net4474;
wire net4476;
wire net4477;
wire net1691;
wire net4478;
wire net4479;
wire net5021;
wire net4481;
wire net5498;
wire net4484;
wire net7430;
wire net4485;
wire net4486;
wire net4490;
wire net5377;
wire net8237;
wire net4492;
wire net6179;
wire net4494;
wire net4496;
wire net173;
wire net4501;
wire net4503;
wire net4637;
wire net3594;
wire net4504;
wire net7382;
wire net4505;
wire net10346;
wire net675;
wire net4506;
wire net5381;
wire net4508;
wire net2551;
wire net5625;
wire net622;
wire net4509;
wire net2947;
wire net4511;
wire net6366;
wire net5926;
wire net4516;
wire net7599;
wire net4522;
wire net4523;
wire net4524;
wire net4525;
wire net8173;
wire net8115;
wire net4526;
wire net2153;
wire net4530;
wire net2306;
wire net4531;
wire net4534;
wire net11167;
wire net268;
wire net1534;
wire net5428;
wire net4536;
wire net5347;
wire net4539;
wire net5573;
wire net1487;
wire net4540;
wire net4541;
wire net4543;
wire net5420;
wire net469;
wire net4546;
wire net10702;
wire net6560;
wire net4722;
wire net7023;
wire net7332;
wire net4547;
wire net4549;
wire net4550;
wire net4552;
wire net4554;
wire net435;
wire net4555;
wire net5711;
wire net7081;
wire net9599;
wire net4556;
wire net4558;
wire net10077;
wire net508;
wire net4559;
wire net4562;
wire net187;
wire net6668;
wire net4567;
wire net7330;
wire net4569;
wire net11369;
wire net6642;
wire net2835;
wire net3206;
wire net4571;
wire net4287;
wire net4572;
wire net4590;
wire net4574;
wire net4575;
wire net10939;
wire net7741;
wire net3373;
wire net4576;
wire net4578;
wire net2095;
wire net6916;
wire net1358;
wire net7321;
wire net4581;
wire net5319;
wire net4583;
wire net6245;
wire net9944;
wire net4585;
wire net3823;
wire net4659;
wire net1590;
wire net4587;
wire net3580;
wire net4592;
wire net5728;
wire net1476;
wire net4593;
wire net4594;
wire net4596;
wire net7735;
wire net6534;
wire net4597;
wire net4598;
wire net7356;
wire net4599;
wire net3976;
wire net4600;
wire net4602;
wire net7048;
wire net4604;
wire net11052;
wire net5322;
wire net6669;
wire net9886;
wire net2676;
wire net4606;
wire net6958;
wire net30;
wire net4611;
wire net4731;
wire net1890;
wire net4613;
wire net6370;
wire net3781;
wire net4614;
wire net4615;
wire net3709;
wire net4616;
wire net4617;
wire net6732;
wire net10542;
wire net4621;
wire net4626;
wire in0;
wire net6919;
wire net3151;
wire net4627;
wire net6001;
wire net2926;
wire net3777;
wire net6932;
wire net3671;
wire net4628;
wire net1363;
wire net4629;
wire net3645;
wire net4630;
wire net4632;
wire net6084;
wire net4634;
wire net4635;
wire net2417;
wire net4050;
wire net4638;
wire net8045;
wire net4838;
wire net4640;
wire net6930;
wire net4641;
wire net4643;
wire net5043;
wire net1808;
wire net6949;
wire net8586;
wire net6572;
wire net4651;
wire net4654;
wire net4655;
wire net9372;
wire net7964;
wire net4656;
wire net5752;
wire net4660;
wire net8182;
wire net4752;
wire net4661;
wire net7419;
wire net4662;
wire net8181;
wire net4663;
wire net4664;
wire net4669;
wire net6152;
wire net4670;
wire net8072;
wire net222;
wire net4672;
wire net4674;
wire net404;
wire out1;
wire net2797;
wire net4675;
wire net4676;
wire net1915;
wire net4677;
wire net4678;
wire net4679;
wire net1274;
wire net4682;
wire net2288;
wire net4686;
wire net4687;
wire net8676;
wire net4688;
wire net4690;
wire net4691;
wire net4755;
wire net8709;
wire net2990;
wire net4693;
wire net4694;
wire net9348;
wire net3700;
wire net4644;
wire net4695;
wire net9468;
wire net4697;
wire net4698;
wire net9340;
wire net4699;
wire net4701;
wire net7827;
wire net4702;
wire net11357;
wire net4703;
wire net7273;
wire net6987;
wire net4705;
wire net992;
wire net4707;
wire net8500;
wire net4711;
wire net4366;
wire net5355;
wire net4712;
wire net4713;
wire net6320;
wire net4714;
wire net1088;
wire net218;
wire net4715;
wire net4257;
wire net4716;
wire net4717;
wire net3264;
wire net5742;
wire net4720;
wire net8807;
wire net2751;
wire net4999;
wire net4721;
wire net7720;
wire net4048;
wire net6839;
wire net5161;
wire net4723;
wire net4724;
wire net4725;
wire net4726;
wire net4727;
wire net7676;
wire net4729;
wire net4730;
wire net3990;
wire net6978;
wire net4732;
wire net4734;
wire net7237;
wire net4739;
wire net4740;
wire net4743;
wire net1933;
wire net2850;
wire net4102;
wire net4744;
wire net4746;
wire net4882;
wire net4166;
wire net4749;
wire net4751;
wire net2998;
wire net4753;
wire net4758;
wire net6067;
wire net4835;
wire net4760;
wire net2606;
wire net4761;
wire net4355;
wire net6393;
wire net4762;
wire net9964;
wire net4765;
wire net10805;
wire net9198;
wire net5598;
wire net4767;
wire net1117;
wire net4769;
wire net743;
wire net4770;
wire net6936;
wire net5190;
wire net4771;
wire net4772;
wire net4404;
wire net4432;
wire net6470;
wire net4009;
wire net4776;
wire net4777;
wire net10029;
wire net7995;
wire net7094;
wire net7718;
wire net4778;
wire net4271;
wire net6410;
wire net1106;
wire net4780;
wire net9627;
wire net4783;
wire net4784;
wire net4785;
wire net4430;
wire net4786;
wire net4788;
wire net4791;
wire net4792;
wire net11253;
wire net2366;
wire net1543;
wire net4795;
wire net4797;
wire net289;
wire net4800;
wire net2808;
wire net4801;
wire net4805;
wire net4324;
wire net7028;
wire net4806;
wire net4807;
wire net2771;
wire net6437;
wire net740;
wire net4809;
wire net11364;
wire net6482;
wire net10354;
wire net470;
wire net4810;
wire net4814;
wire net4816;
wire net4822;
wire net5564;
wire net4823;
wire net10849;
wire net4824;
wire net4519;
wire net4825;
wire net4827;
wire net11430;
wire net4829;
wire net6016;
wire net4830;
wire net9223;
wire net6438;
wire net4831;
wire net2367;
wire net4834;
wire net6417;
wire net4837;
wire net10115;
wire net4845;
wire net5287;
wire net3161;
wire net5986;
wire net6432;
wire net3690;
wire net4214;
wire net4848;
wire net4850;
wire net4851;
wire net4548;
wire net5384;
wire net8847;
wire net4857;
wire net4858;
wire net4860;
wire net4861;
wire net4862;
wire net1517;
wire net4864;
wire net4865;
wire net4867;
wire net509;
wire net4870;
wire net4871;
wire net8415;
wire net4872;
wire net1521;
wire net5129;
wire net9540;
wire net1932;
wire net4817;
wire net4875;
wire net5182;
wire net6699;
wire net4876;
wire net10157;
wire net4877;
wire net4879;
wire net4880;
wire net9920;
wire net4883;
wire net720;
wire net4885;
wire net10708;
wire net4886;
wire net4887;
wire net9532;
wire net4888;
wire net7461;
wire net4889;
wire net7941;
wire net4891;
wire net8333;
wire net4892;
wire net9201;
wire net5730;
wire net6059;
wire net8431;
wire net4894;
wire net4895;
wire net4897;
wire net4092;
wire net4898;
wire net6345;
wire net4900;
wire net2433;
wire net4903;
wire net3205;
wire net4905;
wire net4906;
wire net5635;
wire net4909;
wire net10890;
wire net6191;
wire net1675;
wire net5118;
wire net5154;
wire net6915;
wire net4912;
wire net11561;
wire net7060;
wire net4914;
wire net7388;
wire net4916;
wire net184;
wire net4918;
wire net6687;
wire net4919;
wire net7888;
wire net4277;
wire net5485;
wire net9939;
wire net9359;
wire net7512;
wire net4920;
wire net5176;
wire net4921;
wire net9242;
wire net4923;
wire net4925;
wire net4928;
wire net8160;
wire net5847;
wire net10977;
wire net6242;
wire net4929;
wire net2194;
wire net4932;
wire net5937;
wire net2341;
wire net4934;
wire net6550;
wire net7578;
wire net4935;
wire net4518;
wire net4936;
wire net4938;
wire net4940;
wire net8324;
wire net4941;
wire net2615;
wire net6917;
wire net4942;
wire net4943;
wire net5581;
wire net7210;
wire net4946;
wire net2961;
wire net745;
wire net4149;
wire net6738;
wire net4947;
wire net4950;
wire net4952;
wire net5111;
wire net4953;
wire net4954;
wire net299;
wire net4956;
wire net6887;
wire net4963;
wire net10790;
wire net10450;
wire net4965;
wire net9849;
wire net6681;
wire net7099;
wire net10093;
wire net7312;
wire net4794;
wire net5444;
wire net1325;
wire net4966;
wire net353;
wire net4968;
wire net5995;
wire net11517;
wire net4969;
wire net4974;
wire net4977;
wire net683;
wire net7247;
wire net4980;
wire net5342;
wire net11288;
wire net4981;
wire net2281;
wire net4982;
wire net11529;
wire net6658;
wire net6674;
wire net4983;
wire net4985;
wire net875;
wire net4986;
wire net4989;
wire net6933;
wire net5282;
wire net6486;
wire net11139;
wire net4992;
wire net8936;
wire net4994;
wire net647;
wire net7043;
wire net4995;
wire net4997;
wire net6323;
wire net11480;
wire net8163;
wire net6300;
wire net4115;
wire net5001;
wire net7886;
wire net5606;
wire net3018;
wire net5003;
wire net6426;
wire net11244;
wire net2744;
wire net5006;
wire net9319;
wire net5008;
wire net5011;
wire net4013;
wire net5012;
wire net5014;
wire net4242;
wire net5015;
wire net10352;
wire net4902;
wire net5018;
wire net8566;
wire net5239;
wire net420;
wire net6304;
wire net7293;
wire net41;
wire net5020;
wire net6804;
wire net5023;
wire net3357;
wire net3674;
wire net5028;
wire net10038;
wire net2179;
wire net5029;
wire net9736;
wire net9706;
wire net5032;
wire net5033;
wire net5034;
wire net1539;
wire net5035;
wire net5039;
wire net5041;
wire net303;
wire net6180;
wire net5045;
wire net5046;
wire net5047;
wire net5050;
wire net5051;
wire net10940;
wire net5056;
wire net4561;
wire net5063;
wire net11349;
wire net7263;
wire net6409;
wire net8351;
wire net6540;
wire net3930;
wire net3792;
wire net7433;
wire net5226;
wire net6981;
wire net5073;
wire net5076;
wire net10502;
wire net5078;
wire net5807;
wire net6163;
wire net5079;
wire net5082;
wire net5083;
wire net7736;
wire net5793;
wire net5085;
wire net5089;
wire net9895;
wire net5094;
wire net6646;
wire net5096;
wire net7460;
wire net950;
wire net5101;
wire net5545;
wire net2598;
wire net4201;
wire net5104;
wire net5107;
wire net5109;
wire net8622;
wire net8581;
wire net5113;
wire net5234;
wire net7432;
wire net7747;
wire net548;
wire net5115;
wire net4029;
wire net5233;
wire net5120;
wire net1810;
wire net5121;
wire net5122;
wire net3287;
wire net5124;
wire net5125;
wire net7689;
wire net5127;
wire net5128;
wire net10013;
wire net6132;
wire net7279;
wire net580;
wire net5130;
wire net9837;
wire net5133;
wire net5134;
wire net10133;
wire net5136;
wire net5137;
wire net6913;
wire net1605;
wire net5138;
wire net3677;
wire net5139;
wire net1612;
wire net5141;
wire net39;
wire net5142;
wire net9498;
wire net5103;
wire net5143;
wire net5144;
wire net5145;
wire net7073;
wire net4195;
wire net5146;
wire net5149;
wire net6961;
wire net9329;
wire net820;
wire net5150;
wire net5151;
wire net5155;
wire net5160;
wire net5162;
wire net9817;
wire net2273;
wire net5163;
wire net5296;
wire net6698;
wire net5168;
wire net9539;
wire net5169;
wire net7844;
wire net814;
wire net5707;
wire net11224;
wire net5170;
wire net5171;
wire net5174;
wire net5175;
wire net6844;
wire net6081;
wire net1111;
wire net5179;
wire net10139;
wire net5181;
wire net5185;
wire net5188;
wire net8154;
wire net5189;
wire net5196;
wire net8401;
wire net5197;
wire net8955;
wire net8670;
wire net5201;
wire net6759;
wire net5203;
wire net5204;
wire net2130;
wire net5205;
wire net5206;
wire net1166;
wire net5209;
wire net2910;
wire net6890;
wire net5212;
wire net7976;
wire net6292;
wire net5213;
wire net5219;
wire net5223;
wire net9945;
wire net6112;
wire net206;
wire net2812;
wire net363;
wire net5228;
wire net2483;
wire net6875;
wire net3136;
wire net5232;
wire net5907;
wire net7206;
wire net2467;
wire net5237;
wire net5240;
wire net6362;
wire net4959;
wire net6119;
wire net1779;
wire net5241;
wire net253;
wire net5244;
wire net5246;
wire net5249;
wire net9189;
wire net5251;
wire net1966;
wire net5252;
wire net7037;
wire net5254;
wire net4424;
wire net5256;
wire net5259;
wire net3353;
wire net4308;
wire net5260;
wire net7398;
wire net5266;
wire net11218;
wire net10298;
wire net5270;
wire net5273;
wire net7288;
wire net6106;
wire net5275;
wire net6333;
wire net4595;
wire net5276;
wire net5280;
wire net8294;
wire net5281;
wire net5286;
wire net2837;
wire net5994;
wire net5290;
wire net1445;
wire net6386;
wire net1038;
wire net5291;
wire net6525;
wire net6164;
wire net5297;
wire net5298;
wire net8515;
wire net4473;
wire net5068;
wire net5300;
wire net5301;
wire net10949;
wire net10213;
wire net5304;
wire net5830;
wire net5307;
wire net4878;
wire net5310;
wire net5311;
wire net2300;
wire net3794;
wire net7265;
wire net9400;
wire net5314;
wire net6536;
wire net5317;
wire net3123;
wire net5320;
wire net1979;
wire net6193;
wire net5323;
wire net3825;
wire net5324;
wire net6901;
wire net5325;
wire net11471;
wire net5327;
wire net9094;
wire net3025;
wire net5813;
wire net5328;
wire net5331;
wire net9996;
wire net5333;
wire net5835;
wire net5334;
wire net9719;
wire net355;
wire net5336;
wire net5337;
wire net8999;
wire net8879;
wire net5338;
wire net5339;
wire net1815;
wire net5340;
wire net5627;
wire net5224;
wire net7195;
wire net5557;
wire net5773;
wire net5352;
wire net10616;
wire net4502;
wire net5353;
wire net11297;
wire net5356;
wire net2196;
wire net6211;
wire net5357;
wire net10427;
wire net4100;
wire net5717;
wire net6232;
wire net9572;
wire net5359;
wire net5615;
wire net5361;
wire net5364;
wire net10776;
wire net8435;
wire net531;
wire net1764;
wire net5365;
wire net6631;
wire net11465;
wire net5366;
wire net5370;
wire net7203;
wire net5374;
wire net5383;
wire net5385;
wire net5390;
wire net5391;
wire net6659;
wire net5393;
wire net5395;
wire net5398;
wire net4704;
wire net5402;
wire net5404;
wire net1535;
wire net5405;
wire net5408;
wire net5413;
wire net5416;
wire net10706;
wire net5417;
wire net5418;
wire net1015;
wire net5419;
wire net26;
wire net5424;
wire net10402;
wire net5425;
wire net5426;
wire net5433;
wire net681;
wire net5435;
wire net5437;
wire net5439;
wire net10484;
wire net5775;
wire net5441;
wire net5442;
wire net10284;
wire net5445;
wire net9527;
wire net5448;
wire net5450;
wire net2925;
wire net5451;
wire net4976;
wire net5452;
wire net7283;
wire net5453;
wire net6626;
wire net104;
wire net5454;
wire net4472;
wire net5459;
wire net6216;
wire net6463;
wire net5461;
wire net5072;
wire net5462;
wire net5466;
wire net5467;
wire net5468;
wire net8491;
wire net7445;
wire net319;
wire net5535;
wire net5470;
wire net5471;
wire net6212;
wire net5472;
wire net5475;
wire net5476;
wire net5477;
wire net7316;
wire net5478;
wire net6867;
wire net6295;
wire net1049;
wire net5479;
wire net5486;
wire net5487;
wire net3020;
wire net850;
wire net1505;
wire net5489;
wire net5490;
wire net5491;
wire net9169;
wire net6140;
wire net5495;
wire net5500;
wire net5501;
wire net6617;
wire net5505;
wire net10668;
wire net5506;
wire net9867;
wire net1156;
wire net5509;
wire net9728;
wire net5618;
wire net6800;
wire net10004;
wire net5510;
wire net5511;
wire net10974;
wire net5513;
wire net1972;
wire net5514;
wire net9230;
wire net9179;
wire net5920;
wire net5515;
wire net5516;
wire net5517;
wire net1719;
wire net5522;
wire net2462;
wire net2059;
wire net1873;
wire net5523;
wire net5526;
wire net5527;
wire net5528;
wire net7464;
wire net5531;
wire net3896;
wire net7289;
wire net5532;
wire net6032;
wire net6407;
wire net2181;
wire net5534;
wire net5537;
wire net352;
wire net5540;
wire net4624;
wire net5541;
wire net5542;
wire net5543;
wire net5544;
wire net5547;
wire net5550;
wire net5551;
wire net3942;
wire net5552;
wire net5562;
wire net1312;
wire net5565;
wire net5566;
wire net5567;
wire net5809;
wire out25;
wire net7649;
wire net5677;
wire net7336;
wire net5942;
wire net7438;
wire net5571;
wire net11030;
wire net111;
wire net5574;
wire net947;
wire net5575;
wire net5157;
wire net5295;
wire net5580;
wire net4210;
wire net5584;
wire net10477;
wire net5585;
wire net4779;
wire net6071;
wire net5587;
wire net5591;
wire net6742;
wire net5592;
wire net5593;
wire net9897;
wire net5595;
wire net1309;
wire net5596;
wire net10021;
wire net7835;
wire net1869;
wire net5600;
wire net5106;
wire net5504;
wire net5601;
wire net6230;
wire net5604;
wire net5605;
wire net7090;
wire net9476;
wire net5608;
wire net3506;
wire net562;
wire net267;
wire net1324;
wire net5611;
wire net4435;
wire net5616;
wire net7620;
wire net5619;
wire net3456;
wire net5620;
wire net5059;
wire net5623;
wire net5631;
wire net5636;
wire net11037;
wire net5640;
wire net2168;
wire net1699;
wire net5641;
wire net7829;
wire net2843;
wire net119;
wire net5642;
wire net568;
wire net5643;
wire net9163;
wire net918;
wire net5644;
wire net5646;
wire net1824;
wire net3261;
wire net5650;
wire net8443;
wire net5651;
wire net5652;
wire net6884;
wire net5653;
wire net5654;
wire net5655;
wire net5657;
wire net6440;
wire net5658;
wire net8559;
wire net2166;
wire net5659;
wire net5662;
wire net10888;
wire net6037;
wire net4365;
wire net7001;
wire net4642;
wire net5663;
wire net5665;
wire net7455;
wire net5666;
wire net5671;
wire net7532;
wire net5052;
wire net5672;
wire net32;
wire net5676;
wire net769;
wire net5679;
wire net10366;
wire net3497;
wire net3404;
wire net5684;
wire net5687;
wire net5770;
wire net5691;
wire net6623;
wire net3659;
wire net5693;
wire net5694;
wire net8848;
wire net4913;
wire net5698;
wire net6213;
wire net5804;
wire net5215;
wire net6653;
wire net5703;
wire net1872;
wire net5705;
wire net9559;
wire net2373;
wire net7174;
wire net7807;
wire net865;
wire net5706;
wire net5708;
wire net2443;
wire net5710;
wire net6819;
wire net266;
wire net5713;
wire net5714;
wire net4480;
wire net4991;
wire net5715;
wire net5716;
wire net8250;
wire net3804;
wire net6169;
wire net5718;
wire net5720;
wire net232;
wire net5721;
wire net5722;
wire net5723;
wire net5725;
wire net5726;
wire net6183;
wire net5729;
wire net9307;
wire net6842;
wire net5731;
wire net5632;
wire net5903;
wire net1128;
wire net4544;
wire net6564;
wire net5732;
wire net7348;
wire net5734;
wire net9135;
wire net5736;
wire net5737;
wire net11526;
wire net5738;
wire net5740;
wire net8540;
wire net4623;
wire net5744;
wire net5747;
wire net6686;
wire net9334;
wire net7057;
wire net3313;
wire net5750;
wire net5751;
wire net5754;
wire net3256;
wire net5755;
wire net5757;
wire net590;
wire net5760;
wire net5761;
wire net8373;
wire net7557;
wire net5316;
wire net5762;
wire net6834;
wire net11149;
wire net9846;
wire net5763;
wire net2607;
wire net7272;
wire net3483;
wire net2635;
wire net1995;
wire net5766;
wire net6253;
wire net5772;
wire net5777;
wire net8800;
wire net5781;
wire net7323;
wire net5783;
wire net6845;
wire net7187;
wire net5785;
wire net7885;
wire net2013;
wire net5786;
wire net4420;
wire net5787;
wire net5788;
wire net7819;
wire net5791;
wire net5796;
wire net5797;
wire net2898;
wire net5798;
wire net5915;
wire net5802;
wire net7739;
wire net5054;
wire net6790;
wire net1154;
wire net5803;
wire net5810;
wire net2860;
wire net5811;
wire net708;
wire net2739;
wire net5739;
wire net6413;
wire net10163;
wire net5812;
wire net5817;
wire net6049;
wire net5818;
wire net5819;
wire net9794;
wire net7284;
wire net2319;
wire net5821;
wire net7025;
wire net1474;
wire net5822;
wire net8561;
wire net2748;
wire net5824;
wire net5825;
wire net5826;
wire net5828;
wire net2286;
wire net5831;
wire net2862;
wire net5004;
wire net5832;
wire net5836;
wire net6822;
wire net5840;
wire net156;
wire net5842;
wire net1662;
wire net6516;
wire net5844;
wire net5805;
wire net6977;
wire net5846;
wire net3477;
wire net5850;
wire net2420;
wire net5851;
wire net764;
wire net5852;
wire net11383;
wire net7400;
wire net10481;
wire net3223;
wire net5854;
wire net5855;
wire net4706;
wire net5856;
wire net7117;
wire net5857;
wire net5859;
wire net10737;
wire net5860;
wire net6155;
wire net5861;
wire net5274;
wire net5862;
wire net5865;
wire net5870;
wire net5871;
wire net5872;
wire net5873;
wire net4322;
wire net5875;
wire net6695;
wire net124;
wire net4890;
wire net5880;
wire net1787;
wire net5888;
wire net8053;
wire net5153;
wire net7024;
wire net9811;
wire net1953;
wire net7454;
wire net10584;
wire net5894;
wire net6812;
wire net5895;
wire net1880;
wire net5896;
wire net5897;
wire net11336;
wire net1058;
wire net5898;
wire net8476;
wire net5853;
wire net5899;
wire net1377;
wire net5901;
wire net5902;
wire net11453;
wire net3765;
wire net5904;
wire net8522;
wire net5905;
wire net5909;
wire net4873;
wire net5910;
wire net400;
wire net5911;
wire net5916;
wire net1847;
wire net5917;
wire net5918;
wire net5919;
wire net5921;
wire net5922;
wire net8697;
wire net7118;
wire net5923;
wire net5927;
wire net10964;
wire net10657;
wire net6279;
wire net5929;
wire net2017;
wire net5931;
wire net5932;
wire net11442;
wire net9834;
wire net5934;
wire net3708;
wire net5935;
wire net2901;
wire net6693;
wire net5938;
wire net9697;
wire net5939;
wire net5414;
wire net305;
wire net5940;
wire net11043;
wire net5945;
wire net7093;
wire net5949;
wire net7602;
wire net5261;
wire net5951;
wire net7389;
wire net9078;
wire net840;
wire net5954;
wire net5753;
wire net5955;
wire net6371;
wire net5956;
wire net1649;
wire net1464;
wire net5957;
wire net5958;
wire net7978;
wire net2590;
wire net5959;
wire net8883;
wire net5960;
wire net9140;
wire net3540;
wire net6471;
wire net10397;
wire net5962;
wire net1123;
wire net5964;
wire net6928;
wire net10110;
wire net1919;
wire net5969;
wire net9120;
wire net6865;
wire net5970;
wire out13;
wire net6189;
wire net9542;
wire net5971;
wire net5972;
wire net5973;
wire net11242;
wire net2582;
wire net5975;
wire net2957;
wire net3816;
wire net5978;
wire net5979;
wire net2912;
wire net5981;
wire net6988;
wire net5982;
wire net754;
wire net5983;
wire net5985;
wire net5988;
wire net5992;
wire net9902;
wire net9815;
wire net2183;
wire net6556;
wire net5996;
wire net3213;
wire net6996;
wire net5998;
wire net6000;
wire net6005;
wire net6007;
wire net7421;
wire net2044;
wire net1752;
wire net1949;
wire net6008;
wire net6009;
wire net2470;
wire net6010;
wire net10449;
wire net6011;
wire net2851;
wire net6012;
wire net6013;
wire net10655;
wire net6014;
wire net1229;
wire net6015;
wire net6018;
wire net2905;
wire net1392;
wire net6020;
wire net6021;
wire net8517;
wire net1825;
wire net6022;
wire net6029;
wire net6030;
wire net6031;
wire net10045;
wire net6290;
wire net5269;
wire net6033;
wire net6034;
wire net8402;
wire net6040;
wire net6041;
wire net9670;
wire net2496;
wire net2052;
wire net6042;
wire net6045;
wire net6047;
wire net6050;
wire net3334;
wire net6051;
wire net6052;
wire net6053;
wire net2611;
wire net4158;
wire net6054;
wire net1061;
wire net6055;
wire net6056;
wire net9458;
wire net6060;
wire net4488;
wire net6061;
wire net11097;
wire net4603;
wire net6457;
wire net6512;
wire net5380;
wire net7123;
wire net5329;
wire net6062;
wire net6065;
wire net6066;
wire net6074;
wire net6075;
wire net11506;
wire net228;
wire net5178;
wire net6076;
wire net10062;
wire net6078;
wire net6080;
wire net6082;
wire net6083;
wire net11089;
wire net6085;
wire net6086;
wire net6143;
wire net2619;
wire net2190;
wire net6087;
wire net6090;
wire net3636;
wire net6091;
wire net4056;
wire net6093;
wire net7175;
wire net431;
wire net6098;
wire net3271;
wire net5231;
wire net6100;
wire net7826;
wire net6101;
wire net1294;
wire net6102;
wire net5409;
wire net6628;
wire net8302;
wire net1527;
wire net6158;
wire net6103;
wire net3051;
wire net6104;
wire net1041;
wire net5250;
wire net6105;
wire net7386;
wire net6108;
wire net6109;
wire net4804;
wire net6110;
wire net1263;
wire net1397;
wire net6111;
wire net6113;
wire net6399;
wire net6117;
wire net1349;
wire net6118;
wire net1352;
wire net6121;
wire net6126;
wire net6127;
wire net6129;
wire net1273;
wire net6130;
wire net1561;
wire net6133;
wire net6134;
wire net6135;
wire net4537;
wire net7213;
wire net6136;
wire net6137;
wire net6138;
wire net6139;
wire net6141;
wire net8176;
wire net6144;
wire net6146;
wire net1070;
wire net6888;
wire net10090;
wire net6154;
wire net7097;
wire net8309;
wire net6162;
wire net6902;
wire net6165;
wire net6167;
wire net7191;
wire net11060;
wire net7981;
wire net6289;
wire net6168;
wire net6171;
wire net7299;
wire net7893;
wire net6174;
wire net7903;
wire net7443;
wire net6175;
wire net8258;
wire net6177;
wire net10537;
wire net5110;
wire net6181;
wire net6173;
wire net6182;
wire net10233;
wire net6184;
wire net6185;
wire net10035;
wire net6187;
wire net5474;
wire net1902;
wire net1540;
wire net6190;
wire net2342;
wire net6195;
wire net6196;
wire net9206;
wire net6602;
wire net1715;
wire net6199;
wire net6200;
wire net10457;
wire net6201;
wire net6206;
wire net6208;
wire net9047;
wire net6004;
wire net6209;
wire net7757;
wire net4854;
wire net6210;
wire net6215;
wire net2109;
wire net6217;
wire net3514;
wire net6219;
wire net6220;
wire net11136;
wire net6222;
wire net3412;
wire net341;
wire net6223;
wire net6224;
wire net6227;
wire net4134;
wire net6231;
wire net6233;
wire net5016;
wire net6235;
wire net2546;
wire net6259;
wire net6236;
wire net9590;
wire net1728;
wire net6811;
wire net6238;
wire net7682;
wire net6239;
wire net6241;
wire net6243;
wire net6244;
wire net9123;
wire net1537;
wire net5667;
wire net5570;
wire net6246;
wire net7003;
wire net2035;
wire net1529;
wire net6247;
wire net6250;
wire net2158;
wire net6392;
wire net8147;
wire net6254;
wire net11275;
wire net6257;
wire net6258;
wire net9888;
wire net5686;
wire net4911;
wire net6260;
wire net6261;
wire net9954;
wire net6262;
wire net8647;
wire net8601;
wire net1345;
wire net6263;
wire net4459;
wire net136;
wire net6265;
wire net4718;
wire net6266;
wire net8307;
wire net6269;
wire net6270;
wire net6271;
wire net6273;
wire net6274;
wire net6276;
wire net9048;
wire net6282;
wire net7846;
wire net6283;
wire net6571;
wire net6284;
wire net6285;
wire net6286;
wire net6899;
wire net6287;
wire net6291;
wire net8783;
wire net1647;
wire net6293;
wire net1807;
wire net6294;
wire net2395;
wire net1891;
wire net6301;
wire net6305;
wire net3012;
wire net6306;
wire net2124;
wire net6918;
wire net6308;
wire net11380;
wire net1957;
wire net1096;
wire net2225;
wire net4088;
wire net6309;
wire net2762;
wire net6313;
wire net6314;
wire net9716;
wire net6406;
wire net8349;
wire net6096;
wire net6315;
wire net6317;
wire net6318;
wire net8291;
wire net6319;
wire net6321;
wire net9321;
wire net6325;
wire net2711;
wire net6326;
wire net6327;
wire net8037;
wire net595;
wire net6328;
wire net7125;
wire net6330;
wire net10128;
wire net5081;
wire net6331;
wire net6334;
wire net8180;
wire net6336;
wire net9243;
wire net6338;
wire net4307;
wire net6339;
wire net6341;
wire net8078;
wire net6468;
wire net6342;
wire net6343;
wire net6346;
wire net3583;
wire net2553;
wire net1107;
wire net6347;
wire net6348;
wire net6349;
wire net6352;
wire net6355;
wire net6359;
wire net10443;
wire net6374;
wire net6505;
wire net6364;
wire net7154;
wire net6365;
wire net9413;
wire net427;
wire net6367;
wire net8036;
wire net6369;
wire net11180;
wire net8792;
wire net6372;
wire net6375;
wire net6377;
wire net6378;
wire net2051;
wire net6379;
wire net9460;
wire net6382;
wire net6383;
wire net10495;
wire net6384;
wire net6388;
wire net6389;
wire net169;
wire net6391;
wire net10058;
wire net6394;
wire net3131;
wire net6396;
wire net6739;
wire net11268;
wire net8224;
wire net6397;
wire net6401;
wire net6402;
wire net6405;
wire net8962;
wire net6408;
wire net6491;
wire net6411;
wire net6753;
wire net6412;
wire net8886;
wire net1004;
wire net6415;
wire net6784;
wire net11029;
wire net1047;
wire net6418;
wire net11096;
wire net9655;
wire net6420;
wire net7667;
wire net2685;
wire net6903;
wire net6424;
wire net6428;
wire net7002;
wire net687;
wire net1412;
wire net7179;
wire net3742;
wire net6430;
wire net4121;
wire net6433;
wire net3472;
wire net6439;
wire net4270;
wire net6443;
wire net6444;
wire net6445;
wire net9681;
wire net6446;
wire net8246;
wire net5878;
wire net6447;
wire net3750;
wire net4391;
wire net6452;
wire net6453;
wire net6454;
wire net7039;
wire net6456;
wire net11485;
wire net6459;
wire net6460;
wire net3385;
wire net6469;
wire net6475;
wire net1898;
wire net6477;
wire net6478;
wire net6479;
wire net1546;
wire net6480;
wire net7717;
wire net7161;
wire net4639;
wire net6487;
wire net6489;
wire net6493;
wire net1140;
wire net6494;
wire net6497;
wire net9471;
wire net6499;
wire net6501;
wire net5431;
wire net6503;
wire net5863;
wire net6535;
wire net6603;
wire net6507;
wire net6508;
wire net5733;
wire net7480;
wire net7542;
wire net6511;
wire net10589;
wire net10083;
wire net6513;
wire net6514;
wire net9543;
wire net6515;
wire net6562;
wire net6518;
wire net11207;
wire net2963;
wire net6519;
wire net243;
wire net6520;
wire net1390;
wire net6523;
wire net6524;
wire net7709;
wire net4741;
wire net6823;
wire net6527;
wire net6529;
wire net11539;
wire net8122;
wire net6077;
wire net6533;
wire net10068;
wire net6538;
wire net6544;
wire net6547;
wire net6552;
wire net2348;
wire net6553;
wire net6554;
wire net6685;
wire net7393;
wire net6557;
wire net5634;
wire net6558;
wire net10010;
wire net2820;
wire net6559;
wire net6561;
wire net6563;
wire net6567;
wire net9102;
wire net1583;
wire net5546;
wire net6568;
wire net10471;
wire net6570;
wire net1102;
wire net6575;
wire net4019;
wire net6577;
wire net1138;
wire net6581;
wire net11345;
wire net10459;
wire net10325;
wire net3324;
wire net6582;
wire net9067;
wire net6583;
wire net781;
wire net6599;
wire net6586;
wire net6587;
wire net9702;
wire net6588;
wire net6589;
wire net6202;
wire net6590;
wire net6592;
wire net7534;
wire net6593;
wire net586;
wire net4514;
wire net7391;
wire net5438;
wire net6597;
wire net6605;
wire net6608;
wire net8079;
wire net6609;
wire net6632;
wire net3359;
wire net6610;
wire net10993;
wire net6611;
wire net8248;
wire net471;
wire net6613;
wire net6614;
wire net3614;
wire net4538;
wire net6615;
wire net6616;
wire net6620;
wire net4312;
wire net6621;
wire net6624;
wire net6627;
wire net9558;
wire net6633;
wire net6643;
wire net6648;
wire net6650;
wire net9874;
wire net6656;
wire net8490;
wire net6662;
wire net277;
wire net6665;
wire net5869;
wire net6670;
wire net6672;
wire net6675;
wire net6678;
wire net5848;
wire net6679;
wire net6683;
wire net2350;
wire net6688;
wire net4681;
wire net6690;
wire net6694;
wire net6696;
wire net6704;
wire net1337;
wire net827;
wire net6709;
wire net11117;
wire net7734;
wire net5484;
wire net4984;
wire net6969;
wire net6710;
wire net8892;
wire net3675;
wire net5065;
wire net6711;
wire net3746;
wire net6713;
wire net10392;
wire net6716;
wire net6719;
wire net2410;
wire net6340;
wire net6722;
wire net6726;
wire net7252;
wire net6728;
wire net5521;
wire net6729;
wire net8757;
wire net6734;
wire net4582;
wire net5187;
wire net6736;
wire net547;
wire net6741;
wire net6746;
wire net6747;
wire net9501;
wire net1198;
wire net6748;
wire net6749;
wire net6750;
wire net3253;
wire net6751;
wire net6752;
wire net3190;
wire net1328;
wire net6754;
wire net10188;
wire net9763;
wire net5220;
wire net6755;
wire net6929;
wire net6756;
wire net10643;
wire net6757;
wire net6762;
wire net11226;
wire net10697;
wire net7334;
wire net5318;
wire net6765;
wire net5968;
wire net6768;
wire net2340;
wire net6769;
wire net7232;
wire net6771;
wire net10373;
wire net6772;
wire net2382;
wire net109;
wire net7437;
wire net6773;
wire net1362;
wire net7146;
wire net6775;
wire net6777;
wire net6778;
wire net987;
wire net7236;
wire net6779;
wire net7050;
wire net6780;
wire net5997;
wire net6781;
wire net6794;
wire net6783;
wire net9664;
wire net165;
wire net4573;
wire net6788;
wire net6789;
wire net7062;
wire net6795;
wire net6207;
wire net6798;
wire net6801;
wire net3079;
wire net6802;
wire net7150;
wire net6803;
wire net6805;
wire net6807;
wire net6808;
wire net1659;
wire net6809;
wire net6814;
wire net6815;
wire net8700;
wire net6099;
wire net6817;
wire net6820;
wire net6825;
wire net4353;
wire net6827;
wire net11182;
wire net1782;
wire net6828;
wire net8794;
wire net6829;
wire net1988;
wire net6830;
wire net8583;
wire net6831;
wire net9563;
wire net6833;
wire net6835;
wire net6836;
wire net6837;
wire net806;
wire net6840;
wire net2207;
wire net5795;
wire net6841;
wire net6846;
wire net6847;
wire net6848;
wire net6851;
wire net9024;
wire net6854;
wire net11193;
wire net5569;
wire net6855;
wire net6857;
wire net8944;
wire net6859;
wire net151;
wire net6860;
wire net1905;
wire net6863;
wire net540;
wire net6869;
wire net6870;
wire net8052;
wire net1275;
wire net2315;
wire net6871;
wire net11261;
wire net6873;
wire net5330;
wire net6874;
wire net1582;
wire net6878;
wire net6880;
wire net9593;
wire net6883;
wire net6886;
wire net6889;
wire net6891;
wire net9832;
wire net325;
wire net56;
wire net6893;
wire net6896;
wire net1794;
wire net6898;
wire net5771;
wire net6900;
wire net2148;
wire net4346;
wire net7375;
wire net6904;
wire net11436;
wire net6906;
wire net6910;
wire net705;
wire net6912;
wire net6920;
wire net6925;
wire net10349;
wire net9718;
wire net6926;
wire net6931;
wire net5594;
wire net6935;
wire net4406;
wire net6937;
wire net6938;
wire net6939;
wire net4004;
wire net6942;
wire net1151;
wire net6943;
wire net6944;
wire net4175;
wire net6945;
wire net6947;
wire net399;
wire net6950;
wire net6952;
wire net6953;
wire net2993;
wire net6955;
wire net3863;
wire net6959;
wire net4407;
wire net6962;
wire net6963;
wire net4649;
wire net6964;
wire net2977;
wire net6966;
wire net786;
wire net7114;
wire net6967;
wire net3135;
wire net6970;
wire net2664;
wire net6972;
wire net6974;
wire net6983;
wire net10406;
wire net2682;
wire net6984;
wire net7121;
wire net6027;
wire net6985;
wire net413;
wire net6992;
wire net9842;
wire net7446;
wire net6995;
wire net7580;
wire net3987;
wire net6999;
wire net11055;
wire net7004;
wire net8137;
wire net805;
wire net7005;
wire net1239;
wire net7007;
wire net6024;
wire net5211;
wire net7008;
wire net7010;
wire net7012;
wire net7013;
wire net7014;
wire net7017;
wire net7019;
wire net7697;
wire net7228;
wire net10528;
wire net7020;
wire net7027;
wire net7030;
wire net7032;
wire net7033;
wire net7035;
wire net7036;
wire net7038;
wire net2186;
wire net7096;
wire net7040;
wire net9560;
wire net5868;
wire net7041;
wire net7992;
wire net7045;
wire net7049;
wire net7052;
wire net7055;
wire net23;
wire net7056;
wire net7058;
wire net7063;
wire net3501;
wire net3656;
wire net1805;
wire net7064;
wire net9910;
wire net1334;
wire net7066;
wire net7068;
wire net7077;
wire net7083;
wire net4563;
wire net7086;
wire net10273;
wire net304;
wire net7087;
wire net1370;
wire net7088;
wire net5005;
wire net7089;
wire net7091;
wire net7842;
wire net7098;
wire net7325;
wire net3806;
wire net7100;
wire net7105;
wire net7106;
wire net5102;
wire net7108;
wire net9914;
wire net7110;
wire net8565;
wire net7112;
wire net3553;
wire net7113;
wire net7116;
wire net7119;
wire net7128;
wire net7129;
wire net7133;
wire net11531;
wire net7783;
wire net2727;
wire net7134;
wire net10803;
wire net10441;
wire net7135;
wire net7136;
wire net7138;
wire net10521;
wire net7140;
wire net7141;
wire net7143;
wire net5689;
wire net7144;
wire net7148;
wire net9487;
wire net7149;
wire net7673;
wire net6718;
wire net7152;
wire net9971;
wire net4843;
wire net7157;
wire net11576;
wire net1624;
wire net7160;
wire net1320;
wire net7163;
wire net7851;
wire net7164;
wire net7165;
wire net1290;
wire net7167;
wire net5701;
wire net7168;
wire net7169;
wire net7496;
wire net6192;
wire net7171;
wire net1436;
wire net7172;
wire net9216;
wire net7173;
wire net7180;
wire net8535;
wire net7181;
wire net4320;
wire net7186;
wire net322;
wire net7188;
wire net7197;
wire net1176;
wire net7198;
wire net575;
wire net7199;
wire net1109;
wire net7200;
wire net307;
wire net7201;
wire net3733;
wire net7205;
wire net7207;
wire net7208;
wire net7209;
wire net7211;
wire net1708;
wire net7212;
wire net7076;
wire net7214;
wire net7215;
wire net9428;
wire net7217;
wire net7222;
wire net10975;
wire net9456;
wire net9109;
wire net7224;
wire net7225;
wire net9835;
wire net7067;
wire net7227;
wire net7229;
wire net9915;
wire net5941;
wire net7233;
wire net9395;
wire net3022;
wire net7234;
wire net8270;
wire net4310;
wire net7238;
wire net7240;
wire net7882;
wire net7243;
wire net5293;
wire net7248;
wire net7251;
wire net11066;
wire net7253;
wire net5892;
wire net1812;
wire net7254;
wire net6622;
wire net7255;
wire net5885;
wire net7258;
wire net7264;
wire net7780;
wire net4465;
wire net7266;
wire net7274;
wire net1875;
wire net7275;
wire net6635;
wire net7277;
wire net7280;
wire net7287;
wire net4456;
wire net7291;
wire net9999;
wire net7292;
wire net7297;
wire net7298;
wire net7301;
wire net1877;
wire net7304;
wire net7305;
wire net9008;
wire net7307;
wire net7308;
wire net3865;
wire net7313;
wire net7317;
wire net9564;
wire net7318;
wire net1680;
wire net7322;
wire net10744;
wire net7333;
wire net10740;
wire net7337;
wire net9232;
wire net7339;
wire net7340;
wire net7341;
wire net7342;
wire net7343;
wire net7350;
wire net8364;
wire net6521;
wire net7351;
wire net7352;
wire net1430;
wire net7357;
wire net7360;
wire net7362;
wire net7434;
wire net8473;
wire net7365;
wire net7366;
wire net7367;
wire net7574;
wire net3351;
wire net7369;
wire net11074;
wire net7371;
wire net5765;
wire net7373;
wire net9495;
wire net7376;
wire net8659;
wire net7377;
wire net7380;
wire net5343;
wire net7383;
wire net1019;
wire net7392;
wire net9546;
wire net7394;
wire net10170;
wire net61;
wire net7395;
wire net7397;
wire net7399;
wire net7401;
wire net9552;
wire net7403;
wire net1781;
wire net7404;
wire net7405;
wire net9472;
wire net7407;
wire net3778;
wire net6161;
wire net4468;
wire net3815;
wire net6116;
wire net7409;
wire net11171;
wire net10569;
wire net7411;
wire net7412;
wire net3515;
wire net4566;
wire net7413;
wire net10557;
wire net7420;
wire net6810;
wire net7422;
wire net2063;
wire net3883;
wire net6450;
wire net7424;
wire net11372;
wire net4047;
wire net7426;
wire net4244;
wire net7436;
wire net6495;
wire net7153;
wire net7439;
wire net7442;
wire net7447;
wire net5463;
wire net7448;
wire net7449;
wire net7451;
wire net11525;
wire net2900;
wire net7452;
wire net7856;
wire net7453;
wire net10978;
wire net7456;
wire net7459;
wire net4025;
wire net7468;
wire net10608;
wire net7471;
wire net3281;
wire net7472;
wire net7473;
wire net10832;
wire net5285;
wire net7474;
wire net7477;
wire net2173;
wire net7478;
wire net3606;
wire net7479;
wire net7482;
wire net3368;
wire net7485;
wire net7486;
INV_X32 c26(
.A(in20),
.ZN(net0)
);

INV_X4 c27(
.A(in17),
.ZN(net1)
);

XOR2_X2 c28(
.A(net0),
.B(in11),
.Z(net2)
);

INV_X1 c29(
.A(in10),
.ZN(net3)
);

XNOR2_X1 c30(
.A(net3),
.B(in2),
.ZN(net4)
);

INV_X2 c31(
.A(in8),
.ZN(net5)
);

INV_X8 c32(
.A(in17),
.ZN(net6)
);

INV_X16 c33(
.A(in2),
.ZN(net7)
);

OR3_X2 c34(
.A1(in21),
.A2(in9),
.A3(net0),
.ZN(net8)
);

INV_X32 c35(
.A(net8),
.ZN(net9)
);

OR2_X4 c36(
.A1(in22),
.A2(net2),
.ZN(net10)
);

INV_X4 c37(
.A(in3),
.ZN(net11)
);

OAI21_X2 c38(
.A(net9),
.B1(in6),
.B2(net40),
.ZN(net12)
);

OR2_X1 c39(
.A1(net5),
.A2(net3),
.ZN(net13)
);

XNOR2_X2 c40(
.A(net39),
.B(net2),
.ZN(net14)
);

OAI21_X1 c41(
.A(net7),
.B1(in0),
.B2(in12),
.ZN(net15)
);

INV_X1 c42(
.A(net10),
.ZN(net16)
);

INV_X2 c43(
.A(in15),
.ZN(net17)
);

INV_X8 c44(
.A(net39),
.ZN(net18)
);

INV_X16 c45(
.A(in6),
.ZN(net19)
);

INV_X32 c46(
.A(net17),
.ZN(net20)
);

AND2_X4 c47(
.A1(net18),
.A2(net39),
.ZN(net21)
);

INV_X4 c48(
.A(net14),
.ZN(net22)
);

INV_X1 c49(
.A(net22),
.ZN(net23)
);

INV_X2 c50(
.A(net3),
.ZN(net24)
);

INV_X8 c51(
.A(net8),
.ZN(net25)
);

AND2_X1 c52(
.A1(in0),
.A2(net2),
.ZN(net26)
);

INV_X16 c53(
.A(net23),
.ZN(net27)
);

INV_X32 c54(
.A(net1),
.ZN(net28)
);

AOI21_X2 c55(
.A(net23),
.B1(net27),
.B2(net18),
.ZN(net29)
);

INV_X4 c56(
.A(net28),
.ZN(net30)
);

INV_X1 c57(
.A(net20),
.ZN(net31)
);

AOI21_X1 c58(
.A(net13),
.B1(net1),
.B2(net31),
.ZN(net32)
);

NAND2_X1 c59(
.A1(net30),
.A2(net29),
.ZN(net33)
);

AOI21_X4 c60(
.A(net26),
.B1(net30),
.B2(net33),
.ZN(net34)
);

INV_X2 c61(
.A(net12),
.ZN(net35)
);

NAND2_X2 c62(
.A1(in22),
.A2(net31),
.ZN(net36)
);

NAND2_X4 c63(
.A1(net31),
.A2(net34),
.ZN(net37)
);

INV_X8 c64(
.A(in11),
.ZN(net38)
);

INV_X16 c65(
.A(in1),
.ZN(net39)
);

INV_X32 c66(
.A(in16),
.ZN(net40)
);

AND3_X1 c67(
.A1(net34),
.A2(in5),
.A3(net31),
.ZN(net41)
);

NAND3_X1 c68(
.A1(net2),
.A2(net31),
.A3(net3),
.ZN(net42)
);

INV_X4 c69(
.A(net42),
.ZN(net43)
);

NOR3_X4 c70(
.A1(net16),
.A2(net42),
.A3(net32),
.ZN(net44)
);

INV_X1 c71(
.A(net27),
.ZN(net45)
);

AND2_X2 c72(
.A1(in3),
.A2(net43),
.ZN(net46)
);

NOR3_X2 c73(
.A1(net32),
.A2(in18),
.A3(net45),
.ZN(net47)
);

XOR2_X1 c74(
.A(net40),
.B(net42),
.Z(net48)
);

NOR2_X1 c75(
.A1(net44),
.A2(in20),
.ZN(net49)
);

AND3_X4 c76(
.A1(net38),
.A2(net20),
.A3(net4),
.ZN(net50)
);

NAND3_X2 c77(
.A1(net15),
.A2(net38),
.A3(net12),
.ZN(net51)
);

OR3_X1 c78(
.A1(net4),
.A2(net10),
.A3(net11),
.ZN(net52)
);

MUX2_X1 c79(
.A(net11),
.B(net30),
.S(net49),
.Z(net53)
);

OAI21_X4 c80(
.A(net28),
.B1(net53),
.B2(net39),
.ZN(net54)
);

MUX2_X2 c81(
.A(net54),
.B(net44),
.S(in16),
.Z(net55)
);

NAND3_X4 c82(
.A1(net25),
.A2(net54),
.A3(net39),
.ZN(net56)
);

OR2_X2 c83(
.A1(net43),
.A2(net30),
.ZN(net57)
);

INV_X2 c84(
.A(net9771),
.ZN(net58)
);

INV_X8 c85(
.A(net30),
.ZN(net59)
);

OR3_X4 c86(
.A1(net24),
.A2(net108),
.A3(in13),
.ZN(net60)
);

INV_X16 c87(
.A(net47),
.ZN(net61)
);

NOR2_X4 c88(
.A1(net49),
.A2(net107),
.ZN(net62)
);

INV_X32 c89(
.A(net10535),
.ZN(net63)
);

INV_X4 c90(
.A(in14),
.ZN(net64)
);

INV_X1 c91(
.A(net40),
.ZN(net65)
);

INV_X2 c92(
.A(in13),
.ZN(net66)
);

INV_X8 c93(
.A(net36),
.ZN(net67)
);

INV_X16 c94(
.A(net43),
.ZN(net68)
);

INV_X32 c95(
.A(net9771),
.ZN(net69)
);

DFFR_X1 c96(
.D(net58),
.RN(net108),
.CK(clk),
.Q(net71),
.QN(net70)
);

INV_X4 c97(
.A(net107),
.ZN(net72)
);

INV_X1 c98(
.A(net36),
.ZN(net73)
);

INV_X2 c99(
.A(net106),
.ZN(net74)
);

INV_X8 c100(
.A(net72),
.ZN(net75)
);

NOR2_X2 c101(
.A1(in8),
.A2(net24),
.ZN(net76)
);

XOR2_X2 c102(
.A(net24),
.B(net40),
.Z(net77)
);

XNOR2_X1 c103(
.A(net69),
.B(net74),
.ZN(net78)
);

INV_X16 c104(
.A(net64),
.ZN(net79)
);

INV_X32 c105(
.A(net62),
.ZN(net80)
);

OR2_X4 c106(
.A1(net73),
.A2(net74),
.ZN(net81)
);

INV_X4 c107(
.A(net71),
.ZN(net82)
);

INV_X1 c108(
.A(net65),
.ZN(net83)
);

OR2_X1 c109(
.A1(net81),
.A2(net68),
.ZN(net84)
);

INV_X2 c110(
.A(net61),
.ZN(net85)
);

INV_X8 c111(
.A(net76),
.ZN(net86)
);

XNOR2_X2 c112(
.A(net73),
.B(net83),
.ZN(net87)
);

INV_X16 c113(
.A(net55),
.ZN(net88)
);

INV_X32 c114(
.A(in10),
.ZN(net89)
);

INV_X4 c115(
.A(net89),
.ZN(net90)
);

INV_X1 c116(
.A(net64),
.ZN(net91)
);

AND2_X4 c117(
.A1(net85),
.A2(net106),
.ZN(net92)
);

INV_X2 c118(
.A(net72),
.ZN(net93)
);

INV_X8 c119(
.A(net84),
.ZN(net94)
);

INV_X16 c120(
.A(net87),
.ZN(net95)
);

AND2_X1 c121(
.A1(net61),
.A2(net40),
.ZN(net96)
);

INV_X32 c122(
.A(net63),
.ZN(net97)
);

INV_X4 c123(
.A(net91),
.ZN(net98)
);

DFFR_X2 c124(
.D(net82),
.RN(net37),
.CK(clk),
.Q(net100),
.QN(net99)
);

NAND2_X1 c125(
.A1(net22),
.A2(net99),
.ZN(net101)
);

INV_X1 c126(
.A(in1),
.ZN(net102)
);

NAND2_X2 c127(
.A1(net69),
.A2(net55),
.ZN(net103)
);

DFFRS_X1 c128(
.D(net97),
.RN(net103),
.SN(net91),
.CK(clk),
.Q(net105),
.QN(net104)
);

INV_X2 c129(
.A(net13),
.ZN(net106)
);

INV_X8 c130(
.A(in14),
.ZN(net107)
);

INV_X16 c131(
.A(net55),
.ZN(net108)
);

INV_X32 c132(
.A(in18),
.ZN(net109)
);

INV_X4 c133(
.A(net80),
.ZN(net110)
);

DFFS_X1 c134(
.D(net83),
.SN(net85),
.CK(clk),
.Q(net112),
.QN(net111)
);

INV_X1 c135(
.A(net48),
.ZN(net113)
);

INV_X2 c136(
.A(net94),
.ZN(net114)
);

INV_X8 c137(
.A(net114),
.ZN(net115)
);

DFFS_X2 c138(
.D(net85),
.SN(net88),
.CK(clk),
.Q(net117),
.QN(net116)
);

NAND2_X4 c139(
.A1(net84),
.A2(net91),
.ZN(net118)
);

AND3_X2 c140(
.A1(net114),
.A2(net98),
.A3(net83),
.ZN(net119)
);

DFFR_X1 c141(
.D(net119),
.RN(net91),
.CK(clk),
.Q(net121),
.QN(net120)
);

DFFR_X2 c142(
.D(net115),
.RN(net111),
.CK(clk),
.Q(net123),
.QN(net122)
);

AND2_X2 c143(
.A1(net90),
.A2(net94),
.ZN(net124)
);

XOR2_X1 c144(
.A(net65),
.B(net110),
.Z(net125)
);

NOR2_X1 c145(
.A1(net122),
.A2(net10534),
.ZN(net126)
);

OR2_X2 c146(
.A1(net107),
.A2(net63),
.ZN(net127)
);

DFFRS_X2 c147(
.D(net103),
.RN(net55),
.SN(net75),
.CK(clk),
.Q(net129),
.QN(net128)
);

DFFS_X1 c148(
.D(net75),
.SN(net37),
.CK(clk),
.Q(net131),
.QN(net130)
);

DFFS_X2 c149(
.D(net88),
.SN(net126),
.CK(clk),
.Q(net133),
.QN(net132)
);

NOR2_X4 c150(
.A1(net131),
.A2(net58),
.ZN(net134)
);

NOR2_X2 c151(
.A1(net127),
.A2(net102),
.ZN(net135)
);

DFFR_X1 c152(
.D(net81),
.RN(net119),
.CK(clk),
.Q(net137),
.QN(net136)
);

XOR2_X2 c153(
.A(in18),
.B(net124),
.Z(net138)
);

NOR3_X1 c154(
.A1(net135),
.A2(net120),
.A3(net127),
.ZN(net139)
);

XNOR2_X1 c155(
.A(net98),
.B(net93),
.ZN(net140)
);

OR3_X2 c156(
.A1(net80),
.A2(net134),
.A3(net139),
.ZN(net141)
);

DFFR_X2 c157(
.D(net125),
.RN(net130),
.CK(clk),
.Q(net143),
.QN(net142)
);

OAI21_X2 c158(
.A(net112),
.B1(net128),
.B2(net142),
.ZN(net144)
);

SDFFRS_X1 c159(
.D(net139),
.RN(net141),
.SE(net140),
.SI(net124),
.SN(net88),
.CK(clk),
.Q(net146),
.QN(net145)
);

OAI21_X1 c160(
.A(net143),
.B1(net133),
.B2(net144),
.ZN(net147)
);

AOI21_X2 c161(
.A(net89),
.B1(net135),
.B2(net124),
.ZN(net148)
);

SDFFRS_X2 c162(
.D(net134),
.RN(net82),
.SE(net125),
.SI(net127),
.SN(net124),
.CK(clk),
.Q(net150),
.QN(net149)
);

AOI21_X1 c163(
.A(net129),
.B1(net5),
.B2(net73),
.ZN(net151)
);

AOI21_X4 c164(
.A(net140),
.B1(net104),
.B2(net143),
.ZN(net152)
);

OAI221_X4 c165(
.A(net105),
.B1(net151),
.B2(net147),
.C1(net136),
.C2(net124),
.ZN(net153)
);

INV_X16 c166(
.A(net77),
.ZN(net154)
);

INV_X32 c167(
.A(net48),
.ZN(net155)
);

OR2_X4 c168(
.A1(net155),
.A2(net95),
.ZN(net156)
);

INV_X4 c169(
.A(net9731),
.ZN(net157)
);

INV_X1 c170(
.A(in4),
.ZN(net158)
);

INV_X2 c171(
.A(net146),
.ZN(net159)
);

INV_X8 c172(
.A(net34),
.ZN(net160)
);

INV_X16 c173(
.A(net156),
.ZN(net161)
);

OR2_X1 c174(
.A1(net158),
.A2(net53),
.ZN(net162)
);

INV_X32 c175(
.A(net149),
.ZN(net163)
);

INV_X4 c176(
.A(net59),
.ZN(net164)
);

INV_X1 c177(
.A(net117),
.ZN(net165)
);

INV_X2 c178(
.A(net161),
.ZN(net166)
);

INV_X8 c179(
.A(net79),
.ZN(net167)
);

INV_X16 c180(
.A(net124),
.ZN(net168)
);

INV_X32 c181(
.A(net146),
.ZN(net169)
);

INV_X4 c182(
.A(net9731),
.ZN(net170)
);

INV_X1 c183(
.A(net169),
.ZN(net171)
);

XNOR2_X2 c184(
.A(net123),
.B(net116),
.ZN(net172)
);

AND3_X1 c185(
.A1(net123),
.A2(net116),
.A3(net86),
.ZN(net173)
);

INV_X2 c186(
.A(net152),
.ZN(net174)
);

INV_X8 c187(
.A(net53),
.ZN(net175)
);

AND2_X4 c188(
.A1(net172),
.A2(net136),
.ZN(net176)
);

INV_X16 c189(
.A(net154),
.ZN(net177)
);

INV_X32 c190(
.A(net170),
.ZN(net178)
);

INV_X4 c191(
.A(net101),
.ZN(net179)
);

AND2_X1 c192(
.A1(net151),
.A2(net176),
.ZN(net180)
);

INV_X1 c193(
.A(net178),
.ZN(net181)
);

INV_X2 c194(
.A(net177),
.ZN(net182)
);

INV_X8 c195(
.A(net9860),
.ZN(net183)
);

INV_X16 c196(
.A(net181),
.ZN(net184)
);

NAND2_X1 c197(
.A1(net175),
.A2(net53),
.ZN(net185)
);

NAND2_X2 c198(
.A1(net175),
.A2(net163),
.ZN(net186)
);

INV_X32 c199(
.A(in4),
.ZN(net187)
);

INV_X4 c200(
.A(net117),
.ZN(net188)
);

INV_X1 c201(
.A(net184),
.ZN(net189)
);

INV_X2 c202(
.A(in21),
.ZN(net190)
);

NAND2_X4 c203(
.A1(net77),
.A2(net173),
.ZN(net191)
);

NAND3_X1 c204(
.A1(net186),
.A2(net155),
.A3(net101),
.ZN(net192)
);

INV_X8 c205(
.A(net169),
.ZN(net193)
);

NOR3_X4 c206(
.A1(net150),
.A2(net48),
.A3(net183),
.ZN(net194)
);

AND2_X2 c207(
.A1(net190),
.A2(net165),
.ZN(net195)
);

XOR2_X1 c208(
.A(net183),
.B(net127),
.Z(net196)
);

NOR2_X1 c209(
.A1(net173),
.A2(net86),
.ZN(net197)
);

INV_X16 c210(
.A(net53),
.ZN(net198)
);

INV_X32 c211(
.A(net10931),
.ZN(net199)
);

INV_X4 c212(
.A(net180),
.ZN(net200)
);

OR2_X2 c213(
.A1(net197),
.A2(net164),
.ZN(net201)
);

NOR2_X4 c214(
.A1(net187),
.A2(net178),
.ZN(net202)
);

NOR2_X2 c215(
.A1(net152),
.A2(net157),
.ZN(net203)
);

INV_X1 c216(
.A(net201),
.ZN(net204)
);

INV_X2 c217(
.A(net201),
.ZN(net205)
);

NOR3_X2 c218(
.A1(net200),
.A2(net180),
.A3(net190),
.ZN(net206)
);

XOR2_X2 c219(
.A(net193),
.B(net175),
.Z(net207)
);

XNOR2_X1 c220(
.A(net207),
.B(net124),
.ZN(net208)
);

INV_X8 c221(
.A(net161),
.ZN(net209)
);

INV_X16 c222(
.A(net10892),
.ZN(net210)
);

AND3_X4 c223(
.A1(net205),
.A2(net178),
.A3(net191),
.ZN(net211)
);

INV_X32 c224(
.A(net101),
.ZN(net212)
);

DFFS_X1 c225(
.D(net177),
.SN(net208),
.CK(clk),
.Q(net214),
.QN(net213)
);

OR2_X4 c226(
.A1(net211),
.A2(net175),
.ZN(net215)
);

OR2_X1 c227(
.A1(net164),
.A2(net213),
.ZN(net216)
);

NAND3_X2 c228(
.A1(net79),
.A2(net203),
.A3(net208),
.ZN(net217)
);

INV_X4 c229(
.A(net206),
.ZN(net218)
);

OR3_X1 c230(
.A1(net182),
.A2(net122),
.A3(net10642),
.ZN(net219)
);

XNOR2_X2 c231(
.A(net185),
.B(net180),
.ZN(net220)
);

MUX2_X1 c232(
.A(net93),
.B(net113),
.S(net172),
.Z(net221)
);

OAI21_X4 c233(
.A(net209),
.B1(net197),
.B2(net145),
.ZN(net222)
);

AND2_X4 c234(
.A1(net210),
.A2(net182),
.ZN(net223)
);

AND2_X1 c235(
.A1(net188),
.A2(net10641),
.ZN(net224)
);

INV_X1 c236(
.A(net176),
.ZN(net225)
);

INV_X2 c237(
.A(net212),
.ZN(net226)
);

NAND2_X1 c238(
.A1(net216),
.A2(net162),
.ZN(net227)
);

OAI222_X2 c239(
.A1(net171),
.A2(net227),
.B1(net219),
.B2(net88),
.C1(net191),
.C2(net157),
.ZN(net228)
);

SDFF_X1 c240(
.D(net219),
.SE(net204),
.SI(net209),
.CK(clk),
.Q(net230),
.QN(net229)
);

NAND2_X2 c241(
.A1(net200),
.A2(net11493),
.ZN(net231)
);

MUX2_X2 c242(
.A(net207),
.B(net219),
.S(net11492),
.Z(net232)
);

NAND3_X4 c243(
.A1(net206),
.A2(net10641),
.A3(net11493),
.ZN(net233)
);

INV_X8 c244(
.A(net10435),
.ZN(net234)
);

OR3_X4 c245(
.A1(net234),
.A2(net211),
.A3(net10642),
.ZN(net235)
);

SDFF_X2 c246(
.D(net234),
.SE(net233),
.SI(net11493),
.CK(clk),
.Q(net237),
.QN(net236)
);

AND3_X2 c247(
.A1(net160),
.A2(net233),
.A3(net11492),
.ZN(net238)
);

NOR3_X1 c248(
.A1(net174),
.A2(net234),
.A3(net188),
.ZN(net239)
);

INV_X16 c249(
.A(net159),
.ZN(net240)
);

INV_X32 c250(
.A(net67),
.ZN(net241)
);

INV_X4 c251(
.A(net251),
.ZN(net242)
);

INV_X1 c252(
.A(net184),
.ZN(net243)
);

INV_X2 c253(
.A(net239),
.ZN(net244)
);

INV_X8 c254(
.A(net97),
.ZN(net245)
);

NAND2_X4 c255(
.A1(net240),
.A2(net172),
.ZN(net246)
);

INV_X16 c256(
.A(net11320),
.ZN(net247)
);

INV_X32 c257(
.A(net9701),
.ZN(net248)
);

INV_X4 c258(
.A(net16),
.ZN(net249)
);

INV_X1 c259(
.A(net74),
.ZN(net250)
);

INV_X2 c260(
.A(net95),
.ZN(net251)
);

INV_X8 c261(
.A(net194),
.ZN(net252)
);

INV_X16 c262(
.A(net25),
.ZN(net253)
);

INV_X32 c263(
.A(net74),
.ZN(net254)
);

INV_X4 c264(
.A(net5),
.ZN(net255)
);

INV_X1 c265(
.A(net224),
.ZN(net256)
);

INV_X2 c266(
.A(net249),
.ZN(net257)
);

INV_X8 c267(
.A(net247),
.ZN(net258)
);

AND2_X2 c268(
.A1(net179),
.A2(net242),
.ZN(net259)
);

XOR2_X1 c269(
.A(net163),
.B(net194),
.Z(net260)
);

NOR2_X1 c270(
.A1(net95),
.A2(net203),
.ZN(net261)
);

INV_X16 c271(
.A(net193),
.ZN(net262)
);

INV_X32 c272(
.A(net239),
.ZN(net263)
);

INV_X4 c273(
.A(net260),
.ZN(net264)
);

OR2_X2 c274(
.A1(net264),
.A2(net243),
.ZN(net265)
);

INV_X1 c275(
.A(net225),
.ZN(net266)
);

INV_X2 c276(
.A(net264),
.ZN(net267)
);

INV_X8 c277(
.A(net260),
.ZN(net268)
);

INV_X16 c278(
.A(net9700),
.ZN(net269)
);

OR3_X2 c279(
.A1(net261),
.A2(net256),
.A3(net269),
.ZN(net270)
);

OAI21_X2 c280(
.A(net265),
.B1(net241),
.B2(net268),
.ZN(net271)
);

NOR2_X4 c281(
.A1(net262),
.A2(net225),
.ZN(net272)
);

INV_X32 c282(
.A(net251),
.ZN(net273)
);

OAI21_X1 c283(
.A(net270),
.B1(net244),
.B2(net231),
.ZN(net274)
);

NOR2_X2 c284(
.A1(net273),
.A2(net250),
.ZN(net275)
);

XOR2_X2 c285(
.A(net203),
.B(net172),
.Z(net276)
);

XNOR2_X1 c286(
.A(net252),
.B(net179),
.ZN(net277)
);

INV_X4 c287(
.A(net245),
.ZN(net278)
);

INV_X1 c288(
.A(net243),
.ZN(net279)
);

INV_X2 c289(
.A(net10084),
.ZN(net280)
);

INV_X8 c290(
.A(net11206),
.ZN(net281)
);

INV_X16 c291(
.A(net10832),
.ZN(net282)
);

INV_X32 c292(
.A(net11017),
.ZN(net283)
);

AOI21_X2 c293(
.A(net256),
.B1(net272),
.B2(net185),
.ZN(net284)
);

OR2_X4 c294(
.A1(net263),
.A2(net147),
.ZN(net285)
);

INV_X4 c295(
.A(net172),
.ZN(net286)
);

DFFRS_X1 c296(
.D(net282),
.RN(net277),
.SN(net284),
.CK(clk),
.Q(net288),
.QN(net287)
);

OAI221_X2 c297(
.A(net279),
.B1(net224),
.B2(net184),
.C1(net258),
.C2(net283),
.ZN(net289)
);

INV_X1 c298(
.A(net286),
.ZN(net290)
);

INV_X2 c299(
.A(net289),
.ZN(net291)
);

AOI21_X1 c300(
.A(net159),
.B1(net271),
.B2(net247),
.ZN(net292)
);

OR2_X1 c301(
.A1(net278),
.A2(net242),
.ZN(net293)
);

DFFRS_X2 c302(
.D(net242),
.RN(net293),
.SN(net279),
.CK(clk),
.Q(net295),
.QN(net294)
);

XNOR2_X2 c303(
.A(net267),
.B(net277),
.ZN(net296)
);

AND2_X4 c304(
.A1(net248),
.A2(net287),
.ZN(net297)
);

INV_X8 c305(
.A(net280),
.ZN(net298)
);

INV_X16 c306(
.A(net10327),
.ZN(net299)
);

AND2_X1 c307(
.A1(net295),
.A2(net157),
.ZN(net300)
);

AOI21_X4 c308(
.A(net250),
.B1(net298),
.B2(net269),
.ZN(net301)
);

AND3_X1 c309(
.A1(net301),
.A2(net300),
.A3(net279),
.ZN(net302)
);

NAND2_X1 c310(
.A1(net246),
.A2(net225),
.ZN(net303)
);

NAND3_X1 c311(
.A1(net224),
.A2(net275),
.A3(net67),
.ZN(net304)
);

INV_X32 c312(
.A(net11170),
.ZN(net305)
);

NOR3_X4 c313(
.A1(net269),
.A2(net298),
.A3(net11362),
.ZN(net306)
);

NAND2_X2 c314(
.A1(net306),
.A2(net277),
.ZN(net307)
);

NOR3_X2 c315(
.A1(net300),
.A2(net283),
.A3(net11053),
.ZN(net308)
);

NAND2_X4 c316(
.A1(net244),
.A2(net265),
.ZN(net309)
);

INV_X4 c317(
.A(net11003),
.ZN(net310)
);

AND3_X4 c318(
.A1(net300),
.A2(net310),
.A3(net258),
.ZN(net311)
);

SDFF_X1 c319(
.D(net309),
.SE(net299),
.SI(net185),
.CK(clk),
.Q(net313),
.QN(net312)
);

INV_X1 c320(
.A(net298),
.ZN(net314)
);

AND2_X2 c321(
.A1(net314),
.A2(net264),
.ZN(net315)
);

NAND3_X2 c322(
.A1(net297),
.A2(net307),
.A3(net263),
.ZN(net316)
);

SDFFR_X1 c323(
.D(net247),
.RN(net298),
.SE(net316),
.SI(net284),
.CK(clk),
.Q(net318),
.QN(net317)
);

AOI222_X1 c324(
.A1(net311),
.A2(net318),
.B1(net316),
.B2(net272),
.C1(net258),
.C2(net11362),
.ZN(net319)
);

SDFF_X2 c325(
.D(net231),
.SE(net284),
.SI(net11053),
.CK(clk),
.Q(net321),
.QN(net320)
);

DFFRS_X1 c326(
.D(net271),
.RN(net300),
.SN(net306),
.CK(clk),
.Q(net323),
.QN(net322)
);

INV_X2 c327(
.A(net11048),
.ZN(net324)
);

XOR2_X1 c328(
.A(net307),
.B(net310),
.Z(net325)
);

OR3_X1 c329(
.A1(net325),
.A2(net316),
.ZN(net10531)
);

SDFFRS_X1 c330(
.D(net291),
.RN(net297),
.SE(net197),
.SI(net325),
.SN(net10530),
.CK(clk),
.Q(net328),
.QN(net327)
);

AOI221_X4 c331(
.A(net324),
.B1(net193),
.B2(net327),
.C1(net172),
.C2(net10531),
.ZN(net329)
);

INV_X8 c332(
.A(net310),
.ZN(net330)
);

NOR2_X1 c333(
.A1(net137),
.A2(net290),
.ZN(net331)
);

INV_X16 c334(
.A(net165),
.ZN(net332)
);

INV_X32 c335(
.A(net165),
.ZN(net333)
);

OR2_X2 c336(
.A1(net237),
.A2(net157),
.ZN(net334)
);

NOR2_X4 c337(
.A1(net137),
.A2(net289),
.ZN(net335)
);

INV_X4 c338(
.A(net191),
.ZN(net336)
);

INV_X1 c339(
.A(net127),
.ZN(net337)
);

INV_X2 c340(
.A(net11237),
.ZN(net338)
);

INV_X8 c341(
.A(net11406),
.ZN(net339)
);

INV_X16 c342(
.A(net305),
.ZN(net340)
);

INV_X32 c343(
.A(net289),
.ZN(net341)
);

INV_X4 c344(
.A(net270),
.ZN(net342)
);

INV_X1 c345(
.A(net329),
.ZN(net343)
);

INV_X2 c346(
.A(net288),
.ZN(net344)
);

INV_X8 c347(
.A(net10417),
.ZN(net345)
);

INV_X16 c348(
.A(net323),
.ZN(net346)
);

INV_X32 c349(
.A(net320),
.ZN(net347)
);

INV_X4 c350(
.A(net340),
.ZN(net348)
);

INV_X1 c351(
.A(net269),
.ZN(net349)
);

INV_X2 c352(
.A(net272),
.ZN(net350)
);

NOR2_X2 c353(
.A1(net288),
.A2(net281),
.ZN(net351)
);

INV_X8 c354(
.A(net339),
.ZN(net352)
);

XOR2_X2 c355(
.A(net352),
.B(net345),
.Z(net353)
);

INV_X16 c356(
.A(net227),
.ZN(net354)
);

INV_X32 c357(
.A(net199),
.ZN(net355)
);

INV_X4 c358(
.A(in11),
.ZN(net356)
);

XNOR2_X1 c359(
.A(net356),
.B(net157),
.ZN(net357)
);

OR2_X4 c360(
.A1(net351),
.A2(in11),
.ZN(net358)
);

INV_X1 c361(
.A(net353),
.ZN(net359)
);

OR2_X1 c362(
.A1(net321),
.A2(net185),
.ZN(net360)
);

XNOR2_X2 c363(
.A(net356),
.B(net344),
.ZN(net361)
);

INV_X2 c364(
.A(net11406),
.ZN(net362)
);

AND2_X4 c365(
.A1(net240),
.A2(net355),
.ZN(net363)
);

AND2_X1 c366(
.A1(net348),
.A2(net333),
.ZN(net364)
);

INV_X8 c367(
.A(net363),
.ZN(net365)
);

INV_X16 c368(
.A(net9870),
.ZN(net366)
);

NAND2_X1 c369(
.A1(net362),
.A2(net335),
.ZN(net367)
);

NAND2_X2 c370(
.A1(net364),
.A2(net272),
.ZN(net368)
);

INV_X32 c371(
.A(net339),
.ZN(net369)
);

NAND2_X4 c372(
.A1(net223),
.A2(net358),
.ZN(net370)
);

INV_X4 c373(
.A(net281),
.ZN(net371)
);

MUX2_X1 c374(
.A(net336),
.B(net305),
.S(net330),
.Z(net372)
);

INV_X1 c375(
.A(net335),
.ZN(net373)
);

AND2_X2 c376(
.A1(net347),
.A2(net366),
.ZN(net374)
);

XOR2_X1 c377(
.A(net359),
.B(net363),
.Z(net375)
);

NOR2_X1 c378(
.A1(net366),
.A2(net363),
.ZN(net376)
);

INV_X2 c379(
.A(net10965),
.ZN(net377)
);

INV_X8 c380(
.A(net332),
.ZN(net378)
);

OR2_X2 c381(
.A1(net369),
.A2(net332),
.ZN(net379)
);

NOR2_X4 c382(
.A1(net365),
.A2(net362),
.ZN(net380)
);

NOR2_X2 c383(
.A1(net379),
.A2(net373),
.ZN(net381)
);

INV_X16 c384(
.A(net363),
.ZN(net382)
);

INV_X32 c385(
.A(net380),
.ZN(net383)
);

XOR2_X2 c386(
.A(net333),
.B(net377),
.Z(net384)
);

OAI21_X4 c387(
.A(net381),
.B1(net281),
.B2(net351),
.ZN(net385)
);

XNOR2_X1 c388(
.A(net368),
.B(net322),
.ZN(net386)
);

INV_X4 c389(
.A(net341),
.ZN(net387)
);

INV_X1 c390(
.A(net353),
.ZN(net388)
);

OR2_X4 c391(
.A1(net343),
.A2(net331),
.ZN(net389)
);

OR2_X1 c392(
.A1(net387),
.A2(net350),
.ZN(net390)
);

XNOR2_X2 c393(
.A(net355),
.B(net390),
.ZN(net391)
);

AND2_X4 c394(
.A1(net383),
.A2(net358),
.ZN(net392)
);

MUX2_X2 c395(
.A(net340),
.B(net386),
.S(net191),
.Z(net393)
);

NAND3_X4 c396(
.A1(net379),
.A2(net388),
.A3(net346),
.ZN(net394)
);

AND2_X1 c397(
.A1(net385),
.A2(net371),
.ZN(net395)
);

NAND2_X1 c398(
.A1(net391),
.A2(net338),
.ZN(net396)
);

NAND2_X2 c399(
.A1(net371),
.A2(net394),
.ZN(net397)
);

NAND2_X4 c400(
.A1(net367),
.A2(net10587),
.ZN(net398)
);

OR3_X4 c401(
.A1(net373),
.A2(net365),
.A3(net10587),
.ZN(net399)
);

DFFRS_X2 c402(
.D(net354),
.RN(net384),
.SN(net364),
.CK(clk),
.Q(net401),
.QN(net400)
);

AND3_X2 c403(
.A1(net382),
.A2(net389),
.A3(net392),
.ZN(net402)
);

AND2_X2 c404(
.A1(net381),
.A2(net10588),
.ZN(net403)
);

XOR2_X1 c405(
.A(net402),
.B(net351),
.Z(net404)
);

NOR2_X1 c406(
.A1(net394),
.A2(net403),
.ZN(net405)
);

NOR3_X1 c407(
.A1(net397),
.A2(net333),
.A3(net10588),
.ZN(net406)
);

INV_X2 c408(
.A(net11055),
.ZN(net407)
);

SDFF_X1 c409(
.D(net388),
.SE(net403),
.SI(net407),
.CK(clk),
.Q(net409),
.QN(net408)
);

OR4_X4 c410(
.A1(net407),
.A2(net383),
.A3(net409),
.A4(net404),
.ZN(net410)
);

SDFFR_X2 c411(
.D(net376),
.RN(net410),
.SE(net398),
.SI(net407),
.CK(clk),
.Q(net412),
.QN(net411)
);

OAI22_X2 c412(
.A1(net374),
.A2(net403),
.B1(net404),
.B2(net410),
.ZN(net413)
);

OR3_X2 c413(
.A1(net389),
.A2(net374),
.A3(net10944),
.ZN(net414)
);

OAI211_X4 c414(
.A(net386),
.B(net394),
.C1(net404),
.C2(net407),
.ZN(net415)
);

INV_X8 c415(
.A(net308),
.ZN(net416)
);

INV_X16 c416(
.A(net390),
.ZN(net417)
);

INV_X32 c417(
.A(net416),
.ZN(net418)
);

INV_X4 c418(
.A(net9915),
.ZN(net419)
);

OR2_X2 c419(
.A1(net380),
.A2(net399),
.ZN(net420)
);

OAI21_X2 c420(
.A(net404),
.B1(net416),
.B2(net349),
.ZN(net421)
);

INV_X1 c421(
.A(net418),
.ZN(net422)
);

NOR2_X4 c422(
.A1(net412),
.A2(net392),
.ZN(net423)
);

INV_X2 c423(
.A(net422),
.ZN(net424)
);

INV_X8 c424(
.A(net331),
.ZN(net425)
);

NOR2_X2 c425(
.A1(net147),
.A2(net153),
.ZN(net426)
);

INV_X16 c426(
.A(net331),
.ZN(net427)
);

INV_X32 c427(
.A(net390),
.ZN(net428)
);

XOR2_X2 c428(
.A(net427),
.B(net372),
.Z(net429)
);

OAI211_X1 c429(
.A(net411),
.B(net424),
.C1(net302),
.C2(net345),
.ZN(net430)
);

XNOR2_X1 c430(
.A(net336),
.B(net328),
.ZN(net431)
);

INV_X4 c431(
.A(net257),
.ZN(net432)
);

OR2_X4 c432(
.A1(net414),
.A2(net310),
.ZN(net433)
);

INV_X1 c433(
.A(net432),
.ZN(net434)
);

INV_X2 c434(
.A(net302),
.ZN(net435)
);

INV_X8 c435(
.A(net343),
.ZN(net436)
);

INV_X16 c436(
.A(net33),
.ZN(net437)
);

INV_X32 c437(
.A(net436),
.ZN(net438)
);

INV_X4 c438(
.A(net9653),
.ZN(net439)
);

OR2_X1 c439(
.A1(net290),
.A2(net433),
.ZN(net440)
);

INV_X1 c440(
.A(net378),
.ZN(net441)
);

INV_X2 c441(
.A(net261),
.ZN(net442)
);

INV_X8 c442(
.A(net198),
.ZN(net443)
);

INV_X16 c443(
.A(net439),
.ZN(net444)
);

XNOR2_X2 c444(
.A(net168),
.B(net419),
.ZN(net445)
);

AND2_X4 c445(
.A1(net440),
.A2(net436),
.ZN(net446)
);

AND2_X1 c446(
.A1(net433),
.A2(net308),
.ZN(net447)
);

OAI21_X1 c447(
.A(net424),
.B1(net439),
.B2(net433),
.ZN(net448)
);

NAND2_X1 c448(
.A1(net437),
.A2(net442),
.ZN(net449)
);

INV_X32 c449(
.A(net438),
.ZN(net450)
);

NAND2_X2 c450(
.A1(net406),
.A2(net439),
.ZN(net451)
);

AOI21_X2 c451(
.A(net420),
.B1(net435),
.B2(net447),
.ZN(net452)
);

INV_X4 c452(
.A(net9652),
.ZN(net453)
);

INV_X1 c453(
.A(net10509),
.ZN(net454)
);

INV_X2 c454(
.A(net435),
.ZN(net455)
);

INV_X8 c455(
.A(net10510),
.ZN(net456)
);

NAND2_X4 c456(
.A1(net401),
.A2(net442),
.ZN(net457)
);

INV_X16 c457(
.A(net437),
.ZN(net458)
);

INV_X32 c458(
.A(net11385),
.ZN(net459)
);

INV_X4 c459(
.A(net9912),
.ZN(net460)
);

AOI21_X1 c460(
.A(net302),
.B1(net454),
.B2(net443),
.ZN(net461)
);

INV_X1 c461(
.A(net9912),
.ZN(net462)
);

AOI21_X4 c462(
.A(net329),
.B1(net448),
.B2(net450),
.ZN(net463)
);

AND2_X2 c463(
.A1(net453),
.A2(net308),
.ZN(net464)
);

INV_X2 c464(
.A(net463),
.ZN(net465)
);

INV_X8 c465(
.A(net10069),
.ZN(net466)
);

AND3_X1 c466(
.A1(net451),
.A2(net350),
.A3(net432),
.ZN(net467)
);

XOR2_X1 c467(
.A(net436),
.B(net450),
.Z(net468)
);

NOR2_X1 c468(
.A1(net67),
.A2(net430),
.ZN(net469)
);

OR2_X2 c469(
.A1(net420),
.A2(net442),
.ZN(net470)
);

NOR2_X4 c470(
.A1(net455),
.A2(net460),
.ZN(net471)
);

INV_X16 c471(
.A(net459),
.ZN(net472)
);

INV_X32 c472(
.A(net451),
.ZN(net473)
);

NOR2_X2 c473(
.A1(net471),
.A2(net261),
.ZN(net474)
);

NAND3_X1 c474(
.A1(net431),
.A2(net455),
.A3(net422),
.ZN(net475)
);

NOR3_X4 c475(
.A1(net419),
.A2(net329),
.A3(net456),
.ZN(net476)
);

XOR2_X2 c476(
.A(net427),
.B(net406),
.Z(net477)
);

SDFF_X2 c477(
.D(net458),
.SE(net438),
.SI(net400),
.CK(clk),
.Q(net479),
.QN(net478)
);

INV_X4 c478(
.A(net473),
.ZN(net480)
);

NOR3_X2 c479(
.A1(net480),
.A2(net471),
.A3(net478),
.ZN(net481)
);

AND3_X4 c480(
.A1(net423),
.A2(net369),
.A3(net10759),
.ZN(net482)
);

XNOR2_X1 c481(
.A(net446),
.B(net468),
.ZN(net483)
);

INV_X1 c482(
.A(net349),
.ZN(net484)
);

INV_X2 c483(
.A(net484),
.ZN(net485)
);

INV_X8 c484(
.A(net11015),
.ZN(net486)
);

OR2_X4 c485(
.A1(net485),
.A2(net11169),
.ZN(net487)
);

NAND3_X2 c486(
.A1(net477),
.A2(net485),
.A3(net11015),
.ZN(net488)
);

OR3_X1 c487(
.A1(net429),
.A2(net453),
.A3(net480),
.ZN(net489)
);

MUX2_X1 c488(
.A(net482),
.B(net427),
.S(net441),
.Z(net490)
);

OAI21_X4 c489(
.A(net454),
.B1(net357),
.B2(net446),
.ZN(net491)
);

DFFRS_X1 c490(
.D(net476),
.RN(net447),
.SN(net458),
.CK(clk),
.Q(net493),
.QN(net492)
);

MUX2_X2 c491(
.A(net492),
.B(net439),
.S(net11169),
.Z(net494)
);

SDFFRS_X2 c492(
.D(net490),
.RN(net447),
.SE(net488),
.SI(net410),
.SN(net483),
.CK(clk),
.Q(net496),
.QN(net495)
);

OR2_X1 c493(
.A1(net493),
.A2(net453),
.ZN(net497)
);

INV_X16 c494(
.A(net10260),
.ZN(net498)
);

DFFS_X2 c495(
.D(net475),
.SN(net434),
.CK(clk),
.Q(net500),
.QN(net499)
);

NAND3_X4 c496(
.A1(net498),
.A2(net497),
.A3(net401),
.ZN(net501)
);

OR3_X4 c497(
.A1(net501),
.A2(net497),
.A3(net488),
.ZN(net502)
);

INV_X32 c498(
.A(net9773),
.ZN(net503)
);

INV_X4 c499(
.A(net392),
.ZN(net504)
);

XNOR2_X2 c500(
.A(net496),
.B(net528),
.ZN(net505)
);

AND2_X4 c501(
.A1(net57),
.A2(net518),
.ZN(net506)
);

INV_X1 c502(
.A(net531),
.ZN(net507)
);

INV_X2 c503(
.A(net506),
.ZN(net508)
);

AND2_X1 c504(
.A1(net520),
.A2(net533),
.ZN(net509)
);

INV_X8 c505(
.A(net345),
.ZN(net510)
);

NAND2_X1 c506(
.A1(net509),
.A2(net502),
.ZN(net511)
);

INV_X16 c507(
.A(net520),
.ZN(net512)
);

NAND2_X2 c508(
.A1(net529),
.A2(net504),
.ZN(net513)
);

NAND2_X4 c509(
.A1(net513),
.A2(net532),
.ZN(net514)
);

INV_X32 c510(
.A(net11078),
.ZN(net515)
);

INV_X4 c511(
.A(net157),
.ZN(net516)
);

INV_X1 c512(
.A(net518),
.ZN(net517)
);

INV_X2 c513(
.A(net9772),
.ZN(net518)
);

AND2_X2 c514(
.A1(net473),
.A2(net258),
.ZN(net519)
);

INV_X8 c515(
.A(net157),
.ZN(net520)
);

INV_X16 c516(
.A(net494),
.ZN(net521)
);

INV_X32 c517(
.A(net464),
.ZN(net522)
);

INV_X4 c518(
.A(net398),
.ZN(net523)
);

INV_X1 c519(
.A(net328),
.ZN(net524)
);

INV_X2 c520(
.A(net519),
.ZN(net525)
);

INV_X8 c521(
.A(net467),
.ZN(net526)
);

INV_X16 c522(
.A(net398),
.ZN(net527)
);

INV_X32 c523(
.A(net10024),
.ZN(net528)
);

XOR2_X1 c524(
.A(net453),
.B(net462),
.Z(net529)
);

INV_X4 c525(
.A(net399),
.ZN(net530)
);

INV_X1 c526(
.A(net477),
.ZN(net531)
);

INV_X2 c527(
.A(net345),
.ZN(net532)
);

DFFR_X1 c528(
.D(net360),
.RN(net525),
.CK(clk),
.Q(net534),
.QN(net533)
);

INV_X8 c529(
.A(net505),
.ZN(net535)
);

DFFRS_X2 c530(
.D(net360),
.RN(net399),
.SN(net362),
.CK(clk),
.Q(net537),
.QN(net536)
);

NOR2_X1 c531(
.A1(net531),
.A2(net532),
.ZN(net538)
);

OR2_X2 c532(
.A1(net440),
.A2(net33),
.ZN(net539)
);

NOR2_X4 c533(
.A1(net532),
.A2(net11368),
.ZN(net540)
);

NOR2_X2 c534(
.A1(net368),
.A2(net522),
.ZN(net541)
);

XOR2_X2 c535(
.A(net541),
.B(net517),
.Z(net542)
);

INV_X16 c536(
.A(net537),
.ZN(net543)
);

AND3_X2 c537(
.A1(net516),
.A2(net358),
.A3(net489),
.ZN(net544)
);

XNOR2_X1 c538(
.A(net540),
.B(net517),
.ZN(net545)
);

INV_X32 c539(
.A(net10473),
.ZN(net546)
);

NOR3_X1 c540(
.A1(net491),
.A2(net444),
.A3(net468),
.ZN(net547)
);

OR2_X4 c541(
.A1(net504),
.A2(net517),
.ZN(net548)
);

OR2_X1 c542(
.A1(net392),
.A2(net512),
.ZN(net549)
);

XNOR2_X2 c543(
.A(net453),
.B(net10683),
.ZN(net550)
);

AND2_X4 c544(
.A1(net469),
.A2(net536),
.ZN(net551)
);

AND2_X1 c545(
.A1(net546),
.A2(net540),
.ZN(net552)
);

NAND2_X1 c546(
.A1(net486),
.A2(net499),
.ZN(net553)
);

INV_X4 c547(
.A(net510),
.ZN(net554)
);

NAND2_X2 c548(
.A1(net549),
.A2(net508),
.ZN(net555)
);

NAND2_X4 c549(
.A1(net10682),
.A2(net11368),
.ZN(net556)
);

AND2_X2 c550(
.A1(net553),
.A2(net546),
.ZN(net557)
);

XOR2_X1 c551(
.A(net517),
.B(net543),
.Z(net558)
);

NOR2_X1 c552(
.A1(net558),
.A2(net555),
.ZN(net559)
);

OR2_X2 c553(
.A1(net555),
.A2(net553),
.ZN(net560)
);

NOR2_X4 c554(
.A1(net557),
.A2(net538),
.ZN(net561)
);

NOR2_X2 c555(
.A1(net549),
.A2(net556),
.ZN(net562)
);

XOR2_X2 c556(
.A(net552),
.B(net433),
.Z(net563)
);

SDFFRS_X1 c557(
.D(net515),
.RN(net529),
.SE(net198),
.SI(net559),
.SN(net466),
.CK(clk),
.Q(net565),
.QN(net564)
);

XNOR2_X1 c558(
.A(net532),
.B(net520),
.ZN(net566)
);

DFFR_X2 c559(
.D(net509),
.RN(net561),
.CK(clk),
.Q(net568),
.QN(net567)
);

AOI222_X4 c560(
.A1(net528),
.A2(net540),
.B1(net516),
.B2(net520),
.C1(net559),
.C2(net567),
.ZN(net569)
);

OR3_X2 c561(
.A1(net534),
.A2(net515),
.A3(net466),
.ZN(net570)
);

OR2_X4 c562(
.A1(net521),
.A2(net558),
.ZN(net571)
);

OR2_X1 c563(
.A1(net463),
.A2(net551),
.ZN(net572)
);

XNOR2_X2 c564(
.A(net505),
.B(net555),
.ZN(net573)
);

INV_X1 c565(
.A(net11078),
.ZN(net574)
);

OAI21_X2 c566(
.A(net571),
.B1(net557),
.B2(net570),
.ZN(net575)
);

AND2_X4 c567(
.A1(net542),
.A2(net535),
.ZN(net576)
);

DFFS_X1 c568(
.D(net573),
.SN(net574),
.CK(clk),
.Q(net578),
.QN(net577)
);

AND2_X1 c569(
.A1(net566),
.A2(net532),
.ZN(net579)
);

INV_X2 c570(
.A(net11424),
.ZN(net580)
);

NAND2_X1 c571(
.A1(net444),
.A2(net564),
.ZN(net581)
);

NAND2_X2 c572(
.A1(net539),
.A2(net11495),
.ZN(net582)
);

NAND2_X4 c573(
.A1(net575),
.A2(net581),
.ZN(net583)
);

OAI21_X1 c574(
.A(net565),
.B1(net583),
.B2(net11494),
.ZN(net584)
);

AND2_X2 c575(
.A1(net341),
.A2(net577),
.ZN(net585)
);

INV_X8 c576(
.A(net11380),
.ZN(net586)
);

SDFF_X1 c577(
.D(net502),
.SE(net573),
.SI(net586),
.CK(clk),
.Q(net588),
.QN(net587)
);

AOI21_X2 c578(
.A(net550),
.B1(net486),
.B2(net583),
.ZN(net589)
);

OAI33_X1 c579(
.A1(net580),
.A2(net494),
.A3(net589),
.B1(net586),
.B2(net559),
.B3(net11044),
.ZN(net590)
);

AOI222_X2 c580(
.A1(net503),
.A2(net582),
.B1(net587),
.B2(net517),
.C1(net586),
.C2(net11497),
.ZN(net591)
);

INV_X16 c581(
.A(net519),
.ZN(net592)
);

INV_X32 c582(
.A(net447),
.ZN(net593)
);

INV_X4 c583(
.A(net10097),
.ZN(net594)
);

INV_X1 c584(
.A(net500),
.ZN(net595)
);

INV_X2 c585(
.A(net375),
.ZN(net596)
);

XOR2_X1 c586(
.A(net585),
.B(net563),
.Z(net597)
);

INV_X8 c587(
.A(net9668),
.ZN(net598)
);

NOR2_X1 c588(
.A1(net570),
.A2(net448),
.ZN(net599)
);

INV_X16 c589(
.A(net574),
.ZN(net600)
);

INV_X32 c590(
.A(net510),
.ZN(net601)
);

OR2_X2 c591(
.A1(net554),
.A2(net361),
.ZN(net602)
);

INV_X4 c592(
.A(net86),
.ZN(net603)
);

NOR2_X4 c593(
.A1(net512),
.A2(net554),
.ZN(net604)
);

INV_X1 c594(
.A(net78),
.ZN(net605)
);

NOR2_X2 c595(
.A1(net563),
.A2(net594),
.ZN(net606)
);

XOR2_X2 c596(
.A(net443),
.B(net588),
.Z(net607)
);

INV_X2 c597(
.A(net468),
.ZN(net608)
);

INV_X8 c598(
.A(net361),
.ZN(net609)
);

INV_X16 c599(
.A(net556),
.ZN(net610)
);

INV_X32 c600(
.A(net604),
.ZN(net611)
);

INV_X4 c601(
.A(net594),
.ZN(net612)
);

INV_X1 c602(
.A(net9667),
.ZN(net613)
);

INV_X2 c603(
.A(net512),
.ZN(net614)
);

INV_X8 c604(
.A(net600),
.ZN(net615)
);

INV_X16 c605(
.A(net605),
.ZN(net616)
);

AOI21_X1 c606(
.A(net433),
.B1(net606),
.B2(net609),
.ZN(net617)
);

XNOR2_X1 c607(
.A(net468),
.B(net594),
.ZN(net618)
);

INV_X32 c608(
.A(net500),
.ZN(net619)
);

OR2_X4 c609(
.A1(net611),
.A2(net594),
.ZN(net620)
);

INV_X4 c610(
.A(net609),
.ZN(net621)
);

INV_X1 c611(
.A(net616),
.ZN(net622)
);

INV_X2 c612(
.A(net588),
.ZN(net623)
);

INV_X8 c613(
.A(net9855),
.ZN(net624)
);

INV_X16 c614(
.A(net621),
.ZN(net625)
);

OR2_X1 c615(
.A1(net611),
.A2(net601),
.ZN(net626)
);

XNOR2_X2 c616(
.A(net601),
.B(net581),
.ZN(net627)
);

AND2_X4 c617(
.A1(net615),
.A2(net543),
.ZN(net628)
);

AND2_X1 c618(
.A1(net610),
.A2(net615),
.ZN(net629)
);

NAND2_X1 c619(
.A1(net612),
.A2(net629),
.ZN(net630)
);

INV_X32 c620(
.A(net545),
.ZN(net631)
);

AOI21_X4 c621(
.A(net618),
.B1(net622),
.B2(net609),
.ZN(net632)
);

INV_X4 c622(
.A(net629),
.ZN(net633)
);

NAND2_X2 c623(
.A1(net599),
.A2(net615),
.ZN(net634)
);

INV_X1 c624(
.A(net9889),
.ZN(net635)
);

NAND2_X4 c625(
.A1(net633),
.A2(net361),
.ZN(net636)
);

DFFS_X2 c626(
.D(net607),
.SN(net510),
.CK(clk),
.Q(net638),
.QN(net637)
);

INV_X2 c627(
.A(net593),
.ZN(net639)
);

AND2_X2 c628(
.A1(net608),
.A2(net602),
.ZN(net640)
);

INV_X8 c629(
.A(net615),
.ZN(net641)
);

INV_X16 c630(
.A(net638),
.ZN(net642)
);

XOR2_X1 c631(
.A(net598),
.B(net589),
.Z(net643)
);

AND3_X1 c632(
.A1(net627),
.A2(net568),
.A3(net595),
.ZN(net644)
);

NOR2_X1 c633(
.A1(net448),
.A2(net610),
.ZN(net645)
);

DFFR_X1 c634(
.D(net636),
.RN(net634),
.CK(clk),
.Q(net647),
.QN(net646)
);

INV_X32 c635(
.A(net603),
.ZN(net648)
);

INV_X4 c636(
.A(net9914),
.ZN(net649)
);

NAND3_X1 c637(
.A1(net648),
.A2(net601),
.A3(net634),
.ZN(net650)
);

INV_X1 c638(
.A(net630),
.ZN(net651)
);

INV_X2 c639(
.A(net622),
.ZN(net652)
);

INV_X8 c640(
.A(net10324),
.ZN(net653)
);

INV_X16 c641(
.A(net625),
.ZN(net654)
);

OR2_X2 c642(
.A1(net631),
.A2(net624),
.ZN(net655)
);

NOR2_X4 c643(
.A1(net641),
.A2(net636),
.ZN(net656)
);

NOR3_X4 c644(
.A1(net570),
.A2(net649),
.A3(net641),
.ZN(net657)
);

NOR2_X2 c645(
.A1(net656),
.A2(net632),
.ZN(net658)
);

DFFR_X2 c646(
.D(net625),
.RN(net640),
.CK(clk),
.Q(net660),
.QN(net659)
);

DFFS_X1 c647(
.D(net632),
.SN(net441),
.CK(clk),
.Q(net662),
.QN(net661)
);

XOR2_X2 c648(
.A(net503),
.B(net649),
.Z(net663)
);

DFFS_X2 c649(
.D(net639),
.SN(net635),
.CK(clk),
.Q(net665),
.QN(net664)
);

INV_X32 c650(
.A(net624),
.ZN(net666)
);

NOR3_X2 c651(
.A1(net596),
.A2(net593),
.A3(net375),
.ZN(net667)
);

SDFF_X2 c652(
.D(net667),
.SE(net636),
.SI(net11018),
.CK(clk),
.Q(net669),
.QN(net668)
);

INV_X4 c653(
.A(net663),
.ZN(net670)
);

AND3_X4 c654(
.A1(net670),
.A2(net664),
.A3(net640),
.ZN(net671)
);

INV_X1 c655(
.A(net653),
.ZN(net672)
);

XNOR2_X1 c656(
.A(net651),
.B(net661),
.ZN(net673)
);

NAND3_X2 c657(
.A1(net641),
.A2(net670),
.A3(net673),
.ZN(net674)
);

OR3_X1 c658(
.A1(net443),
.A2(net545),
.A3(net636),
.ZN(net675)
);

AOI221_X2 c659(
.A(net198),
.B1(net667),
.B2(net603),
.C1(net602),
.C2(net615),
.ZN(net676)
);

MUX2_X1 c660(
.A(net597),
.B(net644),
.S(net570),
.Z(net677)
);

DFFRS_X1 c661(
.D(net594),
.RN(net674),
.SN(net617),
.CK(clk),
.Q(net679),
.QN(net678)
);

OAI21_X4 c662(
.A(net358),
.B1(net673),
.B2(net645),
.ZN(net680)
);

NOR4_X4 c663(
.A1(net644),
.A2(net669),
.A3(net666),
.A4(net678),
.ZN(net681)
);

INV_X2 c664(
.A(net11445),
.ZN(net682)
);

INV_X8 c665(
.A(net11497),
.ZN(net683)
);

INV_X16 c666(
.A(net619),
.ZN(net684)
);

OR2_X4 c667(
.A1(net258),
.A2(net660),
.ZN(net685)
);

INV_X32 c668(
.A(net683),
.ZN(net686)
);

INV_X4 c669(
.A(net472),
.ZN(net687)
);

INV_X1 c670(
.A(net657),
.ZN(net688)
);

INV_X2 c671(
.A(net10259),
.ZN(net689)
);

INV_X8 c672(
.A(net685),
.ZN(net690)
);

INV_X16 c673(
.A(net11445),
.ZN(net691)
);

INV_X32 c674(
.A(net619),
.ZN(net692)
);

INV_X4 c675(
.A(net9849),
.ZN(net693)
);

OR2_X1 c676(
.A1(net649),
.A2(net668),
.ZN(net694)
);

INV_X1 c677(
.A(net620),
.ZN(net695)
);

INV_X2 c678(
.A(net11178),
.ZN(net696)
);

INV_X8 c679(
.A(net688),
.ZN(net697)
);

XNOR2_X2 c680(
.A(net670),
.B(net595),
.ZN(net698)
);

INV_X16 c681(
.A(net648),
.ZN(net699)
);

INV_X32 c682(
.A(net372),
.ZN(net700)
);

INV_X4 c683(
.A(net649),
.ZN(net701)
);

INV_X1 c684(
.A(net9918),
.ZN(net702)
);

INV_X2 c685(
.A(net663),
.ZN(net703)
);

AND2_X4 c686(
.A1(net620),
.A2(net11178),
.ZN(net704)
);

INV_X8 c687(
.A(net704),
.ZN(net705)
);

INV_X16 c688(
.A(net683),
.ZN(net706)
);

AND2_X1 c689(
.A1(net654),
.A2(net595),
.ZN(net707)
);

INV_X32 c690(
.A(net595),
.ZN(net708)
);

INV_X4 c691(
.A(net703),
.ZN(net709)
);

INV_X1 c692(
.A(net690),
.ZN(net710)
);

INV_X2 c693(
.A(net532),
.ZN(net711)
);

NAND2_X1 c694(
.A1(net679),
.A2(net684),
.ZN(net712)
);

INV_X8 c695(
.A(net708),
.ZN(net713)
);

INV_X16 c696(
.A(net673),
.ZN(net714)
);

INV_X32 c697(
.A(net704),
.ZN(net715)
);

INV_X4 c698(
.A(net694),
.ZN(net716)
);

INV_X1 c699(
.A(net713),
.ZN(net717)
);

NAND2_X2 c700(
.A1(net689),
.A2(net703),
.ZN(net718)
);

INV_X2 c701(
.A(net702),
.ZN(net719)
);

INV_X8 c702(
.A(net9918),
.ZN(net720)
);

NAND2_X4 c703(
.A1(net709),
.A2(net690),
.ZN(net721)
);

AND2_X2 c704(
.A1(net718),
.A2(net703),
.ZN(net722)
);

INV_X16 c705(
.A(net599),
.ZN(net723)
);

INV_X32 c706(
.A(net699),
.ZN(net724)
);

XOR2_X1 c707(
.A(net717),
.B(net714),
.Z(net725)
);

NOR2_X1 c708(
.A1(net724),
.A2(net686),
.ZN(net726)
);

AOI221_X1 c709(
.A(net669),
.B1(net679),
.B2(net701),
.C1(net720),
.C2(net11496),
.ZN(net727)
);

INV_X4 c710(
.A(net10411),
.ZN(net728)
);

OR2_X2 c711(
.A1(net692),
.A2(net666),
.ZN(net729)
);

INV_X1 c712(
.A(net728),
.ZN(net730)
);

INV_X2 c713(
.A(net718),
.ZN(net731)
);

NOR2_X4 c714(
.A1(net697),
.A2(net721),
.ZN(net732)
);

MUX2_X2 c715(
.A(net730),
.B(net691),
.S(net704),
.Z(net733)
);

NOR2_X2 c716(
.A1(net732),
.A2(net602),
.ZN(net734)
);

XOR2_X2 c717(
.A(net733),
.B(net726),
.Z(net735)
);

INV_X8 c718(
.A(net716),
.ZN(net736)
);

INV_X16 c719(
.A(net727),
.ZN(net737)
);

XNOR2_X1 c720(
.A(net723),
.B(net685),
.ZN(net738)
);

INV_X32 c721(
.A(net687),
.ZN(net739)
);

OR2_X4 c722(
.A1(net712),
.A2(net734),
.ZN(net740)
);

NAND3_X4 c723(
.A1(net441),
.A2(net719),
.A3(net708),
.ZN(net741)
);

OR3_X4 c724(
.A1(net361),
.A2(net729),
.A3(net11498),
.ZN(net742)
);

INV_X4 c725(
.A(net710),
.ZN(net743)
);

AND3_X2 c726(
.A1(net726),
.A2(net628),
.A3(net734),
.ZN(net744)
);

DFFR_X1 c727(
.D(net735),
.RN(net744),
.CK(clk),
.Q(net746),
.QN(net745)
);

SDFFRS_X2 c728(
.D(net635),
.RN(net592),
.SE(net595),
.SI(net722),
.SN(net720),
.CK(clk),
.Q(net748),
.QN(net747)
);

NOR3_X1 c729(
.A1(net729),
.A2(net711),
.A3(net695),
.ZN(net749)
);

INV_X1 c730(
.A(net10248),
.ZN(net750)
);

INV_X2 c731(
.A(net749),
.ZN(net751)
);

OR2_X1 c732(
.A1(net700),
.A2(net742),
.ZN(net752)
);

XNOR2_X2 c733(
.A(net719),
.B(net750),
.ZN(net753)
);

OR3_X2 c734(
.A1(net576),
.A2(net748),
.A3(net686),
.ZN(net754)
);

AND2_X4 c735(
.A1(net684),
.A2(net739),
.ZN(net755)
);

INV_X8 c736(
.A(net725),
.ZN(net756)
);

INV_X16 c737(
.A(net755),
.ZN(net757)
);

INV_X32 c738(
.A(net753),
.ZN(net758)
);

AND2_X1 c739(
.A1(net741),
.A2(net584),
.ZN(net759)
);

OAI21_X2 c740(
.A(net742),
.B1(net759),
.B2(net11213),
.ZN(net760)
);

INV_X4 c741(
.A(net759),
.ZN(net761)
);

OAI21_X1 c742(
.A(net751),
.B1(net724),
.B2(net760),
.ZN(net762)
);

NOR4_X2 c743(
.A1(net761),
.A2(net716),
.A3(net762),
.A4(net727),
.ZN(net763)
);

OAI221_X1 c744(
.A(net754),
.B1(net747),
.B2(net761),
.C1(net699),
.C2(net666),
.ZN(net764)
);

OAI221_X4 c745(
.A(net740),
.B1(net763),
.B2(net756),
.C1(net762),
.C2(net742),
.ZN(net765)
);

NAND2_X1 c746(
.A1(net760),
.A2(net11213),
.ZN(net766)
);

NAND2_X2 c747(
.A1(net344),
.A2(net714),
.ZN(net767)
);

INV_X1 c748(
.A(net9966),
.ZN(net768)
);

INV_X2 c749(
.A(net731),
.ZN(net769)
);

INV_X8 c750(
.A(net666),
.ZN(net770)
);

NAND2_X4 c751(
.A1(net507),
.A2(net769),
.ZN(net771)
);

INV_X16 c752(
.A(net756),
.ZN(net772)
);

AND2_X2 c753(
.A1(net318),
.A2(net722),
.ZN(net773)
);

INV_X32 c754(
.A(net722),
.ZN(net774)
);

INV_X4 c755(
.A(net628),
.ZN(net775)
);

INV_X1 c756(
.A(net662),
.ZN(net776)
);

AOI21_X2 c757(
.A(net285),
.B1(net538),
.B2(net776),
.ZN(net777)
);

INV_X2 c758(
.A(net770),
.ZN(net778)
);

AOI21_X1 c759(
.A(net760),
.B1(net646),
.B2(net698),
.ZN(net779)
);

INV_X8 c760(
.A(net628),
.ZN(net780)
);

INV_X16 c761(
.A(net775),
.ZN(net781)
);

INV_X32 c762(
.A(net746),
.ZN(net782)
);

XOR2_X1 c763(
.A(net71),
.B(net770),
.Z(net783)
);

NOR2_X1 c764(
.A1(net769),
.A2(net720),
.ZN(net784)
);

INV_X4 c765(
.A(net623),
.ZN(net785)
);

INV_X1 c766(
.A(net785),
.ZN(net786)
);

INV_X2 c767(
.A(net11499),
.ZN(net787)
);

INV_X8 c768(
.A(net657),
.ZN(net788)
);

INV_X16 c769(
.A(net736),
.ZN(net789)
);

INV_X32 c770(
.A(net623),
.ZN(net790)
);

INV_X4 c771(
.A(net714),
.ZN(net791)
);

INV_X1 c772(
.A(net782),
.ZN(net792)
);

OR2_X2 c773(
.A1(net57),
.A2(net791),
.ZN(net793)
);

NOR2_X4 c774(
.A1(net780),
.A2(net788),
.ZN(net794)
);

INV_X2 c775(
.A(net776),
.ZN(net795)
);

INV_X8 c776(
.A(net743),
.ZN(net796)
);

INV_X16 c777(
.A(net787),
.ZN(net797)
);

NOR2_X2 c778(
.A1(net773),
.A2(net778),
.ZN(net798)
);

INV_X32 c779(
.A(net9770),
.ZN(net799)
);

XOR2_X2 c780(
.A(net647),
.B(net790),
.Z(net800)
);

XNOR2_X1 c781(
.A(net794),
.B(net731),
.ZN(net801)
);

INV_X4 c782(
.A(net791),
.ZN(net802)
);

OR2_X4 c783(
.A1(net796),
.A2(net797),
.ZN(net803)
);

INV_X1 c784(
.A(net790),
.ZN(net804)
);

AOI21_X4 c785(
.A(net802),
.B1(net793),
.B2(net731),
.ZN(net805)
);

INV_X2 c786(
.A(net786),
.ZN(net806)
);

OR2_X1 c787(
.A1(net647),
.A2(net744),
.ZN(net807)
);

XNOR2_X2 c788(
.A(net721),
.B(net799),
.ZN(net808)
);

AND2_X4 c789(
.A1(net801),
.A2(net10546),
.ZN(net809)
);

INV_X8 c790(
.A(net788),
.ZN(net810)
);

INV_X16 c791(
.A(net806),
.ZN(net811)
);

INV_X32 c792(
.A(net11469),
.ZN(net812)
);

INV_X4 c793(
.A(net800),
.ZN(net813)
);

AND2_X1 c794(
.A1(net786),
.A2(net772),
.ZN(net814)
);

NAND2_X1 c795(
.A1(net722),
.A2(net743),
.ZN(net815)
);

INV_X1 c796(
.A(net792),
.ZN(net816)
);

INV_X2 c797(
.A(net802),
.ZN(net817)
);

NAND2_X2 c798(
.A1(net768),
.A2(net790),
.ZN(net818)
);

INV_X8 c799(
.A(net11051),
.ZN(net819)
);

DFFR_X2 c800(
.D(net797),
.RN(net817),
.CK(clk),
.Q(net821),
.QN(net820)
);

INV_X16 c801(
.A(net9770),
.ZN(net822)
);

NAND2_X4 c802(
.A1(net801),
.A2(net806),
.ZN(net823)
);

INV_X32 c803(
.A(net767),
.ZN(net824)
);

AOI211_X4 c804(
.A(net809),
.B(net818),
.C1(net797),
.C2(net819),
.ZN(net825)
);

AND2_X2 c805(
.A1(net775),
.A2(net815),
.ZN(net826)
);

XOR2_X1 c806(
.A(net781),
.B(net657),
.Z(net827)
);

INV_X4 c807(
.A(net10547),
.ZN(net828)
);

INV_X1 c808(
.A(net804),
.ZN(net829)
);

NOR2_X1 c809(
.A1(net715),
.A2(net826),
.ZN(net830)
);

OR2_X2 c810(
.A1(net793),
.A2(net826),
.ZN(net831)
);

NOR4_X1 c811(
.A1(net796),
.A2(net819),
.A3(net793),
.A4(net825),
.ZN(net832)
);

OAI221_X2 c812(
.A(net818),
.B1(net825),
.B2(net657),
.C1(net790),
.C2(net823),
.ZN(net833)
);

NOR2_X4 c813(
.A1(net780),
.A2(net822),
.ZN(net834)
);

INV_X2 c814(
.A(net10021),
.ZN(net835)
);

NOR2_X2 c815(
.A1(net693),
.A2(net823),
.ZN(net836)
);

XOR2_X2 c816(
.A(net803),
.B(net829),
.Z(net837)
);

XNOR2_X1 c817(
.A(net837),
.B(net834),
.ZN(net838)
);

DFFS_X1 c818(
.D(net833),
.SN(net835),
.CK(clk),
.Q(net840),
.QN(net839)
);

OR2_X4 c819(
.A1(net829),
.A2(net714),
.ZN(net841)
);

DFFRS_X2 c820(
.D(net831),
.RN(net838),
.SN(net784),
.CK(clk),
.Q(net843),
.QN(net842)
);

AOI221_X4 c821(
.A(net838),
.B1(net816),
.B2(net802),
.C1(net825),
.C2(net837),
.ZN(net844)
);

AND3_X1 c822(
.A1(net811),
.A2(net826),
.A3(net839),
.ZN(net845)
);

SDFF_X1 c823(
.D(net844),
.SE(net813),
.SI(net804),
.CK(clk),
.Q(net847),
.QN(net846)
);

NAND3_X1 c824(
.A1(net847),
.A2(net666),
.A3(net799),
.ZN(net848)
);

AOI221_X2 c825(
.A(net830),
.B1(net842),
.B2(net845),
.C1(net778),
.C2(net839),
.ZN(net849)
);

AOI211_X2 c826(
.A(net832),
.B(net801),
.C1(net844),
.C2(net825),
.ZN(net850)
);

OR2_X1 c827(
.A1(net836),
.A2(net809),
.ZN(net851)
);

XNOR2_X2 c828(
.A(net841),
.B(net816),
.ZN(net852)
);

SDFFRS_X1 c829(
.D(net852),
.RN(net845),
.SE(net851),
.SI(net825),
.SN(net774),
.CK(clk),
.Q(net854),
.QN(net853)
);

INV_X8 c830(
.A(net825),
.ZN(net855)
);

INV_X16 c831(
.A(net9705),
.ZN(net856)
);

INV_X32 c832(
.A(net466),
.ZN(net857)
);

AND2_X4 c833(
.A1(net589),
.A2(net556),
.ZN(net858)
);

INV_X4 c834(
.A(net358),
.ZN(net859)
);

INV_X1 c835(
.A(net857),
.ZN(net860)
);

INV_X2 c836(
.A(net857),
.ZN(net861)
);

INV_X8 c837(
.A(net859),
.ZN(net862)
);

INV_X16 c838(
.A(net858),
.ZN(net863)
);

AND2_X1 c839(
.A1(net824),
.A2(net823),
.ZN(net864)
);

INV_X32 c840(
.A(net861),
.ZN(net865)
);

INV_X4 c841(
.A(net820),
.ZN(net866)
);

NAND2_X1 c842(
.A1(net866),
.A2(net864),
.ZN(net867)
);

INV_X1 c843(
.A(net10564),
.ZN(net868)
);

INV_X2 c844(
.A(net9706),
.ZN(net869)
);

INV_X8 c845(
.A(net827),
.ZN(net870)
);

NAND2_X2 c846(
.A1(net756),
.A2(net637),
.ZN(net871)
);

SDFF_X2 c847(
.D(net871),
.SE(net827),
.SI(net853),
.CK(clk),
.Q(net873),
.QN(net872)
);

INV_X16 c848(
.A(net859),
.ZN(net874)
);

INV_X32 c849(
.A(net762),
.ZN(net875)
);

DFFRS_X1 c850(
.D(net862),
.RN(net873),
.SN(net772),
.CK(clk),
.Q(net877),
.QN(net876)
);

INV_X4 c851(
.A(net789),
.ZN(net878)
);

NOR3_X4 c852(
.A1(net854),
.A2(net872),
.A3(net788),
.ZN(net879)
);

INV_X1 c853(
.A(net815),
.ZN(net880)
);

INV_X2 c854(
.A(net878),
.ZN(net881)
);

INV_X8 c855(
.A(net868),
.ZN(net882)
);

INV_X16 c856(
.A(net865),
.ZN(net883)
);

INV_X32 c857(
.A(net778),
.ZN(net884)
);

INV_X4 c858(
.A(net824),
.ZN(net885)
);

INV_X1 c859(
.A(net858),
.ZN(net886)
);

NAND2_X4 c860(
.A1(net706),
.A2(net778),
.ZN(net887)
);

AND2_X2 c861(
.A1(net731),
.A2(net779),
.ZN(net888)
);

XOR2_X1 c862(
.A(net868),
.B(net816),
.Z(net889)
);

NOR2_X1 c863(
.A1(net884),
.A2(net825),
.ZN(net890)
);

OR2_X2 c864(
.A1(net522),
.A2(net784),
.ZN(net891)
);

NOR2_X4 c865(
.A1(net889),
.A2(net784),
.ZN(net892)
);

INV_X2 c866(
.A(net883),
.ZN(net893)
);

INV_X8 c867(
.A(net9907),
.ZN(net894)
);

NOR3_X2 c868(
.A1(net860),
.A2(net893),
.A3(net749),
.ZN(net895)
);

AOI22_X1 c869(
.A1(net883),
.A2(net857),
.B1(net495),
.B2(net839),
.ZN(net896)
);

INV_X16 c870(
.A(net749),
.ZN(net897)
);

INV_X32 c871(
.A(net10337),
.ZN(net898)
);

NOR2_X2 c872(
.A1(net882),
.A2(net866),
.ZN(net899)
);

INV_X4 c873(
.A(net870),
.ZN(net900)
);

INV_X1 c874(
.A(net866),
.ZN(net901)
);

XOR2_X2 c875(
.A(net893),
.B(net900),
.Z(net902)
);

INV_X2 c876(
.A(net9907),
.ZN(net903)
);

INV_X8 c877(
.A(net896),
.ZN(net904)
);

AND3_X4 c878(
.A1(net878),
.A2(net900),
.A3(net883),
.ZN(net905)
);

DFFS_X2 c879(
.D(net890),
.SN(net903),
.CK(clk),
.Q(net907),
.QN(net906)
);

NAND3_X2 c880(
.A1(net559),
.A2(net840),
.A3(net637),
.ZN(net908)
);

INV_X16 c881(
.A(net897),
.ZN(net909)
);

INV_X32 c882(
.A(net898),
.ZN(net910)
);

XNOR2_X1 c883(
.A(net904),
.B(net891),
.ZN(net911)
);

OR2_X4 c884(
.A1(net886),
.A2(net854),
.ZN(net912)
);

OR2_X1 c885(
.A1(net910),
.A2(net882),
.ZN(net913)
);

XNOR2_X2 c886(
.A(net856),
.B(net815),
.ZN(net914)
);

INV_X4 c887(
.A(net874),
.ZN(net915)
);

AND2_X4 c888(
.A1(net881),
.A2(net789),
.ZN(net916)
);

INV_X1 c889(
.A(net916),
.ZN(net917)
);

INV_X2 c890(
.A(net869),
.ZN(net918)
);

OR3_X1 c891(
.A1(net880),
.A2(net823),
.A3(net911),
.ZN(net919)
);

MUX2_X1 c892(
.A(net825),
.B(net896),
.S(net883),
.Z(net920)
);

INV_X8 c893(
.A(net913),
.ZN(net921)
);

INV_X16 c894(
.A(net10563),
.ZN(net922)
);

INV_X32 c895(
.A(net9849),
.ZN(net923)
);

INV_X4 c896(
.A(net10258),
.ZN(net924)
);

OAI21_X4 c897(
.A(net919),
.B1(net900),
.B2(net788),
.ZN(net925)
);

AND2_X1 c898(
.A1(net788),
.A2(net891),
.ZN(net926)
);

MUX2_X2 c899(
.A(net873),
.B(net762),
.S(net11114),
.Z(net927)
);

NAND2_X1 c900(
.A1(net918),
.A2(net11114),
.ZN(net928)
);

INV_X1 c901(
.A(net10347),
.ZN(net929)
);

OAI222_X1 c902(
.A1(net923),
.A2(net925),
.B1(net893),
.B2(net900),
.C1(net889),
.C2(net878),
.ZN(net930)
);

NAND2_X2 c903(
.A1(net928),
.A2(net926),
.ZN(net931)
);

INV_X2 c904(
.A(net931),
.ZN(net932)
);

INV_X8 c905(
.A(net11318),
.ZN(net933)
);

NAND3_X4 c906(
.A1(net924),
.A2(net933),
.A3(net899),
.ZN(net934)
);

NAND2_X4 c907(
.A1(net895),
.A2(net816),
.ZN(net935)
);

OR3_X4 c908(
.A1(net929),
.A2(net932),
.A3(net922),
.ZN(net936)
);

AOI221_X1 c909(
.A(net902),
.B1(net877),
.B2(net934),
.C1(net889),
.C2(net559),
.ZN(net937)
);

DFFRS_X2 c910(
.D(net918),
.RN(net933),
.SN(net890),
.CK(clk),
.Q(net939),
.QN(net938)
);

AND3_X2 c911(
.A1(net899),
.A2(net917),
.A3(net10805),
.ZN(net940)
);

AND2_X2 c912(
.A1(net940),
.A2(net10773),
.ZN(net941)
);

INV_X16 c913(
.A(net35),
.ZN(net942)
);

INV_X32 c914(
.A(net9),
.ZN(net943)
);

INV_X4 c915(
.A(net50),
.ZN(net944)
);

INV_X1 c916(
.A(net26),
.ZN(net945)
);

INV_X2 c917(
.A(net47),
.ZN(net946)
);

INV_X8 c918(
.A(net6),
.ZN(net947)
);

INV_X16 c919(
.A(net46),
.ZN(net948)
);

INV_X32 c920(
.A(in23),
.ZN(net949)
);

INV_X4 c921(
.A(in5),
.ZN(net950)
);

INV_X1 c922(
.A(net19),
.ZN(net951)
);

INV_X2 c923(
.A(net6),
.ZN(net952)
);

XOR2_X1 c924(
.A(in12),
.B(net50),
.Z(net953)
);

INV_X8 c925(
.A(net946),
.ZN(net954)
);

INV_X16 c926(
.A(net9785),
.ZN(net955)
);

INV_X32 c927(
.A(net51),
.ZN(net956)
);

INV_X4 c928(
.A(net9785),
.ZN(net957)
);

NOR2_X1 c929(
.A1(in19),
.A2(net952),
.ZN(net958)
);

INV_X1 c930(
.A(net953),
.ZN(net959)
);

INV_X2 c931(
.A(in13),
.ZN(net960)
);

INV_X8 c932(
.A(net953),
.ZN(net961)
);

INV_X16 c933(
.A(net957),
.ZN(net962)
);

INV_X32 c934(
.A(in19),
.ZN(net963)
);

INV_X4 c935(
.A(net960),
.ZN(net964)
);

OR2_X2 c936(
.A1(net959),
.A2(net961),
.ZN(net965)
);

INV_X1 c937(
.A(net957),
.ZN(net966)
);

INV_X2 c938(
.A(net966),
.ZN(net967)
);

NOR2_X4 c939(
.A1(net19),
.A2(net958),
.ZN(net968)
);

INV_X8 c940(
.A(net46),
.ZN(net969)
);

INV_X16 c941(
.A(in7),
.ZN(net970)
);

INV_X32 c942(
.A(net951),
.ZN(net971)
);

INV_X4 c943(
.A(net971),
.ZN(net972)
);

INV_X1 c944(
.A(net950),
.ZN(net973)
);

INV_X2 c945(
.A(net49),
.ZN(net974)
);

INV_X8 c946(
.A(net974),
.ZN(net975)
);

NOR3_X1 c947(
.A1(net961),
.A2(net966),
.A3(net973),
.ZN(net976)
);

INV_X16 c948(
.A(net972),
.ZN(net977)
);

NOR2_X2 c949(
.A1(net51),
.A2(net963),
.ZN(net978)
);

INV_X32 c950(
.A(in9),
.ZN(net979)
);

INV_X4 c951(
.A(net958),
.ZN(net980)
);

INV_X1 c952(
.A(net50),
.ZN(net981)
);

INV_X2 c953(
.A(net979),
.ZN(net982)
);

XOR2_X2 c954(
.A(net945),
.B(net981),
.Z(net983)
);

XNOR2_X1 c955(
.A(net980),
.B(net983),
.ZN(net984)
);

INV_X8 c956(
.A(net975),
.ZN(net985)
);

OR2_X4 c957(
.A1(net976),
.A2(net982),
.ZN(net986)
);

OR2_X1 c958(
.A1(net951),
.A2(net971),
.ZN(net987)
);

OR3_X2 c959(
.A1(net959),
.A2(net974),
.A3(net976),
.ZN(net988)
);

XNOR2_X2 c960(
.A(net970),
.B(net964),
.ZN(net989)
);

INV_X16 c961(
.A(net977),
.ZN(net990)
);

OAI21_X2 c962(
.A(in15),
.B1(net6),
.B2(net949),
.ZN(net991)
);

INV_X32 c963(
.A(net989),
.ZN(net992)
);

AND2_X4 c964(
.A1(net988),
.A2(net6),
.ZN(net993)
);

INV_X4 c965(
.A(net978),
.ZN(net994)
);

AND2_X1 c966(
.A1(net987),
.A2(net977),
.ZN(net995)
);

NAND2_X1 c967(
.A1(net955),
.A2(net990),
.ZN(net996)
);

NAND2_X2 c968(
.A1(net952),
.A2(in23),
.ZN(net997)
);

NAND2_X4 c969(
.A1(net943),
.A2(net992),
.ZN(net998)
);

AND2_X2 c970(
.A1(net985),
.A2(net994),
.ZN(net999)
);

OAI21_X1 c971(
.A(net976),
.B1(net955),
.B2(net966),
.ZN(net1000)
);

XOR2_X1 c972(
.A(net946),
.B(net967),
.Z(net1001)
);

NOR2_X1 c973(
.A1(net998),
.A2(net989),
.ZN(net1002)
);

INV_X1 c974(
.A(net967),
.ZN(net1003)
);

INV_X2 c975(
.A(net997),
.ZN(net1004)
);

INV_X8 c976(
.A(net1002),
.ZN(net1005)
);

INV_X16 c977(
.A(in9),
.ZN(net1006)
);

AOI21_X2 c978(
.A(net1004),
.B1(net1005),
.B2(net970),
.ZN(net1007)
);

OR2_X2 c979(
.A1(net964),
.A2(net976),
.ZN(net1008)
);

INV_X32 c980(
.A(in12),
.ZN(net1009)
);

INV_X4 c981(
.A(net994),
.ZN(net1010)
);

NOR2_X4 c982(
.A1(net983),
.A2(net985),
.ZN(net1011)
);

NOR2_X2 c983(
.A1(net1010),
.A2(net1002),
.ZN(net1012)
);

XOR2_X2 c984(
.A(net1011),
.B(net1008),
.Z(net1013)
);

AOI21_X1 c985(
.A(net981),
.B1(net35),
.B2(net1001),
.ZN(net1014)
);

XNOR2_X1 c986(
.A(net992),
.B(net971),
.ZN(net1015)
);

OR2_X4 c987(
.A1(net1003),
.A2(net10625),
.ZN(net1016)
);

OAI222_X4 c988(
.A1(net1004),
.A2(net949),
.B1(net991),
.B2(net1016),
.C1(net973),
.C2(net10626),
.ZN(net1017)
);

OR2_X1 c989(
.A1(net948),
.A2(net10626),
.ZN(net1018)
);

OAI221_X1 c990(
.A(net1012),
.B1(net1017),
.B2(net973),
.C1(net949),
.C2(net10625),
.ZN(net1019)
);

DFFR_X1 c991(
.D(net1001),
.RN(net1015),
.CK(clk),
.Q(net1021),
.QN(net1020)
);

XNOR2_X2 c992(
.A(net1015),
.B(net979),
.ZN(net1022)
);

AND4_X4 c993(
.A1(net1017),
.A2(net1022),
.A3(net1012),
.A4(net1016),
.ZN(net1023)
);

NAND4_X1 c994(
.A1(net1022),
.A2(net1008),
.A3(net1012),
.A4(net966),
.ZN(net1024)
);

OR4_X1 c995(
.A1(net996),
.A2(net1000),
.A3(net1022),
.A4(net966),
.ZN(net1025)
);

AOI21_X4 c996(
.A(net1087),
.B1(net1085),
.B2(net954),
.ZN(net1026)
);

INV_X1 c997(
.A(net995),
.ZN(net1027)
);

AND2_X4 c998(
.A1(net1089),
.A2(net52),
.ZN(net1028)
);

AND2_X1 c999(
.A1(net110),
.A2(net990),
.ZN(net1029)
);

INV_X2 c1000(
.A(net1074),
.ZN(net1030)
);

INV_X8 c1001(
.A(net121),
.ZN(net1031)
);

NAND2_X1 c1002(
.A1(net1018),
.A2(net1091),
.ZN(net1032)
);

NAND2_X2 c1003(
.A1(net1088),
.A2(net1027),
.ZN(net1033)
);

INV_X16 c1004(
.A(net10705),
.ZN(net1034)
);

INV_X32 c1005(
.A(net1062),
.ZN(net1035)
);

INV_X4 c1006(
.A(net1030),
.ZN(net1036)
);

SDFF_X1 c1007(
.D(net1027),
.SE(net1031),
.SI(net1033),
.CK(clk),
.Q(net1038),
.QN(net1037)
);

INV_X1 c1008(
.A(net984),
.ZN(net1039)
);

INV_X2 c1009(
.A(net950),
.ZN(net1040)
);

AND3_X1 c1010(
.A1(net1034),
.A2(net987),
.A3(net1008),
.ZN(net1041)
);

NAND2_X4 c1011(
.A1(net1060),
.A2(net1072),
.ZN(net1042)
);

AND2_X2 c1012(
.A1(net1071),
.A2(net1082),
.ZN(net1043)
);

XOR2_X1 c1013(
.A(net1028),
.B(net1061),
.Z(net1044)
);

NOR2_X1 c1014(
.A1(net1078),
.A2(net1060),
.ZN(net1045)
);

INV_X8 c1015(
.A(net1083),
.ZN(net1046)
);

INV_X16 c1016(
.A(net1073),
.ZN(net1047)
);

OR2_X2 c1017(
.A1(net1046),
.A2(in25),
.ZN(net1048)
);

INV_X32 c1018(
.A(net10535),
.ZN(net1049)
);

SDFF_X2 c1019(
.D(net1031),
.SE(net138),
.SI(net962),
.CK(clk),
.Q(net1051),
.QN(net1050)
);

OAI222_X2 c1020(
.A1(net1049),
.A2(net1043),
.B1(net1075),
.B2(net1067),
.C1(net973),
.C2(net954),
.ZN(net1052)
);

INV_X4 c1021(
.A(net1081),
.ZN(net1053)
);

DFFR_X2 c1022(
.D(net1076),
.RN(net1091),
.CK(clk),
.Q(net1055),
.QN(net1054)
);

NOR2_X4 c1023(
.A1(net1059),
.A2(net11500),
.ZN(net1056)
);

NOR2_X2 c1024(
.A1(net100),
.A2(net996),
.ZN(net1057)
);

XOR2_X2 c1025(
.A(net1018),
.B(net144),
.Z(net1058)
);

XNOR2_X1 c1026(
.A(net133),
.B(net49),
.ZN(net1059)
);

OR2_X4 c1027(
.A1(net990),
.A2(net126),
.ZN(net1060)
);

OR2_X1 c1028(
.A1(net109),
.A2(net986),
.ZN(net1061)
);

NAND3_X1 c1029(
.A1(net52),
.A2(net144),
.A3(net17),
.ZN(net1062)
);

DFFRS_X1 c1030(
.D(net37),
.RN(net1062),
.SN(net110),
.CK(clk),
.Q(net1064),
.QN(net1063)
);

XNOR2_X2 c1031(
.A(net144),
.B(net141),
.ZN(net1065)
);

INV_X1 c1032(
.A(net9675),
.ZN(net1066)
);

INV_X2 c1033(
.A(net965),
.ZN(net1067)
);

DFFS_X1 c1034(
.D(net115),
.SN(net984),
.CK(clk),
.Q(net1069),
.QN(net1068)
);

AND2_X4 c1035(
.A1(net1063),
.A2(net52),
.ZN(net1070)
);

INV_X8 c1036(
.A(net62),
.ZN(net1071)
);

DFFS_X2 c1037(
.D(net1058),
.SN(net96),
.CK(clk),
.Q(net1073),
.QN(net1072)
);

AND2_X1 c1038(
.A1(net986),
.A2(net66),
.ZN(net1074)
);

DFFR_X1 c1039(
.D(net944),
.RN(net138),
.CK(clk),
.Q(net1076),
.QN(net1075)
);

INV_X16 c1040(
.A(net965),
.ZN(net1077)
);

INV_X32 c1041(
.A(net52),
.ZN(net1078)
);

INV_X4 c1042(
.A(net1077),
.ZN(net1079)
);

INV_X1 c1043(
.A(net1058),
.ZN(net1080)
);

INV_X2 c1044(
.A(net1061),
.ZN(net1081)
);

NAND2_X1 c1045(
.A1(net76),
.A2(net70),
.ZN(net1082)
);

INV_X8 c1046(
.A(net10058),
.ZN(net1083)
);

NAND2_X2 c1047(
.A1(net126),
.A2(net1079),
.ZN(net1084)
);

NAND2_X4 c1048(
.A1(net1082),
.A2(net995),
.ZN(net1085)
);

INV_X16 c1049(
.A(net1003),
.ZN(net1086)
);

INV_X32 c1050(
.A(net66),
.ZN(net1087)
);

INV_X4 c1051(
.A(net1079),
.ZN(net1088)
);

INV_X1 c1052(
.A(net973),
.ZN(net1089)
);

INV_X2 c1053(
.A(net1078),
.ZN(net1090)
);

AND2_X2 c1054(
.A1(net1084),
.A2(net1061),
.ZN(net1091)
);

INV_X8 c1055(
.A(net1085),
.ZN(net1092)
);

INV_X16 c1056(
.A(net141),
.ZN(net1093)
);

XOR2_X1 c1057(
.A(net1043),
.B(net141),
.Z(net1094)
);

DFFR_X2 c1058(
.D(net1036),
.RN(net966),
.CK(clk),
.Q(net1096),
.QN(net1095)
);

INV_X32 c1059(
.A(net9676),
.ZN(net1097)
);

NOR3_X4 c1060(
.A1(net1053),
.A2(net1009),
.A3(net1096),
.ZN(net1098)
);

NOR2_X1 c1061(
.A1(net1064),
.A2(net1056),
.ZN(net1099)
);

OAI22_X1 c1062(
.A1(net1055),
.A2(net1034),
.B1(net1083),
.B2(net1067),
.ZN(net1100)
);

OR2_X2 c1063(
.A1(net1048),
.A2(net973),
.ZN(net1101)
);

NOR2_X4 c1064(
.A1(net126),
.A2(net10704),
.ZN(net1102)
);

DFFS_X1 c1065(
.D(net96),
.SN(net1099),
.CK(clk),
.Q(net1104),
.QN(net1103)
);

NOR2_X2 c1066(
.A1(net1096),
.A2(net10691),
.ZN(net1105)
);

XOR2_X2 c1067(
.A(net1104),
.B(net1037),
.Z(net1106)
);

AND4_X2 c1068(
.A1(net1057),
.A2(net1028),
.A3(net1067),
.A4(net1095),
.ZN(net1107)
);

XNOR2_X1 c1069(
.A(net1096),
.B(net1107),
.ZN(net1108)
);

OR2_X4 c1070(
.A1(net1107),
.A2(net1097),
.ZN(net1109)
);

OAI221_X4 c1071(
.A(net1099),
.B1(net1083),
.B2(net965),
.C1(net1035),
.C2(net1107),
.ZN(net1110)
);

INV_X4 c1072(
.A(net10893),
.ZN(net1111)
);

SDFFS_X1 c1073(
.D(net1106),
.SE(net1110),
.SI(net1095),
.SN(net1107),
.CK(clk),
.Q(net1113),
.QN(net1112)
);

OR2_X1 c1074(
.A1(net138),
.A2(net1111),
.ZN(net1114)
);

XNOR2_X2 c1075(
.A(net1111),
.B(net1045),
.ZN(net1115)
);

AOI222_X1 c1076(
.A1(net1033),
.A2(net1103),
.B1(net1056),
.B2(net1100),
.C1(net1107),
.C2(net11500),
.ZN(net1116)
);

SDFFS_X2 c1077(
.D(net1093),
.SE(net1115),
.SI(net1086),
.SN(net11502),
.CK(clk),
.Q(net1118),
.QN(net1117)
);

AOI222_X4 c1078(
.A1(net984),
.A2(net1117),
.B1(net1107),
.B2(net1086),
.C1(net10704),
.C2(net11502),
.ZN(net1119)
);

INV_X1 c1079(
.A(net9814),
.ZN(net1120)
);

INV_X2 c1080(
.A(net9790),
.ZN(net1121)
);

INV_X8 c1081(
.A(net158),
.ZN(net1122)
);

INV_X16 c1082(
.A(net189),
.ZN(net1123)
);

INV_X32 c1083(
.A(net9790),
.ZN(net1124)
);

INV_X4 c1084(
.A(net1105),
.ZN(net1125)
);

AND2_X4 c1085(
.A1(in25),
.A2(net59),
.ZN(net1126)
);

INV_X1 c1086(
.A(net196),
.ZN(net1127)
);

INV_X2 c1087(
.A(net90),
.ZN(net1128)
);

AND2_X1 c1088(
.A1(net1096),
.A2(net1126),
.ZN(net1129)
);

INV_X8 c1089(
.A(net1047),
.ZN(net1130)
);

INV_X16 c1090(
.A(net1022),
.ZN(net1131)
);

INV_X32 c1091(
.A(net1084),
.ZN(net1132)
);

INV_X4 c1092(
.A(net181),
.ZN(net1133)
);

NOR3_X2 c1093(
.A1(net1133),
.A2(net987),
.A3(net1123),
.ZN(net1134)
);

INV_X1 c1094(
.A(net1066),
.ZN(net1135)
);

INV_X2 c1095(
.A(net9813),
.ZN(net1136)
);

INV_X8 c1096(
.A(net1042),
.ZN(net1137)
);

INV_X16 c1097(
.A(net962),
.ZN(net1138)
);

INV_X32 c1098(
.A(net226),
.ZN(net1139)
);

INV_X4 c1099(
.A(net1044),
.ZN(net1140)
);

INV_X1 c1100(
.A(net221),
.ZN(net1141)
);

INV_X2 c1101(
.A(net1124),
.ZN(net1142)
);

INV_X8 c1102(
.A(net1122),
.ZN(net1143)
);

INV_X16 c1103(
.A(net10300),
.ZN(net1144)
);

NAND2_X1 c1104(
.A1(net1127),
.A2(net11503),
.ZN(net1145)
);

INV_X32 c1105(
.A(net9845),
.ZN(net1146)
);

INV_X4 c1106(
.A(net10832),
.ZN(net1147)
);

INV_X1 c1107(
.A(net9951),
.ZN(net1148)
);

NAND2_X2 c1108(
.A1(net1136),
.A2(net1145),
.ZN(net1149)
);

INV_X2 c1109(
.A(net987),
.ZN(net1150)
);

DFFRS_X2 c1110(
.D(net232),
.RN(net202),
.SN(net944),
.CK(clk),
.Q(net1152),
.QN(net1151)
);

NAND2_X4 c1111(
.A1(net113),
.A2(net1066),
.ZN(net1153)
);

AND2_X2 c1112(
.A1(net1149),
.A2(net1137),
.ZN(net1154)
);

AND3_X4 c1113(
.A1(net1042),
.A2(net1145),
.A3(net11503),
.ZN(net1155)
);

INV_X8 c1114(
.A(net204),
.ZN(net1156)
);

XOR2_X1 c1115(
.A(net1126),
.B(net1148),
.Z(net1157)
);

INV_X16 c1116(
.A(net10827),
.ZN(net1158)
);

INV_X32 c1117(
.A(net167),
.ZN(net1159)
);

SDFF_X1 c1118(
.D(net1159),
.SE(net1154),
.SI(net1137),
.CK(clk),
.Q(net1161),
.QN(net1160)
);

NOR2_X1 c1119(
.A1(net1087),
.A2(net1137),
.ZN(net1162)
);

OR2_X2 c1120(
.A1(net162),
.A2(net1133),
.ZN(net1163)
);

NAND3_X2 c1121(
.A1(net109),
.A2(net1160),
.A3(net1100),
.ZN(net1164)
);

INV_X4 c1122(
.A(net167),
.ZN(net1165)
);

NOR2_X4 c1123(
.A1(net196),
.A2(net90),
.ZN(net1166)
);

DFFS_X2 c1124(
.D(net230),
.SN(net1162),
.CK(clk),
.Q(net1168),
.QN(net1167)
);

NOR2_X2 c1125(
.A1(net1122),
.A2(net1127),
.ZN(net1169)
);

INV_X1 c1126(
.A(net113),
.ZN(net1170)
);

XOR2_X2 c1127(
.A(net68),
.B(net1161),
.Z(net1171)
);

XNOR2_X1 c1128(
.A(net1156),
.B(net1164),
.ZN(net1172)
);

INV_X2 c1129(
.A(net1170),
.ZN(net1173)
);

OR3_X1 c1130(
.A1(net1092),
.A2(net1006),
.A3(net11503),
.ZN(net1174)
);

MUX2_X1 c1131(
.A(net1150),
.B(net1166),
.S(net1135),
.Z(net1175)
);

OR2_X4 c1132(
.A1(net195),
.A2(net221),
.ZN(net1176)
);

INV_X8 c1133(
.A(net11054),
.ZN(net1177)
);

OR2_X1 c1134(
.A1(net1147),
.A2(net229),
.ZN(net1178)
);

XNOR2_X2 c1135(
.A(net1178),
.B(net1166),
.ZN(net1179)
);

AND2_X4 c1136(
.A1(net202),
.A2(net1100),
.ZN(net1180)
);

INV_X16 c1137(
.A(net1143),
.ZN(net1181)
);

OAI21_X4 c1138(
.A(net1131),
.B1(net1181),
.B2(net87),
.ZN(net1182)
);

AND2_X1 c1139(
.A1(net59),
.A2(net1157),
.ZN(net1183)
);

NAND2_X1 c1140(
.A1(net1146),
.A2(net1176),
.ZN(net1184)
);

MUX2_X2 c1141(
.A(net1125),
.B(net1130),
.S(net1022),
.Z(net1185)
);

NAND2_X2 c1142(
.A1(net1123),
.A2(net1183),
.ZN(net1186)
);

NAND3_X4 c1143(
.A1(net1136),
.A2(net1176),
.A3(net109),
.ZN(net1187)
);

SDFF_X2 c1144(
.D(net1172),
.SE(net1181),
.SI(net1182),
.CK(clk),
.Q(net1189),
.QN(net1188)
);

OR3_X4 c1145(
.A1(net1187),
.A2(net1178),
.A3(net1186),
.ZN(net1190)
);

NAND2_X4 c1146(
.A1(net1183),
.A2(net1177),
.ZN(net1191)
);

INV_X32 c1147(
.A(net1173),
.ZN(net1192)
);

AND3_X2 c1148(
.A1(net183),
.A2(net1145),
.A3(net1182),
.ZN(net1193)
);

AND2_X2 c1149(
.A1(net1157),
.A2(net1144),
.ZN(net1194)
);

NOR3_X1 c1150(
.A1(net1192),
.A2(net226),
.A3(net1194),
.ZN(net1195)
);

OAI221_X2 c1151(
.A(net1174),
.B1(net1184),
.B2(net1182),
.C1(net954),
.C2(net1195),
.ZN(net1196)
);

OR3_X2 c1152(
.A1(net1182),
.A2(net1138),
.A3(net1167),
.ZN(net1197)
);

OAI21_X2 c1153(
.A(net1184),
.B1(net1195),
.B2(net1131),
.ZN(net1198)
);

OAI21_X1 c1154(
.A(net1168),
.B1(net1195),
.B2(net11129),
.ZN(net1199)
);

XOR2_X1 c1155(
.A(net197),
.B(net11129),
.Z(net1200)
);

NOR2_X1 c1156(
.A1(net1194),
.A2(net1193),
.ZN(net1201)
);

DFFR_X1 c1157(
.D(net1201),
.RN(net195),
.CK(clk),
.Q(net1203),
.QN(net1202)
);

DFFRS_X1 c1158(
.D(net1200),
.RN(net1195),
.SN(net1201),
.CK(clk),
.Q(net1205),
.QN(net1204)
);

AOI21_X2 c1159(
.A(net1148),
.B1(net1192),
.B2(net1125),
.ZN(net1206)
);

AOI21_X1 c1160(
.A(net1171),
.B1(net1197),
.B2(net1191),
.ZN(net1207)
);

OAI33_X1 c1161(
.A1(net949),
.A2(net1207),
.A3(net1195),
.B1(net1095),
.B2(net1066),
.B3(net10696),
.ZN(net1208)
);

INV_X4 c1162(
.A(net9869),
.ZN(net1209)
);

INV_X1 c1163(
.A(net266),
.ZN(net1210)
);

INV_X2 c1164(
.A(net254),
.ZN(net1211)
);

INV_X8 c1165(
.A(net1138),
.ZN(net1212)
);

INV_X16 c1166(
.A(net1006),
.ZN(net1213)
);

INV_X32 c1167(
.A(net11085),
.ZN(net1214)
);

INV_X4 c1168(
.A(net11085),
.ZN(net1215)
);

INV_X1 c1169(
.A(net1212),
.ZN(net1216)
);

INV_X2 c1170(
.A(net1216),
.ZN(net1217)
);

INV_X8 c1171(
.A(net11336),
.ZN(net1218)
);

INV_X16 c1172(
.A(net1197),
.ZN(net1219)
);

OR2_X2 c1173(
.A1(net214),
.A2(net1186),
.ZN(net1220)
);

INV_X32 c1174(
.A(net266),
.ZN(net1221)
);

INV_X4 c1175(
.A(net10111),
.ZN(net1222)
);

INV_X1 c1176(
.A(net1039),
.ZN(net1223)
);

INV_X2 c1177(
.A(net10370),
.ZN(net1224)
);

NOR2_X4 c1178(
.A1(net1100),
.A2(net1086),
.ZN(net1225)
);

NOR2_X2 c1179(
.A1(net1219),
.A2(net1195),
.ZN(net1226)
);

XOR2_X2 c1180(
.A(net1166),
.B(net241),
.Z(net1227)
);

XNOR2_X1 c1181(
.A(net1039),
.B(net1210),
.ZN(net1228)
);

INV_X8 c1182(
.A(net1152),
.ZN(net1229)
);

INV_X16 c1183(
.A(net10112),
.ZN(net1230)
);

INV_X32 c1184(
.A(net255),
.ZN(net1231)
);

INV_X4 c1185(
.A(net10534),
.ZN(net1232)
);

AOI21_X4 c1186(
.A(net1187),
.B1(net1154),
.B2(net1228),
.ZN(net1233)
);

INV_X1 c1187(
.A(net1129),
.ZN(net1234)
);

INV_X2 c1188(
.A(net1222),
.ZN(net1235)
);

OR2_X4 c1189(
.A1(net1153),
.A2(net1214),
.ZN(net1236)
);

AND3_X1 c1190(
.A1(net197),
.A2(net1068),
.A3(net1121),
.ZN(net1237)
);

OR2_X1 c1191(
.A1(net325),
.A2(net1213),
.ZN(net1238)
);

INV_X8 c1192(
.A(net1232),
.ZN(net1239)
);

INV_X16 c1193(
.A(net1232),
.ZN(net1240)
);

INV_X32 c1194(
.A(net1231),
.ZN(net1241)
);

XNOR2_X2 c1195(
.A(net1069),
.B(net57),
.ZN(net1242)
);

AND2_X4 c1196(
.A1(net1215),
.A2(net1224),
.ZN(net1243)
);

AND2_X1 c1197(
.A1(net1234),
.A2(net1243),
.ZN(net1244)
);

INV_X4 c1198(
.A(net1134),
.ZN(net1245)
);

INV_X1 c1199(
.A(net1133),
.ZN(net1246)
);

NAND2_X1 c1200(
.A1(net1209),
.A2(net11131),
.ZN(net1247)
);

NAND2_X2 c1201(
.A1(net1181),
.A2(net1243),
.ZN(net1248)
);

INV_X2 c1202(
.A(net1245),
.ZN(net1249)
);

DFFR_X2 c1203(
.D(net1154),
.RN(net315),
.CK(clk),
.Q(net1251),
.QN(net1250)
);

INV_X8 c1204(
.A(net9845),
.ZN(net1252)
);

INV_X16 c1205(
.A(net1251),
.ZN(net1253)
);

INV_X32 c1206(
.A(net1223),
.ZN(net1254)
);

NAND2_X4 c1207(
.A1(net944),
.A2(net1243),
.ZN(net1255)
);

NAND3_X1 c1208(
.A1(net1249),
.A2(net1228),
.A3(net1230),
.ZN(net1256)
);

NOR3_X4 c1209(
.A1(net241),
.A2(net1256),
.A3(net1210),
.ZN(net1257)
);

INV_X4 c1210(
.A(net1246),
.ZN(net1258)
);

AND2_X2 c1211(
.A1(net1242),
.A2(net1215),
.ZN(net1259)
);

INV_X1 c1212(
.A(net1235),
.ZN(net1260)
);

AND4_X1 c1213(
.A1(net1176),
.A2(net313),
.A3(net45),
.A4(net1086),
.ZN(net1261)
);

XOR2_X1 c1214(
.A(net1120),
.B(net1246),
.Z(net1262)
);

NOR2_X1 c1215(
.A1(net1248),
.A2(net1255),
.ZN(net1263)
);

INV_X2 c1216(
.A(net11157),
.ZN(net1264)
);

OR2_X2 c1217(
.A1(net1243),
.A2(net1258),
.ZN(net1265)
);

INV_X8 c1218(
.A(net1261),
.ZN(net1266)
);

NOR2_X4 c1219(
.A1(net1219),
.A2(net1248),
.ZN(net1267)
);

NOR2_X2 c1220(
.A1(net1237),
.A2(net1234),
.ZN(net1268)
);

XOR2_X2 c1221(
.A(net1258),
.B(net1243),
.Z(net1269)
);

INV_X16 c1222(
.A(net10120),
.ZN(net1270)
);

XNOR2_X1 c1223(
.A(net1231),
.B(net1255),
.ZN(net1271)
);

OR2_X4 c1224(
.A1(net1244),
.A2(net1245),
.ZN(net1272)
);

NOR3_X2 c1225(
.A1(net1139),
.A2(net312),
.A3(net1272),
.ZN(net1273)
);

AND3_X4 c1226(
.A1(net313),
.A2(net1265),
.A3(net1242),
.ZN(net1274)
);

OR2_X1 c1227(
.A1(net1211),
.A2(net1235),
.ZN(net1275)
);

XNOR2_X2 c1228(
.A(net1268),
.B(net1006),
.ZN(net1276)
);

AND2_X4 c1229(
.A1(net1274),
.A2(net10538),
.ZN(net1277)
);

AND2_X1 c1230(
.A1(net1273),
.A2(net1228),
.ZN(net1278)
);

NAND2_X1 c1231(
.A1(net17),
.A2(net1244),
.ZN(net1279)
);

NAND3_X2 c1232(
.A1(net1264),
.A2(net1277),
.A3(net1269),
.ZN(net1280)
);

NAND2_X2 c1233(
.A1(net253),
.A2(net1246),
.ZN(net1281)
);

OR3_X1 c1234(
.A1(net1276),
.A2(net1251),
.A3(net1224),
.ZN(net1282)
);

DFFRS_X2 c1235(
.D(net1256),
.RN(net1231),
.SN(net1219),
.CK(clk),
.Q(net1284),
.QN(net1283)
);

MUX2_X1 c1236(
.A(net1281),
.B(net1268),
.S(net1282),
.Z(net1285)
);

OAI21_X4 c1237(
.A(net1239),
.B1(net1137),
.B2(net11158),
.ZN(net1286)
);

MUX2_X2 c1238(
.A(net1265),
.B(net1259),
.S(net1232),
.Z(net1287)
);

AOI222_X2 c1239(
.A1(net1264),
.A2(net1100),
.B1(net1217),
.B2(net1247),
.C1(net258),
.C2(net11361),
.ZN(net1288)
);

AOI22_X4 c1240(
.A1(net1259),
.A2(net1268),
.B1(net1166),
.B2(net1212),
.ZN(net1289)
);

OAI22_X4 c1241(
.A1(net1287),
.A2(net1256),
.B1(net1282),
.B2(net1251),
.ZN(net1290)
);

OAI222_X1 c1242(
.A1(net303),
.A2(net1260),
.B1(net253),
.B2(net1250),
.C1(net1212),
.C2(net258),
.ZN(net1291)
);

NAND2_X4 c1243(
.A1(net1271),
.A2(net1289),
.ZN(net1292)
);

AND2_X2 c1244(
.A1(net1274),
.A2(net1281),
.ZN(net1293)
);

INV_X32 c1245(
.A(net11073),
.ZN(net1294)
);

INV_X4 c1246(
.A(net338),
.ZN(net1295)
);

INV_X1 c1247(
.A(net1179),
.ZN(net1296)
);

INV_X2 c1248(
.A(net10539),
.ZN(net1297)
);

XOR2_X1 c1249(
.A(net305),
.B(net1163),
.Z(net1298)
);

INV_X8 c1250(
.A(net1228),
.ZN(net1299)
);

INV_X16 c1251(
.A(net1121),
.ZN(net1300)
);

INV_X32 c1252(
.A(net11398),
.ZN(net1301)
);

NOR2_X1 c1253(
.A1(net1297),
.A2(net10833),
.ZN(net1302)
);

INV_X4 c1254(
.A(net9714),
.ZN(net1303)
);

INV_X1 c1255(
.A(net11073),
.ZN(net1304)
);

INV_X2 c1256(
.A(net1299),
.ZN(net1305)
);

OR2_X2 c1257(
.A1(net185),
.A2(net408),
.ZN(net1306)
);

INV_X8 c1258(
.A(net9714),
.ZN(net1307)
);

INV_X16 c1259(
.A(net1303),
.ZN(net1308)
);

INV_X32 c1260(
.A(net1258),
.ZN(net1309)
);

NOR2_X4 c1261(
.A1(net45),
.A2(net1277),
.ZN(net1310)
);

DFFS_X1 c1262(
.D(net403),
.SN(net1193),
.CK(clk),
.Q(net1312),
.QN(net1311)
);

NAND3_X4 c1263(
.A1(net1260),
.A2(net1217),
.A3(net10944),
.ZN(net1313)
);

INV_X4 c1264(
.A(net1137),
.ZN(net1314)
);

INV_X1 c1265(
.A(net323),
.ZN(net1315)
);

INV_X2 c1266(
.A(net1301),
.ZN(net1316)
);

INV_X8 c1267(
.A(net1138),
.ZN(net1317)
);

INV_X16 c1268(
.A(net1300),
.ZN(net1318)
);

AOI221_X4 c1269(
.A(net227),
.B1(net1317),
.B2(net1212),
.C1(net1086),
.C2(net1247),
.ZN(net1319)
);

INV_X32 c1270(
.A(net269),
.ZN(net1320)
);

INV_X4 c1271(
.A(net1260),
.ZN(net1321)
);

NOR2_X2 c1272(
.A1(net1209),
.A2(net1224),
.ZN(net1322)
);

INV_X1 c1273(
.A(net1158),
.ZN(net1323)
);

INV_X2 c1274(
.A(net1163),
.ZN(net1324)
);

INV_X8 c1275(
.A(net9902),
.ZN(net1325)
);

XOR2_X2 c1276(
.A(net1217),
.B(net11131),
.Z(net1326)
);

INV_X16 c1277(
.A(net389),
.ZN(net1327)
);

INV_X32 c1278(
.A(net1180),
.ZN(net1328)
);

INV_X4 c1279(
.A(net1308),
.ZN(net1329)
);

INV_X1 c1280(
.A(net1322),
.ZN(net1330)
);

SDFFR_X1 c1281(
.D(net1295),
.RN(net1286),
.SE(net1303),
.SI(net408),
.CK(clk),
.Q(net1332),
.QN(net1331)
);

INV_X2 c1282(
.A(net1323),
.ZN(net1333)
);

INV_X8 c1283(
.A(net1330),
.ZN(net1334)
);

XNOR2_X1 c1284(
.A(net1332),
.B(net290),
.ZN(net1335)
);

INV_X16 c1285(
.A(net1302),
.ZN(net1336)
);

OR3_X4 c1286(
.A1(net1328),
.A2(net1228),
.A3(net1317),
.ZN(net1337)
);

INV_X32 c1287(
.A(net1320),
.ZN(net1338)
);

INV_X4 c1288(
.A(net11039),
.ZN(net1339)
);

INV_X1 c1289(
.A(net9885),
.ZN(net1340)
);

INV_X2 c1290(
.A(net11158),
.ZN(net1341)
);

AOI22_X2 c1291(
.A1(net330),
.A2(net1317),
.B1(net1297),
.B2(net10833),
.ZN(net1342)
);

OR2_X4 c1292(
.A1(net1335),
.A2(net1341),
.ZN(net1343)
);

INV_X8 c1293(
.A(net11336),
.ZN(net1344)
);

INV_X16 c1294(
.A(net1321),
.ZN(net1345)
);

INV_X32 c1295(
.A(net1345),
.ZN(net1346)
);

OR2_X1 c1296(
.A1(net1305),
.A2(net1225),
.ZN(net1347)
);

INV_X4 c1297(
.A(net9902),
.ZN(net1348)
);

XNOR2_X2 c1298(
.A(net1329),
.B(net1330),
.ZN(net1349)
);

AND2_X4 c1299(
.A1(net1349),
.A2(net1323),
.ZN(net1350)
);

INV_X1 c1300(
.A(net10931),
.ZN(net1351)
);

AND2_X1 c1301(
.A1(net337),
.A2(net1343),
.ZN(net1352)
);

INV_X2 c1302(
.A(net393),
.ZN(net1353)
);

AND3_X2 c1303(
.A1(net377),
.A2(net1323),
.A3(net11039),
.ZN(net1354)
);

NAND2_X1 c1304(
.A1(net1168),
.A2(net1349),
.ZN(net1355)
);

NAND2_X2 c1305(
.A1(net1296),
.A2(net1351),
.ZN(net1356)
);

NAND2_X4 c1306(
.A1(net1352),
.A2(net1212),
.ZN(net1357)
);

AND2_X2 c1307(
.A1(net1315),
.A2(net1340),
.ZN(net1358)
);

INV_X8 c1308(
.A(net1356),
.ZN(net1359)
);

SDFFR_X2 c1309(
.D(net1313),
.RN(net409),
.SE(net415),
.SI(net1247),
.CK(clk),
.Q(net1361),
.QN(net1360)
);

INV_X16 c1310(
.A(net1342),
.ZN(net1362)
);

INV_X32 c1311(
.A(net11221),
.ZN(net1363)
);

XOR2_X1 c1312(
.A(net370),
.B(net1179),
.Z(net1364)
);

NOR2_X1 c1313(
.A1(net1218),
.A2(net1351),
.ZN(net1365)
);

NOR3_X1 c1314(
.A1(net1363),
.A2(net1358),
.A3(net999),
.ZN(net1366)
);

OR2_X2 c1315(
.A1(net1346),
.A2(net1311),
.ZN(net1367)
);

INV_X4 c1316(
.A(net11055),
.ZN(net1368)
);

NAND4_X4 c1317(
.A1(net1367),
.A2(net1323),
.A3(net1343),
.A4(net10839),
.ZN(net1369)
);

OR3_X2 c1318(
.A1(net1325),
.A2(net1308),
.A3(net1329),
.ZN(net1370)
);

OAI211_X2 c1319(
.A(net1266),
.B(net1212),
.C1(net350),
.C2(net1351),
.ZN(net1371)
);

NOR2_X4 c1320(
.A1(net1331),
.A2(net11245),
.ZN(net1372)
);

OAI21_X2 c1321(
.A(net1368),
.B1(net1369),
.B2(net11245),
.ZN(net1373)
);

NOR2_X2 c1322(
.A1(net1362),
.A2(net1373),
.ZN(net1374)
);

OAI21_X1 c1323(
.A(net1284),
.B1(net1329),
.B2(net10840),
.ZN(net1375)
);

AOI221_X2 c1324(
.A(net1357),
.B1(net1358),
.B2(net1351),
.C1(net1374),
.C2(net1353),
.ZN(net1376)
);

SDFF_X1 c1325(
.D(net1221),
.SE(net1266),
.SI(net1319),
.CK(clk),
.Q(net1378),
.QN(net1377)
);

XOR2_X2 c1326(
.A(net1370),
.B(net1354),
.Z(net1379)
);

AOI21_X2 c1327(
.A(net1376),
.B1(net1377),
.B2(net1379),
.ZN(net1380)
);

INV_X1 c1328(
.A(net9870),
.ZN(net1381)
);

INV_X2 c1329(
.A(net1372),
.ZN(net1382)
);

XNOR2_X1 c1330(
.A(net310),
.B(net423),
.ZN(net1383)
);

INV_X8 c1331(
.A(net11215),
.ZN(net1384)
);

OR2_X4 c1332(
.A1(net1284),
.A2(net1277),
.ZN(net1385)
);

INV_X16 c1333(
.A(net1149),
.ZN(net1386)
);

OR2_X1 c1334(
.A1(net168),
.A2(net1353),
.ZN(net1387)
);

SDFF_X2 c1335(
.D(net308),
.SE(net1225),
.SI(net1314),
.CK(clk),
.Q(net1389),
.QN(net1388)
);

XNOR2_X2 c1336(
.A(net156),
.B(net450),
.ZN(net1390)
);

INV_X32 c1337(
.A(net442),
.ZN(net1391)
);

AND2_X4 c1338(
.A1(net423),
.A2(net327),
.ZN(net1392)
);

AND2_X1 c1339(
.A1(net1390),
.A2(net1317),
.ZN(net1393)
);

INV_X4 c1340(
.A(net501),
.ZN(net1394)
);

NAND2_X1 c1341(
.A1(net1227),
.A2(net1378),
.ZN(net1395)
);

OR4_X2 c1342(
.A1(net431),
.A2(net1395),
.A3(net1336),
.A4(net1373),
.ZN(net1396)
);

INV_X1 c1343(
.A(net1277),
.ZN(net1397)
);

AOI21_X1 c1344(
.A(net1361),
.B1(net1294),
.B2(net449),
.ZN(net1398)
);

INV_X2 c1345(
.A(net439),
.ZN(net1399)
);

INV_X8 c1346(
.A(net456),
.ZN(net1400)
);

NAND2_X2 c1347(
.A1(net1237),
.A2(net1340),
.ZN(net1401)
);

NAND2_X4 c1348(
.A1(net1275),
.A2(net479),
.ZN(net1402)
);

INV_X16 c1349(
.A(net350),
.ZN(net1403)
);

DFFS_X2 c1350(
.D(net1314),
.SN(net483),
.CK(clk),
.Q(net1405),
.QN(net1404)
);

INV_X32 c1351(
.A(net10490),
.ZN(net1406)
);

INV_X4 c1352(
.A(net1304),
.ZN(net1407)
);

INV_X1 c1353(
.A(net11234),
.ZN(net1408)
);

INV_X2 c1354(
.A(net1395),
.ZN(net1409)
);

AND2_X2 c1355(
.A1(net1283),
.A2(net10960),
.ZN(net1410)
);

INV_X8 c1356(
.A(net1407),
.ZN(net1411)
);

INV_X16 c1357(
.A(net1344),
.ZN(net1412)
);

INV_X32 c1358(
.A(net414),
.ZN(net1413)
);

XOR2_X1 c1359(
.A(net430),
.B(net1402),
.Z(net1414)
);

INV_X4 c1360(
.A(net1392),
.ZN(net1415)
);

NOR2_X1 c1361(
.A1(net1312),
.A2(net1364),
.ZN(net1416)
);

OR2_X2 c1362(
.A1(net460),
.A2(net1412),
.ZN(net1417)
);

NOR2_X4 c1363(
.A1(net487),
.A2(net1414),
.ZN(net1418)
);

NOR2_X2 c1364(
.A1(net434),
.A2(net1360),
.ZN(net1419)
);

INV_X1 c1365(
.A(net11016),
.ZN(net1420)
);

INV_X2 c1366(
.A(net285),
.ZN(net1421)
);

INV_X8 c1367(
.A(net1420),
.ZN(net1422)
);

AOI211_X1 c1368(
.A(net1422),
.B(net1400),
.C1(net462),
.C2(net1086),
.ZN(net1423)
);

AOI21_X4 c1369(
.A(net1381),
.B1(net1394),
.B2(net1405),
.ZN(net1424)
);

INV_X16 c1370(
.A(net11286),
.ZN(net1425)
);

XOR2_X2 c1371(
.A(net479),
.B(net1408),
.Z(net1426)
);

XNOR2_X1 c1372(
.A(net1340),
.B(net442),
.ZN(net1427)
);

INV_X32 c1373(
.A(net1355),
.ZN(net1428)
);

INV_X4 c1374(
.A(net1424),
.ZN(net1429)
);

OR2_X4 c1375(
.A1(net1386),
.A2(net1360),
.ZN(net1430)
);

AND3_X1 c1376(
.A1(net1384),
.A2(net1301),
.A3(net1401),
.ZN(net1431)
);

OR2_X1 c1377(
.A1(net1416),
.A2(net434),
.ZN(net1432)
);

XNOR2_X2 c1378(
.A(net1429),
.B(net431),
.ZN(net1433)
);

INV_X1 c1379(
.A(net1301),
.ZN(net1434)
);

INV_X2 c1380(
.A(net11234),
.ZN(net1435)
);

INV_X8 c1381(
.A(net1396),
.ZN(net1436)
);

INV_X16 c1382(
.A(net1425),
.ZN(net1437)
);

SDFFRS_X2 c1383(
.D(net1397),
.RN(net1407),
.SE(net1420),
.SI(net1225),
.SN(net1412),
.CK(clk),
.Q(net1439),
.QN(net1438)
);

NAND3_X1 c1384(
.A1(net1378),
.A2(net1438),
.A3(net1409),
.ZN(net1440)
);

NAND4_X2 c1385(
.A1(net1440),
.A2(net1410),
.A3(net1428),
.A4(net1399),
.ZN(net1441)
);

DFFRS_X1 c1386(
.D(net1424),
.RN(net457),
.SN(net10840),
.CK(clk),
.Q(net1443),
.QN(net1442)
);

INV_X32 c1387(
.A(net10306),
.ZN(net1444)
);

AND2_X4 c1388(
.A1(net1408),
.A2(net1404),
.ZN(net1445)
);

INV_X4 c1389(
.A(net10016),
.ZN(net1446)
);

INV_X1 c1390(
.A(net10061),
.ZN(net1447)
);

AND2_X1 c1391(
.A1(net1447),
.A2(net1428),
.ZN(net1448)
);

NAND2_X1 c1392(
.A1(net1445),
.A2(net1353),
.ZN(net1449)
);

NOR3_X4 c1393(
.A1(net1417),
.A2(net1373),
.A3(net1442),
.ZN(net1450)
);

NAND2_X2 c1394(
.A1(net1444),
.A2(net11275),
.ZN(net1451)
);

NAND2_X4 c1395(
.A1(net1435),
.A2(net487),
.ZN(net1452)
);

AND2_X2 c1396(
.A1(net1450),
.A2(net1283),
.ZN(net1453)
);

XOR2_X1 c1397(
.A(net1452),
.B(net1374),
.Z(net1454)
);

NOR2_X1 c1398(
.A1(net1433),
.A2(net1408),
.ZN(net1455)
);

OR2_X2 c1399(
.A1(net1437),
.A2(net1431),
.ZN(net1456)
);

NOR3_X2 c1400(
.A1(net1439),
.A2(net1372),
.A3(net11275),
.ZN(net1457)
);

INV_X2 c1401(
.A(net11215),
.ZN(net1458)
);

AOI221_X1 c1402(
.A(net1457),
.B1(net1427),
.B2(net1411),
.C1(net350),
.C2(net1386),
.ZN(net1459)
);

OAI221_X1 c1403(
.A(net1449),
.B1(net1444),
.B2(net1365),
.C1(net1412),
.C2(net1428),
.ZN(net1460)
);

SDFFS_X1 c1404(
.D(net1336),
.SE(net1453),
.SI(net1440),
.SN(net1401),
.CK(clk),
.Q(net1462),
.QN(net1461)
);

OR4_X4 c1405(
.A1(net1419),
.A2(net1456),
.A3(net1461),
.A4(net1317),
.ZN(net1463)
);

INV_X8 c1406(
.A(net11367),
.ZN(net1464)
);

SDFFS_X2 c1407(
.D(net1456),
.SE(net1451),
.SI(net1418),
.SN(net11116),
.CK(clk),
.Q(net1466),
.QN(net1465)
);

AND3_X4 c1408(
.A1(net1365),
.A2(net1464),
.A3(net1445),
.ZN(net1467)
);

NAND3_X2 c1409(
.A1(net1467),
.A2(net283),
.A3(net1457),
.ZN(net1468)
);

OAI222_X4 c1410(
.A1(net1383),
.A2(net1467),
.B1(net1465),
.B2(net1212),
.C1(net1412),
.C2(net11116),
.ZN(net1469)
);

INV_X16 c1411(
.A(net9934),
.ZN(net1470)
);

INV_X32 c1412(
.A(net9733),
.ZN(net1471)
);

NOR2_X4 c1413(
.A1(net551),
.A2(net1399),
.ZN(net1472)
);

NOR2_X2 c1414(
.A1(net399),
.A2(net1403),
.ZN(net1473)
);

OR3_X1 c1415(
.A1(net579),
.A2(net562),
.A3(net1309),
.ZN(net1474)
);

INV_X4 c1416(
.A(net9941),
.ZN(net1475)
);

XOR2_X2 c1417(
.A(net1436),
.B(net10758),
.Z(net1476)
);

XNOR2_X1 c1418(
.A(net1405),
.B(net1364),
.ZN(net1477)
);

INV_X1 c1419(
.A(net11423),
.ZN(net1478)
);

INV_X2 c1420(
.A(net1413),
.ZN(net1479)
);

INV_X8 c1421(
.A(net1439),
.ZN(net1480)
);

OR2_X4 c1422(
.A1(net578),
.A2(net465),
.ZN(net1481)
);

INV_X16 c1423(
.A(net1406),
.ZN(net1482)
);

OAI22_X2 c1424(
.A1(net530),
.A2(net524),
.B1(net375),
.B2(net1412),
.ZN(net1483)
);

MUX2_X1 c1425(
.A(net526),
.B(net508),
.S(net1451),
.Z(net1484)
);

INV_X32 c1426(
.A(net11408),
.ZN(net1485)
);

INV_X4 c1427(
.A(net548),
.ZN(net1486)
);

INV_X1 c1428(
.A(net1409),
.ZN(net1487)
);

INV_X2 c1429(
.A(net11408),
.ZN(net1488)
);

INV_X8 c1430(
.A(net257),
.ZN(net1489)
);

INV_X16 c1431(
.A(net11477),
.ZN(net1490)
);

INV_X32 c1432(
.A(net9885),
.ZN(net1491)
);

OR2_X1 c1433(
.A1(net1488),
.A2(net466),
.ZN(net1492)
);

INV_X4 c1434(
.A(net9889),
.ZN(net1493)
);

XNOR2_X2 c1435(
.A(net1213),
.B(net1294),
.ZN(net1494)
);

INV_X1 c1436(
.A(net1493),
.ZN(net1495)
);

DFFRS_X2 c1437(
.D(net1477),
.RN(net1492),
.SN(net11347),
.CK(clk),
.Q(net1497),
.QN(net1496)
);

INV_X2 c1438(
.A(net541),
.ZN(net1498)
);

INV_X8 c1439(
.A(net1490),
.ZN(net1499)
);

INV_X16 c1440(
.A(net11424),
.ZN(net1500)
);

AND2_X4 c1441(
.A1(net1486),
.A2(net257),
.ZN(net1501)
);

INV_X32 c1442(
.A(net513),
.ZN(net1502)
);

INV_X4 c1443(
.A(net1448),
.ZN(net1503)
);

AND2_X1 c1444(
.A1(net1478),
.A2(net1488),
.ZN(net1504)
);

NAND2_X1 c1445(
.A1(net362),
.A2(net1496),
.ZN(net1505)
);

INV_X1 c1446(
.A(net11407),
.ZN(net1506)
);

OAI21_X4 c1447(
.A(net1502),
.B1(net1482),
.B2(net526),
.ZN(net1507)
);

INV_X2 c1448(
.A(net9933),
.ZN(net1508)
);

MUX2_X2 c1449(
.A(net1473),
.B(net1503),
.S(net538),
.Z(net1509)
);

INV_X8 c1450(
.A(net11307),
.ZN(net1510)
);

OAI211_X4 c1451(
.A(net1294),
.B(net1438),
.C1(net1436),
.C2(net11075),
.ZN(net1511)
);

NAND2_X2 c1452(
.A1(net1471),
.A2(net586),
.ZN(net1512)
);

NAND2_X4 c1453(
.A1(net1462),
.A2(net1489),
.ZN(net1513)
);

INV_X16 c1454(
.A(net1451),
.ZN(net1514)
);

DFFR_X1 c1455(
.D(net1503),
.RN(net525),
.CK(clk),
.Q(net1516),
.QN(net1515)
);

NAND3_X4 c1456(
.A1(net1505),
.A2(net1490),
.A3(net1479),
.ZN(net1517)
);

AND2_X2 c1457(
.A1(net1317),
.A2(net1515),
.ZN(net1518)
);

INV_X32 c1458(
.A(net1410),
.ZN(net1519)
);

XOR2_X1 c1459(
.A(net447),
.B(net1513),
.Z(net1520)
);

INV_X4 c1460(
.A(net11347),
.ZN(net1521)
);

INV_X1 c1461(
.A(net1485),
.ZN(net1522)
);

NOR2_X1 c1462(
.A1(net1494),
.A2(net522),
.ZN(net1523)
);

OR2_X2 c1463(
.A1(net1508),
.A2(net450),
.ZN(net1524)
);

INV_X2 c1464(
.A(net1364),
.ZN(net1525)
);

NOR2_X4 c1465(
.A1(net1519),
.A2(net586),
.ZN(net1526)
);

NOR2_X2 c1466(
.A1(net508),
.A2(net589),
.ZN(net1527)
);

INV_X8 c1467(
.A(net9732),
.ZN(net1528)
);

INV_X16 c1468(
.A(net450),
.ZN(net1529)
);

XOR2_X2 c1469(
.A(net1495),
.B(net1488),
.Z(net1530)
);

OAI222_X2 c1470(
.A1(net562),
.A2(net1502),
.B1(net1530),
.B2(net543),
.C1(net1517),
.C2(net559),
.ZN(net1531)
);

OR3_X4 c1471(
.A1(net1498),
.A2(net586),
.A3(net1388),
.ZN(net1532)
);

XNOR2_X1 c1472(
.A(net1516),
.B(net1454),
.ZN(net1533)
);

AND3_X2 c1473(
.A1(net1203),
.A2(net579),
.A3(net258),
.ZN(net1534)
);

NOR3_X1 c1474(
.A1(net1512),
.A2(net1462),
.A3(net562),
.ZN(net1535)
);

OR2_X4 c1475(
.A1(net1492),
.A2(net1517),
.ZN(net1536)
);

OR3_X2 c1476(
.A1(net525),
.A2(net1524),
.A3(net1528),
.ZN(net1537)
);

OR2_X1 c1477(
.A1(net1536),
.A2(net1517),
.ZN(net1538)
);

OAI21_X2 c1478(
.A(net1497),
.B1(net530),
.B2(net1528),
.ZN(net1539)
);

XNOR2_X2 c1479(
.A(net1510),
.B(net11308),
.ZN(net1540)
);

AND2_X4 c1480(
.A1(net1500),
.A2(net1506),
.ZN(net1541)
);

AND2_X1 c1481(
.A1(net1520),
.A2(net1526),
.ZN(net1542)
);

SDFF_X1 c1482(
.D(net1517),
.SE(net1410),
.SI(net1542),
.CK(clk),
.Q(net1544),
.QN(net1543)
);

OAI21_X1 c1483(
.A(net1516),
.B1(net1543),
.B2(net11397),
.ZN(net1545)
);

AOI222_X1 c1484(
.A1(net1480),
.A2(net1532),
.B1(net1519),
.B2(net1217),
.C1(net1513),
.C2(net586),
.ZN(net1546)
);

SDFF_X2 c1485(
.D(net1385),
.SE(net1497),
.SI(net1542),
.CK(clk),
.Q(net1548),
.QN(net1547)
);

DFFRS_X1 c1486(
.D(net1547),
.RN(net1542),
.SN(net11074),
.CK(clk),
.Q(net1550),
.QN(net1549)
);

DFFRS_X2 c1487(
.D(net1524),
.RN(net1490),
.SN(net1542),
.CK(clk),
.Q(net1552),
.QN(net1551)
);

OAI211_X1 c1488(
.A(net1528),
.B(net1512),
.C1(net1534),
.C2(net1517),
.ZN(net1553)
);

AOI222_X4 c1489(
.A1(net1389),
.A2(net1506),
.B1(net1522),
.B2(net1542),
.C1(net586),
.C2(net559),
.ZN(net1554)
);

AOI21_X2 c1490(
.A(net1534),
.B1(net1551),
.B2(net11059),
.ZN(net1555)
);

SDFF_X1 c1491(
.D(net1521),
.SE(net1542),
.SI(net1555),
.CK(clk),
.Q(net1557),
.QN(net1556)
);

AOI21_X1 c1492(
.A(net1556),
.B1(net1541),
.B2(net11059),
.ZN(net1558)
);

AOI21_X4 c1493(
.A(net1546),
.B1(net1553),
.B2(net11307),
.ZN(net1559)
);

NAND2_X1 c1494(
.A1(net1055),
.A2(net642),
.ZN(net1560)
);

INV_X32 c1495(
.A(net11450),
.ZN(net1561)
);

INV_X4 c1496(
.A(net9906),
.ZN(net1562)
);

NOR4_X4 c1497(
.A1(net581),
.A2(net656),
.A3(net507),
.A4(net659),
.ZN(net1563)
);

INV_X1 c1498(
.A(net1558),
.ZN(net1564)
);

INV_X2 c1499(
.A(net614),
.ZN(net1565)
);

INV_X8 c1500(
.A(net665),
.ZN(net1566)
);

INV_X16 c1501(
.A(net672),
.ZN(net1567)
);

INV_X32 c1502(
.A(net681),
.ZN(net1568)
);

INV_X4 c1503(
.A(net586),
.ZN(net1569)
);

NAND2_X2 c1504(
.A1(net328),
.A2(net626),
.ZN(net1570)
);

INV_X1 c1505(
.A(net1565),
.ZN(net1571)
);

INV_X2 c1506(
.A(net568),
.ZN(net1572)
);

INV_X8 c1507(
.A(net1567),
.ZN(net1573)
);

AND3_X1 c1508(
.A1(net1565),
.A2(net642),
.A3(net1569),
.ZN(net1574)
);

NAND2_X4 c1509(
.A1(net655),
.A2(net346),
.ZN(net1575)
);

AND2_X2 c1510(
.A1(net606),
.A2(net1549),
.ZN(net1576)
);

INV_X16 c1511(
.A(net11450),
.ZN(net1577)
);

INV_X32 c1512(
.A(net1555),
.ZN(net1578)
);

INV_X4 c1513(
.A(net11057),
.ZN(net1579)
);

INV_X1 c1514(
.A(net11057),
.ZN(net1580)
);

INV_X2 c1515(
.A(net11360),
.ZN(net1581)
);

DFFR_X2 c1516(
.D(net1563),
.RN(net462),
.CK(clk),
.Q(net1583),
.QN(net1582)
);

INV_X8 c1517(
.A(net1567),
.ZN(net1584)
);

NAND3_X1 c1518(
.A1(net1574),
.A2(net1582),
.A3(net1560),
.ZN(net1585)
);

XOR2_X1 c1519(
.A(net1326),
.B(net1565),
.Z(net1586)
);

INV_X16 c1520(
.A(net11397),
.ZN(net1587)
);

NOR2_X1 c1521(
.A1(net643),
.A2(net462),
.ZN(net1588)
);

INV_X32 c1522(
.A(net1540),
.ZN(net1589)
);

INV_X4 c1523(
.A(net1550),
.ZN(net1590)
);

DFFS_X1 c1524(
.D(net1576),
.SN(net1583),
.CK(clk),
.Q(net1592),
.QN(net1591)
);

INV_X1 c1525(
.A(net642),
.ZN(net1593)
);

INV_X2 c1526(
.A(net1544),
.ZN(net1594)
);

INV_X8 c1527(
.A(net9906),
.ZN(net1595)
);

OR2_X2 c1528(
.A1(net1570),
.A2(net1447),
.ZN(net1596)
);

NOR2_X4 c1529(
.A1(net1560),
.A2(net613),
.ZN(net1597)
);

NOR2_X2 c1530(
.A1(net674),
.A2(net1373),
.ZN(net1598)
);

XOR2_X2 c1531(
.A(net1561),
.B(net1595),
.Z(net1599)
);

INV_X16 c1532(
.A(net1588),
.ZN(net1600)
);

INV_X32 c1533(
.A(net1585),
.ZN(net1601)
);

INV_X4 c1534(
.A(net633),
.ZN(net1602)
);

INV_X1 c1535(
.A(net375),
.ZN(net1603)
);

XNOR2_X1 c1536(
.A(net1600),
.B(net1529),
.ZN(net1604)
);

OR2_X4 c1537(
.A1(net645),
.A2(net1326),
.ZN(net1605)
);

OR2_X1 c1538(
.A1(net1578),
.A2(net1522),
.ZN(net1606)
);

INV_X2 c1539(
.A(net10212),
.ZN(net1607)
);

XNOR2_X2 c1540(
.A(net1577),
.B(net1604),
.ZN(net1608)
);

AND2_X4 c1541(
.A1(net1529),
.A2(net1578),
.ZN(net1609)
);

AND2_X1 c1542(
.A1(net1598),
.A2(net1601),
.ZN(net1610)
);

NAND2_X1 c1543(
.A1(net1569),
.A2(net1603),
.ZN(net1611)
);

INV_X8 c1544(
.A(net10282),
.ZN(net1612)
);

NOR4_X2 c1545(
.A1(net1593),
.A2(net1603),
.A3(net674),
.A4(net1599),
.ZN(net1613)
);

NAND2_X2 c1546(
.A1(net1579),
.A2(net1605),
.ZN(net1614)
);

OAI221_X4 c1547(
.A(net1426),
.B1(net1609),
.B2(net1590),
.C1(net466),
.C2(net634),
.ZN(net1615)
);

INV_X16 c1548(
.A(net1602),
.ZN(net1616)
);

NAND2_X4 c1549(
.A1(net1482),
.A2(net1550),
.ZN(net1617)
);

AND2_X2 c1550(
.A1(net1597),
.A2(net1565),
.ZN(net1618)
);

INV_X32 c1551(
.A(net1606),
.ZN(net1619)
);

XOR2_X1 c1552(
.A(net1596),
.B(net1426),
.Z(net1620)
);

NOR2_X1 c1553(
.A1(net462),
.A2(net1594),
.ZN(net1621)
);

INV_X4 c1554(
.A(net1575),
.ZN(net1622)
);

OR2_X2 c1555(
.A1(net1566),
.A2(net11004),
.ZN(net1623)
);

NOR2_X4 c1556(
.A1(net613),
.A2(net1590),
.ZN(net1624)
);

NOR2_X2 c1557(
.A1(net1590),
.A2(net1611),
.ZN(net1625)
);

NOR3_X4 c1558(
.A1(net1592),
.A2(net1623),
.A3(net483),
.ZN(net1626)
);

XOR2_X2 c1559(
.A(net1611),
.B(net1597),
.Z(net1627)
);

SDFFR_X1 c1560(
.D(net1617),
.RN(net1546),
.SE(net634),
.SI(net1599),
.CK(clk),
.Q(net1629),
.QN(net1628)
);

NOR3_X2 c1561(
.A1(net1622),
.A2(net1596),
.A3(net1600),
.ZN(net1630)
);

INV_X1 c1562(
.A(net9989),
.ZN(net1631)
);

AND3_X4 c1563(
.A1(net1620),
.A2(net1624),
.A3(net1591),
.ZN(net1632)
);

XNOR2_X1 c1564(
.A(net1612),
.B(net1426),
.ZN(net1633)
);

OR2_X4 c1565(
.A1(net1623),
.A2(net1630),
.ZN(net1634)
);

INV_X2 c1566(
.A(net1625),
.ZN(net1635)
);

SDFFR_X2 c1567(
.D(net1601),
.RN(net1627),
.SE(net1630),
.SI(net1635),
.CK(clk),
.Q(net1637),
.QN(net1636)
);

SDFFRS_X1 c1568(
.D(net1566),
.RN(net1574),
.SE(net1054),
.SI(net1586),
.SN(net1604),
.CK(clk),
.Q(net1639),
.QN(net1638)
);

OR2_X1 c1569(
.A1(net1631),
.A2(net10697),
.ZN(net1640)
);

AOI211_X4 c1570(
.A(net1630),
.B(net1639),
.C1(net1589),
.C2(net1635),
.ZN(net1641)
);

XNOR2_X2 c1571(
.A(net1620),
.B(net10698),
.ZN(net1642)
);

NAND3_X2 c1572(
.A1(net584),
.A2(net1640),
.A3(net11004),
.ZN(net1643)
);

OR3_X1 c1573(
.A1(net1572),
.A2(net1643),
.A3(net1599),
.ZN(net1644)
);

NOR4_X1 c1574(
.A1(net1616),
.A2(net1640),
.A3(net1584),
.A4(net1599),
.ZN(net1645)
);

AND2_X4 c1575(
.A1(net1627),
.A2(net1638),
.ZN(net1646)
);

MUX2_X1 c1576(
.A(net1589),
.B(net1499),
.S(net1644),
.Z(net1647)
);

INV_X8 c1577(
.A(net585),
.ZN(net1648)
);

INV_X16 c1578(
.A(net666),
.ZN(net1649)
);

OAI21_X4 c1579(
.A(net346),
.B1(net1373),
.B2(net1577),
.ZN(net1650)
);

INV_X32 c1580(
.A(net696),
.ZN(net1651)
);

INV_X4 c1581(
.A(net710),
.ZN(net1652)
);

INV_X1 c1582(
.A(net662),
.ZN(net1653)
);

INV_X2 c1583(
.A(net1217),
.ZN(net1654)
);

INV_X8 c1584(
.A(net1654),
.ZN(net1655)
);

AND2_X1 c1585(
.A1(net689),
.A2(net711),
.ZN(net1656)
);

AOI211_X2 c1586(
.A(net357),
.B(net1654),
.C1(net727),
.C2(net1599),
.ZN(net1657)
);

INV_X16 c1587(
.A(net1656),
.ZN(net1658)
);

INV_X32 c1588(
.A(net1639),
.ZN(net1659)
);

INV_X4 c1589(
.A(net739),
.ZN(net1660)
);

INV_X1 c1590(
.A(net600),
.ZN(net1661)
);

INV_X2 c1591(
.A(net1506),
.ZN(net1662)
);

NAND2_X1 c1592(
.A1(net1648),
.A2(net1645),
.ZN(net1663)
);

INV_X8 c1593(
.A(net673),
.ZN(net1664)
);

INV_X16 c1594(
.A(net1577),
.ZN(net1665)
);

NAND2_X2 c1595(
.A1(net1665),
.A2(net1643),
.ZN(net1666)
);

INV_X32 c1596(
.A(net1573),
.ZN(net1667)
);

INV_X4 c1597(
.A(net11256),
.ZN(net1668)
);

INV_X1 c1598(
.A(net1586),
.ZN(net1669)
);

INV_X2 c1599(
.A(net535),
.ZN(net1670)
);

INV_X8 c1600(
.A(net1649),
.ZN(net1671)
);

INV_X16 c1601(
.A(net734),
.ZN(net1672)
);

INV_X32 c1602(
.A(net11256),
.ZN(net1673)
);

INV_X4 c1603(
.A(net1568),
.ZN(net1674)
);

INV_X1 c1604(
.A(net716),
.ZN(net1675)
);

NAND2_X4 c1605(
.A1(net602),
.A2(net734),
.ZN(net1676)
);

MUX2_X2 c1606(
.A(net739),
.B(net698),
.S(net11005),
.Z(net1677)
);

INV_X2 c1607(
.A(net1676),
.ZN(net1678)
);

AND2_X2 c1608(
.A1(net1650),
.A2(net1675),
.ZN(net1679)
);

INV_X8 c1609(
.A(net1648),
.ZN(net1680)
);

INV_X16 c1610(
.A(net1672),
.ZN(net1681)
);

XOR2_X1 c1611(
.A(net1624),
.B(net1651),
.Z(net1682)
);

NOR2_X1 c1612(
.A1(net1612),
.A2(net1655),
.ZN(net1683)
);

OR2_X2 c1613(
.A1(net1564),
.A2(net760),
.ZN(net1684)
);

INV_X32 c1614(
.A(net1654),
.ZN(net1685)
);

INV_X4 c1615(
.A(net543),
.ZN(net1686)
);

NOR2_X4 c1616(
.A1(net1603),
.A2(net1640),
.ZN(net1687)
);

INV_X1 c1617(
.A(net9958),
.ZN(net1688)
);

NOR2_X2 c1618(
.A1(net1659),
.A2(net522),
.ZN(net1689)
);

XOR2_X2 c1619(
.A(net1671),
.B(net1672),
.Z(net1690)
);

INV_X2 c1620(
.A(net11393),
.ZN(net1691)
);

INV_X8 c1621(
.A(net11346),
.ZN(net1692)
);

INV_X16 c1622(
.A(net742),
.ZN(net1693)
);

INV_X32 c1623(
.A(net1664),
.ZN(net1694)
);

INV_X4 c1624(
.A(net9967),
.ZN(net1695)
);

DFFS_X2 c1625(
.D(net1678),
.SN(net1681),
.CK(clk),
.Q(net1697),
.QN(net1696)
);

INV_X1 c1626(
.A(net1652),
.ZN(net1698)
);

XNOR2_X1 c1627(
.A(net1682),
.B(net1683),
.ZN(net1699)
);

NAND3_X4 c1628(
.A1(net1661),
.A2(net1681),
.A3(net763),
.ZN(net1700)
);

OR3_X4 c1629(
.A1(net1669),
.A2(net1686),
.A3(net1698),
.ZN(net1701)
);

OR2_X4 c1630(
.A1(net737),
.A2(net1686),
.ZN(net1702)
);

OR2_X1 c1631(
.A1(net757),
.A2(net1701),
.ZN(net1703)
);

DFFR_X1 c1632(
.D(net1694),
.RN(net1681),
.CK(clk),
.Q(net1705),
.QN(net1704)
);

XNOR2_X2 c1633(
.A(net1665),
.B(net1651),
.ZN(net1706)
);

INV_X2 c1634(
.A(net10377),
.ZN(net1707)
);

AND2_X4 c1635(
.A1(net1587),
.A2(net1650),
.ZN(net1708)
);

AOI22_X1 c1636(
.A1(net1688),
.A2(net1254),
.B1(net705),
.B2(net666),
.ZN(net1709)
);

AND2_X1 c1637(
.A1(net660),
.A2(net1603),
.ZN(net1710)
);

DFFR_X2 c1638(
.D(net1709),
.RN(net1669),
.CK(clk),
.Q(net1712),
.QN(net1711)
);

NAND2_X1 c1639(
.A1(net1684),
.A2(net747),
.ZN(net1713)
);

AND3_X2 c1640(
.A1(net1674),
.A2(net1418),
.A3(net758),
.ZN(net1714)
);

INV_X8 c1641(
.A(net10495),
.ZN(net1715)
);

NAND2_X2 c1642(
.A1(net1655),
.A2(net1712),
.ZN(net1716)
);

INV_X16 c1643(
.A(net9970),
.ZN(net1717)
);

AND4_X4 c1644(
.A1(net1653),
.A2(net1715),
.A3(net1698),
.A4(net701),
.ZN(net1718)
);

NAND2_X4 c1645(
.A1(net1683),
.A2(net1582),
.ZN(net1719)
);

AND2_X2 c1646(
.A1(net1715),
.A2(net11299),
.ZN(net1720)
);

INV_X32 c1647(
.A(net1668),
.ZN(net1721)
);

XOR2_X1 c1648(
.A(net1676),
.B(net1701),
.Z(net1722)
);

NOR3_X1 c1649(
.A1(net1719),
.A2(net1707),
.A3(net1721),
.ZN(net1723)
);

NOR2_X1 c1650(
.A1(net1720),
.A2(net1693),
.ZN(net1724)
);

OR3_X2 c1651(
.A1(net1710),
.A2(net1716),
.A3(net659),
.ZN(net1725)
);

OAI21_X2 c1652(
.A(net1657),
.B1(net543),
.B2(net1719),
.ZN(net1726)
);

OAI21_X1 c1653(
.A(net695),
.B1(net1720),
.B2(net1581),
.ZN(net1727)
);

OR2_X2 c1654(
.A1(net1717),
.A2(net1650),
.ZN(net1728)
);

NOR2_X4 c1655(
.A1(net1727),
.A2(net1612),
.ZN(net1729)
);

NOR2_X2 c1656(
.A1(net1721),
.A2(net686),
.ZN(net1730)
);

DFFS_X1 c1657(
.D(net1726),
.SN(net1707),
.CK(clk),
.Q(net1732),
.QN(net1731)
);

OAI33_X1 c1658(
.A1(net1725),
.A2(net1676),
.A3(net1731),
.B1(net1414),
.B2(net720),
.B3(net1635),
.ZN(net1733)
);

NAND4_X1 c1659(
.A1(net584),
.A2(net1729),
.A3(net1672),
.A4(net1701),
.ZN(net1734)
);

AOI21_X2 c1660(
.A(net806),
.B1(net834),
.B2(net1686),
.ZN(net1735)
);

INV_X4 c1661(
.A(net1516),
.ZN(net1736)
);

XOR2_X2 c1662(
.A(net816),
.B(net11423),
.Z(net1737)
);

XNOR2_X1 c1663(
.A(net1621),
.B(net846),
.ZN(net1738)
);

AOI21_X1 c1664(
.A(net1718),
.B1(net774),
.B2(net11499),
.ZN(net1739)
);

INV_X1 c1665(
.A(net1670),
.ZN(net1740)
);

OR2_X4 c1666(
.A1(net1518),
.A2(net1414),
.ZN(net1741)
);

OR2_X1 c1667(
.A1(net684),
.A2(net779),
.ZN(net1742)
);

INV_X2 c1668(
.A(net11031),
.ZN(net1743)
);

INV_X8 c1669(
.A(net1640),
.ZN(net1744)
);

INV_X16 c1670(
.A(net1583),
.ZN(net1745)
);

INV_X32 c1671(
.A(net1744),
.ZN(net1746)
);

INV_X4 c1672(
.A(net9674),
.ZN(net1747)
);

XNOR2_X2 c1673(
.A(net845),
.B(net1595),
.ZN(net1748)
);

OAI221_X2 c1674(
.A(net750),
.B1(net626),
.B2(net1515),
.C1(net1599),
.C2(net1743),
.ZN(net1749)
);

INV_X1 c1675(
.A(net1581),
.ZN(net1750)
);

SDFF_X2 c1676(
.D(net851),
.SE(net1704),
.SI(net813),
.CK(clk),
.Q(net1752),
.QN(net1751)
);

AND2_X4 c1677(
.A1(net1747),
.A2(net1647),
.ZN(net1753)
);

INV_X2 c1678(
.A(net1694),
.ZN(net1754)
);

INV_X8 c1679(
.A(net1754),
.ZN(net1755)
);

INV_X16 c1680(
.A(net11340),
.ZN(net1756)
);

INV_X32 c1681(
.A(net9882),
.ZN(net1757)
);

INV_X4 c1682(
.A(net795),
.ZN(net1758)
);

SDFFS_X1 c1683(
.D(net1756),
.SE(net1757),
.SI(net771),
.SN(net834),
.CK(clk),
.Q(net1760),
.QN(net1759)
);

DFFRS_X1 c1684(
.D(net771),
.RN(net1757),
.SN(net745),
.CK(clk),
.Q(net1762),
.QN(net1761)
);

AND2_X1 c1685(
.A1(net1745),
.A2(net1716),
.ZN(net1763)
);

INV_X1 c1686(
.A(net770),
.ZN(net1764)
);

INV_X2 c1687(
.A(net808),
.ZN(net1765)
);

AOI21_X4 c1688(
.A(net847),
.B1(net1628),
.B2(net1751),
.ZN(net1766)
);

NAND2_X1 c1689(
.A1(net1765),
.A2(net1730),
.ZN(net1767)
);

NAND2_X2 c1690(
.A1(net1724),
.A2(net826),
.ZN(net1768)
);

NAND2_X4 c1691(
.A1(net1740),
.A2(net834),
.ZN(net1769)
);

INV_X8 c1692(
.A(net1739),
.ZN(net1770)
);

AND2_X2 c1693(
.A1(net1698),
.A2(net1755),
.ZN(net1771)
);

INV_X16 c1694(
.A(net813),
.ZN(net1772)
);

INV_X32 c1695(
.A(net9882),
.ZN(net1773)
);

INV_X4 c1696(
.A(net1746),
.ZN(net1774)
);

XOR2_X1 c1697(
.A(net1770),
.B(net1767),
.Z(net1775)
);

INV_X1 c1698(
.A(net799),
.ZN(net1776)
);

INV_X2 c1699(
.A(net1748),
.ZN(net1777)
);

INV_X8 c1700(
.A(net1757),
.ZN(net1778)
);

INV_X16 c1701(
.A(net1773),
.ZN(net1779)
);

INV_X32 c1702(
.A(net9913),
.ZN(net1780)
);

AOI222_X2 c1703(
.A1(net1699),
.A2(net795),
.B1(net1757),
.B2(net1750),
.C1(net1715),
.C2(net1743),
.ZN(net1781)
);

INV_X4 c1704(
.A(net9913),
.ZN(net1782)
);

INV_X1 c1705(
.A(net9888),
.ZN(net1783)
);

NOR2_X1 c1706(
.A1(net1705),
.A2(net1670),
.ZN(net1784)
);

AOI221_X4 c1707(
.A(net1780),
.B1(net1784),
.B2(net1217),
.C1(net1743),
.C2(net10591),
.ZN(net1785)
);

INV_X2 c1708(
.A(net11062),
.ZN(net1786)
);

INV_X8 c1709(
.A(net1778),
.ZN(net1787)
);

INV_X16 c1710(
.A(net1772),
.ZN(net1788)
);

OR2_X2 c1711(
.A1(net1786),
.A2(net694),
.ZN(net1789)
);

NOR2_X4 c1712(
.A1(net1763),
.A2(net1761),
.ZN(net1790)
);

INV_X32 c1713(
.A(net1749),
.ZN(net1791)
);

INV_X4 c1714(
.A(net822),
.ZN(net1792)
);

NOR2_X2 c1715(
.A1(net1649),
.A2(net1789),
.ZN(net1793)
);

AND3_X1 c1716(
.A1(net748),
.A2(net1780),
.A3(net662),
.ZN(net1794)
);

OR4_X1 c1717(
.A1(net1766),
.A2(net1749),
.A3(net1687),
.A4(net1743),
.ZN(net1795)
);

INV_X1 c1718(
.A(net1787),
.ZN(net1796)
);

NAND3_X1 c1719(
.A1(net1768),
.A2(net1499),
.A3(net10592),
.ZN(net1797)
);

INV_X2 c1720(
.A(net1707),
.ZN(net1798)
);

XOR2_X2 c1721(
.A(net1798),
.B(net1789),
.Z(net1799)
);

INV_X8 c1722(
.A(net1783),
.ZN(net1800)
);

XNOR2_X1 c1723(
.A(net1629),
.B(net1768),
.ZN(net1801)
);

OR2_X4 c1724(
.A1(net1789),
.A2(net1786),
.ZN(net1802)
);

INV_X16 c1725(
.A(net1735),
.ZN(net1803)
);

NOR3_X4 c1726(
.A1(net1736),
.A2(net1786),
.A3(net495),
.ZN(net1804)
);

NOR3_X2 c1727(
.A1(net1774),
.A2(net1803),
.A3(net783),
.ZN(net1805)
);

OR2_X1 c1728(
.A1(net1797),
.A2(net1764),
.ZN(net1806)
);

INV_X32 c1729(
.A(net9888),
.ZN(net1807)
);

XNOR2_X2 c1730(
.A(net1784),
.B(net1804),
.ZN(net1808)
);

AND2_X4 c1731(
.A1(net1795),
.A2(net1792),
.ZN(net1809)
);

AND2_X1 c1732(
.A1(net1793),
.A2(net1621),
.ZN(net1810)
);

INV_X4 c1733(
.A(net9674),
.ZN(net1811)
);

AND3_X4 c1734(
.A1(net1808),
.A2(net1699),
.A3(net1791),
.ZN(net1812)
);

NAND2_X1 c1735(
.A1(net1796),
.A2(net1779),
.ZN(net1813)
);

NAND3_X2 c1736(
.A1(net1769),
.A2(net1813),
.A3(net1788),
.ZN(net1814)
);

NAND2_X2 c1737(
.A1(net1813),
.A2(net1786),
.ZN(net1815)
);

OR3_X1 c1738(
.A1(net1595),
.A2(net1737),
.A3(net661),
.ZN(net1816)
);

NAND2_X4 c1739(
.A1(net798),
.A2(net1805),
.ZN(net1817)
);

MUX2_X1 c1740(
.A(net1804),
.B(net1817),
.S(net1789),
.Z(net1818)
);

OAI21_X4 c1741(
.A(net1811),
.B1(net1812),
.B2(net1817),
.ZN(net1819)
);

INV_X1 c1742(
.A(net11188),
.ZN(net1820)
);

INV_X2 c1743(
.A(net1799),
.ZN(net1821)
);

INV_X8 c1744(
.A(net1785),
.ZN(net1822)
);

AND2_X2 c1745(
.A1(net1788),
.A2(net1635),
.ZN(net1823)
);

INV_X16 c1746(
.A(net1814),
.ZN(net1824)
);

INV_X32 c1747(
.A(net1414),
.ZN(net1825)
);

XOR2_X1 c1748(
.A(net1755),
.B(net940),
.Z(net1826)
);

INV_X4 c1749(
.A(net10385),
.ZN(net1827)
);

INV_X1 c1750(
.A(net1804),
.ZN(net1828)
);

DFFS_X2 c1751(
.D(net941),
.SN(net901),
.CK(clk),
.Q(net1830),
.QN(net1829)
);

NOR2_X1 c1752(
.A1(net1830),
.A2(net1764),
.ZN(net1831)
);

OR2_X2 c1753(
.A1(net1825),
.A2(net1788),
.ZN(net1832)
);

NOR2_X4 c1754(
.A1(net816),
.A2(net887),
.ZN(net1833)
);

NOR2_X2 c1755(
.A1(net1833),
.A2(net905),
.ZN(net1834)
);

INV_X2 c1756(
.A(net9651),
.ZN(net1835)
);

INV_X8 c1757(
.A(net892),
.ZN(net1836)
);

XOR2_X2 c1758(
.A(net1827),
.B(net819),
.Z(net1837)
);

INV_X16 c1759(
.A(net848),
.ZN(net1838)
);

XNOR2_X1 c1760(
.A(net891),
.B(net1835),
.ZN(net1839)
);

OR2_X4 c1761(
.A1(net821),
.A2(net906),
.ZN(net1840)
);

INV_X32 c1762(
.A(net861),
.ZN(net1841)
);

OR2_X1 c1763(
.A1(net1835),
.A2(net1594),
.ZN(net1842)
);

SDFFS_X2 c1764(
.D(net1822),
.SE(net941),
.SI(net863),
.SN(net889),
.CK(clk),
.Q(net1844),
.QN(net1843)
);

XNOR2_X2 c1765(
.A(net905),
.B(net1715),
.ZN(net1845)
);

INV_X4 c1766(
.A(net1842),
.ZN(net1846)
);

AND2_X4 c1767(
.A1(net885),
.A2(net1824),
.ZN(net1847)
);

AND2_X1 c1768(
.A1(net915),
.A2(net1823),
.ZN(net1848)
);

INV_X1 c1769(
.A(net10930),
.ZN(net1849)
);

NAND2_X1 c1770(
.A1(net1764),
.A2(net1843),
.ZN(net1850)
);

MUX2_X2 c1771(
.A(net706),
.B(net899),
.S(net1824),
.Z(net1851)
);

SDFFR_X1 c1772(
.D(net927),
.RN(net1834),
.SE(net905),
.SI(net1824),
.CK(clk),
.Q(net1853),
.QN(net1852)
);

NAND2_X2 c1773(
.A1(net1738),
.A2(net1840),
.ZN(net1854)
);

NAND2_X4 c1774(
.A1(net886),
.A2(net1830),
.ZN(net1855)
);

AND2_X2 c1775(
.A1(net935),
.A2(net1838),
.ZN(net1856)
);

INV_X2 c1776(
.A(net887),
.ZN(net1857)
);

INV_X8 c1777(
.A(net1716),
.ZN(net1858)
);

XOR2_X1 c1778(
.A(net1839),
.B(net1843),
.Z(net1859)
);

NOR2_X1 c1779(
.A1(net1853),
.A2(net915),
.ZN(net1860)
);

NAND3_X4 c1780(
.A1(net1309),
.A2(net1799),
.A3(net784),
.ZN(net1861)
);

INV_X16 c1781(
.A(net1850),
.ZN(net1862)
);

OR2_X2 c1782(
.A1(net894),
.A2(net934),
.ZN(net1863)
);

INV_X32 c1783(
.A(net9650),
.ZN(net1864)
);

NOR2_X4 c1784(
.A1(net1715),
.A2(net1846),
.ZN(net1865)
);

OR3_X4 c1785(
.A1(net1846),
.A2(net1829),
.A3(net861),
.ZN(net1866)
);

NOR2_X2 c1786(
.A1(net1866),
.A2(net1837),
.ZN(net1867)
);

XOR2_X2 c1787(
.A(net1855),
.B(net848),
.Z(net1868)
);

AND3_X2 c1788(
.A1(net1856),
.A2(net1841),
.A3(net1849),
.ZN(net1869)
);

XNOR2_X1 c1789(
.A(net1861),
.B(net1837),
.ZN(net1870)
);

OR2_X4 c1790(
.A1(net698),
.A2(net1830),
.ZN(net1871)
);

OR2_X1 c1791(
.A1(net889),
.A2(net11061),
.ZN(net1872)
);

XNOR2_X2 c1792(
.A(net1848),
.B(net849),
.ZN(net1873)
);

AND2_X4 c1793(
.A1(net901),
.A2(net10929),
.ZN(net1874)
);

AND2_X1 c1794(
.A1(net1862),
.A2(net1849),
.ZN(net1875)
);

NAND2_X1 c1795(
.A1(net1758),
.A2(net1755),
.ZN(net1876)
);

NOR3_X1 c1796(
.A1(net911),
.A2(net940),
.A3(net1857),
.ZN(net1877)
);

NAND2_X2 c1797(
.A1(net1821),
.A2(net823),
.ZN(net1878)
);

NAND2_X4 c1798(
.A1(net1842),
.A2(net11061),
.ZN(net1879)
);

AND2_X2 c1799(
.A1(net766),
.A2(net1841),
.ZN(net1880)
);

INV_X4 c1800(
.A(net10060),
.ZN(net1881)
);

OAI222_X1 c1801(
.A1(net1845),
.A2(net938),
.B1(net876),
.B2(net863),
.C1(net1824),
.C2(net10990),
.ZN(net1882)
);

XOR2_X1 c1802(
.A(net1875),
.B(net1842),
.Z(net1883)
);

OR3_X2 c1803(
.A1(net1854),
.A2(net1518),
.A3(net1868),
.ZN(net1884)
);

DFFR_X1 c1804(
.D(net1849),
.RN(net1755),
.CK(clk),
.Q(net1886),
.QN(net1885)
);

DFFRS_X2 c1805(
.D(net940),
.RN(net1880),
.SN(net1844),
.CK(clk),
.Q(net1888),
.QN(net1887)
);

OAI21_X2 c1806(
.A(net1878),
.B1(net1866),
.B2(net927),
.ZN(net1889)
);

NOR2_X1 c1807(
.A1(net1518),
.A2(net1872),
.ZN(net1890)
);

OAI21_X1 c1808(
.A(net1883),
.B1(net1814),
.B2(net1885),
.ZN(net1891)
);

SDFF_X1 c1809(
.D(net1891),
.SE(net907),
.SI(net1880),
.CK(clk),
.Q(net1893),
.QN(net1892)
);

AOI21_X2 c1810(
.A(net935),
.B1(net1890),
.B2(net10774),
.ZN(net1894)
);

AOI221_X2 c1811(
.A(net1859),
.B1(net1824),
.B2(net1890),
.C1(net914),
.C2(net876),
.ZN(net1895)
);

AOI21_X1 c1812(
.A(net1879),
.B1(net1892),
.B2(net11267),
.ZN(net1896)
);

AOI21_X4 c1813(
.A(net1894),
.B1(net1888),
.B2(net1881),
.ZN(net1897)
);

OR2_X2 c1814(
.A1(net1894),
.A2(net10996),
.ZN(net1898)
);

OAI22_X1 c1815(
.A1(net1896),
.A2(net1837),
.B1(net1887),
.B2(net876),
.ZN(net1899)
);

NOR2_X4 c1816(
.A1(net1872),
.A2(net1758),
.ZN(net1900)
);

NOR2_X2 c1817(
.A1(net1900),
.A2(net1846),
.ZN(net1901)
);

AND4_X2 c1818(
.A1(net1899),
.A2(net1852),
.A3(net1833),
.A4(net1870),
.ZN(net1902)
);

XOR2_X2 c1819(
.A(net1836),
.B(net11508),
.Z(net1903)
);

AOI221_X1 c1820(
.A(net1823),
.B1(net894),
.B2(net1886),
.C1(net1829),
.C2(net876),
.ZN(net1904)
);

XNOR2_X1 c1821(
.A(net865),
.B(net1868),
.ZN(net1905)
);

OR2_X4 c1822(
.A1(net1904),
.A2(net10804),
.ZN(net1906)
);

AND4_X1 c1823(
.A1(net1890),
.A2(net1902),
.A3(net1881),
.A4(net1840),
.ZN(net1907)
);

SDFF_X2 c1824(
.D(net1907),
.SE(net1904),
.SI(net11267),
.CK(clk),
.Q(net1909),
.QN(net1908)
);

DFFRS_X1 c1825(
.D(net1834),
.RN(net1908),
.SN(net10756),
.CK(clk),
.Q(net1911),
.QN(net1910)
);

INV_X1 c1826(
.A(net956),
.ZN(net1912)
);

INV_X2 c1827(
.A(net1912),
.ZN(net1913)
);

INV_X8 c1828(
.A(net15),
.ZN(net1914)
);

INV_X16 c1829(
.A(net1914),
.ZN(net1915)
);

INV_X32 c1830(
.A(net56),
.ZN(net1916)
);

INV_X4 c1831(
.A(net9799),
.ZN(net1917)
);

DFFR_X2 c1832(
.D(net943),
.RN(net954),
.CK(clk),
.Q(net1919),
.QN(net1918)
);

INV_X1 c1833(
.A(net7),
.ZN(net1920)
);

INV_X2 c1834(
.A(net1913),
.ZN(net1921)
);

INV_X8 c1835(
.A(net1920),
.ZN(net1922)
);

INV_X16 c1836(
.A(net1025),
.ZN(net1923)
);

INV_X32 c1837(
.A(net9798),
.ZN(net1924)
);

INV_X4 c1838(
.A(net993),
.ZN(net1925)
);

INV_X1 c1839(
.A(net1007),
.ZN(net1926)
);

OR2_X1 c1840(
.A1(net1009),
.A2(net1926),
.ZN(net1927)
);

INV_X2 c1841(
.A(net1924),
.ZN(net1928)
);

XNOR2_X2 c1842(
.A(net978),
.B(net1927),
.ZN(net1929)
);

INV_X8 c1843(
.A(net1919),
.ZN(net1930)
);

AND2_X4 c1844(
.A1(net968),
.A2(net1913),
.ZN(net1931)
);

AND3_X1 c1845(
.A1(net1924),
.A2(net7),
.A3(net10533),
.ZN(net1932)
);

INV_X16 c1846(
.A(net9879),
.ZN(net1933)
);

AND2_X1 c1847(
.A1(net1007),
.A2(net1920),
.ZN(net1934)
);

INV_X32 c1848(
.A(net947),
.ZN(net1935)
);

INV_X4 c1849(
.A(net56),
.ZN(net1936)
);

NAND3_X1 c1850(
.A1(net956),
.A2(net1930),
.A3(net996),
.ZN(net1937)
);

INV_X1 c1851(
.A(net1928),
.ZN(net1938)
);

NAND2_X1 c1852(
.A1(net980),
.A2(net1923),
.ZN(net1939)
);

NAND2_X2 c1853(
.A1(net969),
.A2(net1926),
.ZN(net1940)
);

NAND2_X4 c1854(
.A1(net1025),
.A2(net1923),
.ZN(net1941)
);

INV_X2 c1855(
.A(net21),
.ZN(net1942)
);

NOR3_X4 c1856(
.A1(net1936),
.A2(net1934),
.A3(net954),
.ZN(net1943)
);

NOR3_X2 c1857(
.A1(net1926),
.A2(net1012),
.A3(net29),
.ZN(net1944)
);

DFFS_X1 c1858(
.D(net1941),
.SN(net1918),
.CK(clk),
.Q(net1946),
.QN(net1945)
);

AND2_X2 c1859(
.A1(net1923),
.A2(net1945),
.ZN(net1947)
);

INV_X8 c1860(
.A(net9993),
.ZN(net1948)
);

DFFRS_X2 c1861(
.D(net1925),
.RN(net1916),
.SN(net1019),
.CK(clk),
.Q(net1950),
.QN(net1949)
);

INV_X16 c1862(
.A(net1950),
.ZN(net1951)
);

XOR2_X1 c1863(
.A(net1940),
.B(net10532),
.Z(net1952)
);

DFFS_X2 c1864(
.D(net1939),
.SN(net1948),
.CK(clk),
.Q(net1954),
.QN(net1953)
);

DFFR_X1 c1865(
.D(net1913),
.RN(net1947),
.CK(clk),
.Q(net1956),
.QN(net1955)
);

INV_X32 c1866(
.A(net9994),
.ZN(net1957)
);

NOR2_X1 c1867(
.A1(net1942),
.A2(net1948),
.ZN(net1958)
);

INV_X4 c1868(
.A(net1931),
.ZN(net1959)
);

INV_X1 c1869(
.A(net993),
.ZN(net1960)
);

OR2_X2 c1870(
.A1(net1937),
.A2(net949),
.ZN(net1961)
);

INV_X2 c1871(
.A(net1938),
.ZN(net1962)
);

NOR2_X4 c1872(
.A1(net1917),
.A2(net947),
.ZN(net1963)
);

NOR2_X2 c1873(
.A1(net1934),
.A2(net1007),
.ZN(net1964)
);

INV_X8 c1874(
.A(net1912),
.ZN(net1965)
);

DFFR_X2 c1875(
.D(net1941),
.RN(net1016),
.CK(clk),
.Q(net1967),
.QN(net1966)
);

XOR2_X2 c1876(
.A(net1953),
.B(net1963),
.Z(net1968)
);

XNOR2_X1 c1877(
.A(net1963),
.B(net1928),
.ZN(net1969)
);

AND3_X4 c1878(
.A1(net982),
.A2(net1963),
.A3(net1926),
.ZN(net1970)
);

INV_X16 c1879(
.A(net9861),
.ZN(net1971)
);

DFFS_X1 c1880(
.D(net1965),
.SN(net1970),
.CK(clk),
.Q(net1973),
.QN(net1972)
);

NAND3_X2 c1881(
.A1(net1948),
.A2(net1928),
.A3(net1011),
.ZN(net1974)
);

INV_X32 c1882(
.A(net1969),
.ZN(net1975)
);

DFFS_X2 c1883(
.D(net1960),
.SN(net1945),
.CK(clk),
.Q(net1977),
.QN(net1976)
);

DFFR_X1 c1884(
.D(net1925),
.RN(net1976),
.CK(clk),
.Q(net1979),
.QN(net1978)
);

OR2_X4 c1885(
.A1(net1975),
.A2(net1937),
.ZN(net1980)
);

INV_X4 c1886(
.A(net1969),
.ZN(net1981)
);

INV_X1 c1887(
.A(net1971),
.ZN(net1982)
);

OR2_X1 c1888(
.A1(net1919),
.A2(net1948),
.ZN(net1983)
);

XNOR2_X2 c1889(
.A(net1935),
.B(net1938),
.ZN(net1984)
);

AND2_X4 c1890(
.A1(net1983),
.A2(net1980),
.ZN(net1985)
);

OR3_X1 c1891(
.A1(net1984),
.A2(net1975),
.A3(net1012),
.ZN(net1986)
);

DFFR_X2 c1892(
.D(net1012),
.RN(net1964),
.CK(clk),
.Q(net1988),
.QN(net1987)
);

DFFS_X1 c1893(
.D(net1964),
.SN(net1957),
.CK(clk),
.Q(net1990),
.QN(net1989)
);

AND2_X1 c1894(
.A1(net1990),
.A2(net1966),
.ZN(net1991)
);

OAI221_X1 c1895(
.A(net972),
.B1(net1986),
.B2(net56),
.C1(net1961),
.C2(net45),
.ZN(net1992)
);

MUX2_X1 c1896(
.A(net1962),
.B(net1949),
.S(net10711),
.Z(net1993)
);

SDFF_X1 c1897(
.D(net1981),
.SE(net1947),
.SI(net1993),
.CK(clk),
.Q(net1995),
.QN(net1994)
);

NAND2_X1 c1898(
.A1(net21),
.A2(net1981),
.ZN(net1996)
);

SDFF_X2 c1899(
.D(net1967),
.SE(net1995),
.SI(net1941),
.CK(clk),
.Q(net1998),
.QN(net1997)
);

OAI21_X4 c1900(
.A(net1997),
.B1(net1968),
.B2(net10866),
.ZN(net1999)
);

DFFS_X2 c1901(
.D(net1916),
.SN(net1960),
.CK(clk),
.Q(net2001),
.QN(net2000)
);

DFFRS_X1 c1902(
.D(net1998),
.RN(net1985),
.SN(net1996),
.CK(clk),
.Q(net2003),
.QN(net2002)
);

NAND2_X2 c1903(
.A1(net1985),
.A2(net2003),
.ZN(net2004)
);

DFFRS_X2 c1904(
.D(net1954),
.RN(net1983),
.SN(net1986),
.CK(clk),
.Q(net2006),
.QN(net2005)
);

NAND2_X4 c1905(
.A1(net1957),
.A2(net10699),
.ZN(net2007)
);

OAI222_X4 c1906(
.A1(in25),
.A2(net1983),
.B1(net2002),
.B2(net954),
.C1(net966),
.C2(net1922),
.ZN(net2008)
);

MUX2_X2 c1907(
.A(net1962),
.B(net1977),
.S(net2007),
.Z(net2009)
);

AOI22_X4 c1908(
.A1(net2003),
.A2(net1999),
.B1(net2009),
.B2(net1944),
.ZN(net2010)
);

INV_X2 c1909(
.A(net1102),
.ZN(net2011)
);

AND2_X2 c1910(
.A1(net45),
.A2(net57),
.ZN(net2012)
);

INV_X8 c1911(
.A(net1963),
.ZN(net2013)
);

XOR2_X1 c1912(
.A(net2007),
.B(net1050),
.Z(net2014)
);

INV_X16 c1913(
.A(net102),
.ZN(net2015)
);

INV_X32 c1914(
.A(net2013),
.ZN(net2016)
);

INV_X4 c1915(
.A(net118),
.ZN(net2017)
);

NOR2_X1 c1916(
.A1(net2014),
.A2(net11501),
.ZN(net2018)
);

INV_X1 c1917(
.A(net9809),
.ZN(net2019)
);

OR2_X2 c1918(
.A1(net966),
.A2(net2007),
.ZN(net2020)
);

INV_X2 c1919(
.A(net9718),
.ZN(net2021)
);

NOR2_X4 c1920(
.A1(net2021),
.A2(net1115),
.ZN(net2022)
);

INV_X8 c1921(
.A(net9717),
.ZN(net2023)
);

INV_X16 c1922(
.A(net1958),
.ZN(net2024)
);

INV_X32 c1923(
.A(net2001),
.ZN(net2025)
);

INV_X4 c1924(
.A(net2015),
.ZN(net2026)
);

INV_X1 c1925(
.A(net2009),
.ZN(net2027)
);

SDFF_X1 c1926(
.D(net102),
.SE(net1091),
.SI(net2018),
.CK(clk),
.Q(net2029),
.QN(net2028)
);

INV_X2 c1927(
.A(net9831),
.ZN(net2030)
);

NOR2_X2 c1928(
.A1(net1991),
.A2(net2025),
.ZN(net2031)
);

XOR2_X2 c1929(
.A(net1091),
.B(net1958),
.Z(net2032)
);

INV_X8 c1930(
.A(net9832),
.ZN(net2033)
);

INV_X16 c1931(
.A(net9832),
.ZN(net2034)
);

XNOR2_X1 c1932(
.A(net2014),
.B(net996),
.ZN(net2035)
);

OR2_X4 c1933(
.A1(net1090),
.A2(net45),
.ZN(net2036)
);

INV_X32 c1934(
.A(net1977),
.ZN(net2037)
);

OR2_X1 c1935(
.A1(net2017),
.A2(net2000),
.ZN(net2038)
);

INV_X4 c1936(
.A(net996),
.ZN(net2039)
);

DFFR_X1 c1937(
.D(net1090),
.RN(net2038),
.CK(clk),
.Q(net2041),
.QN(net2040)
);

INV_X1 c1938(
.A(net10303),
.ZN(net2042)
);

INV_X2 c1939(
.A(net2024),
.ZN(net2043)
);

INV_X8 c1940(
.A(net10057),
.ZN(net2044)
);

NAND3_X4 c1941(
.A1(net2039),
.A2(net2043),
.A3(net1041),
.ZN(net2045)
);

OR3_X4 c1942(
.A1(net2012),
.A2(net2031),
.A3(net1996),
.ZN(net2046)
);

INV_X16 c1943(
.A(net2019),
.ZN(net2047)
);

INV_X32 c1944(
.A(net2018),
.ZN(net2048)
);

XNOR2_X2 c1945(
.A(net1926),
.B(net87),
.ZN(net2049)
);

SDFF_X2 c1946(
.D(net2025),
.SE(net1940),
.SI(net10700),
.CK(clk),
.Q(net2051),
.QN(net2050)
);

INV_X4 c1947(
.A(net2036),
.ZN(net2052)
);

INV_X1 c1948(
.A(net2045),
.ZN(net2053)
);

INV_X2 c1949(
.A(net1115),
.ZN(net2054)
);

AND2_X4 c1950(
.A1(net2034),
.A2(net2015),
.ZN(net2055)
);

AND3_X2 c1951(
.A1(net990),
.A2(net2013),
.A3(net1991),
.ZN(net2056)
);

INV_X8 c1952(
.A(net2035),
.ZN(net2057)
);

INV_X16 c1953(
.A(net2036),
.ZN(net2058)
);

INV_X32 c1954(
.A(net1008),
.ZN(net2059)
);

INV_X4 c1955(
.A(net10134),
.ZN(net2060)
);

INV_X1 c1956(
.A(net2031),
.ZN(net2061)
);

AND2_X1 c1957(
.A1(net2061),
.A2(net10866),
.ZN(net2062)
);

INV_X2 c1958(
.A(net1921),
.ZN(net2063)
);

DFFR_X2 c1959(
.D(net2055),
.RN(net1024),
.CK(clk),
.Q(net2065),
.QN(net2064)
);

INV_X8 c1960(
.A(net1041),
.ZN(net2066)
);

NOR3_X1 c1961(
.A1(net2060),
.A2(net1090),
.A3(net1976),
.ZN(net2067)
);

DFFS_X1 c1962(
.D(net2043),
.SN(net1944),
.CK(clk),
.Q(net2069),
.QN(net2068)
);

NAND2_X1 c1963(
.A1(net2016),
.A2(net2025),
.ZN(net2070)
);

NAND2_X2 c1964(
.A1(net2063),
.A2(net2066),
.ZN(net2071)
);

INV_X16 c1965(
.A(net2039),
.ZN(net2072)
);

NAND2_X4 c1966(
.A1(net2025),
.A2(net2064),
.ZN(net2073)
);

AND2_X2 c1967(
.A1(net1102),
.A2(net2028),
.ZN(net2074)
);

XOR2_X1 c1968(
.A(net2065),
.B(net2046),
.Z(net2075)
);

NOR2_X1 c1969(
.A1(net2059),
.A2(net2068),
.ZN(net2076)
);

INV_X32 c1970(
.A(net2046),
.ZN(net2077)
);

INV_X4 c1971(
.A(net10893),
.ZN(net2078)
);

DFFS_X2 c1972(
.D(net2075),
.SN(net2011),
.CK(clk),
.Q(net2080),
.QN(net2079)
);

OR2_X2 c1973(
.A1(net2011),
.A2(net2068),
.ZN(net2081)
);

OR3_X2 c1974(
.A1(net2049),
.A2(net2079),
.A3(net2074),
.ZN(net2082)
);

NOR2_X4 c1975(
.A1(net2070),
.A2(net2072),
.ZN(net2083)
);

NOR2_X2 c1976(
.A1(net2074),
.A2(net2068),
.ZN(net2084)
);

DFFR_X1 c1977(
.D(net2054),
.RN(net2067),
.CK(clk),
.Q(net2086),
.QN(net2085)
);

OAI21_X2 c1978(
.A(net2037),
.B1(net2081),
.B2(net966),
.ZN(net2087)
);

OAI21_X1 c1979(
.A(net2026),
.B1(net2065),
.B2(net1993),
.ZN(net2088)
);

XOR2_X2 c1980(
.A(net2080),
.B(net10932),
.Z(net2089)
);

OAI222_X2 c1981(
.A1(net2087),
.A2(net2078),
.B1(net2014),
.B2(net1932),
.C1(net1035),
.C2(net2016),
.ZN(net2090)
);

XNOR2_X1 c1982(
.A(net2030),
.B(net2086),
.ZN(net2091)
);

AOI21_X2 c1983(
.A(net2084),
.B1(net2090),
.B2(net2067),
.ZN(net2092)
);

AOI21_X1 c1984(
.A(net1040),
.B1(net2090),
.B2(net2064),
.ZN(net2093)
);

AOI21_X4 c1985(
.A(net124),
.B1(net2085),
.B2(net2088),
.ZN(net2094)
);

OR2_X4 c1986(
.A1(net2093),
.A2(net1112),
.ZN(net2095)
);

OR2_X1 c1987(
.A1(net2073),
.A2(net2088),
.ZN(net2096)
);

XNOR2_X2 c1988(
.A(net2062),
.B(net2095),
.ZN(net2097)
);

AND3_X1 c1989(
.A1(net2012),
.A2(net2096),
.A3(net2088),
.ZN(net2098)
);

NAND3_X1 c1990(
.A1(net2053),
.A2(net2098),
.A3(net11501),
.ZN(net2099)
);

NOR3_X4 c1991(
.A1(net2098),
.A2(net2086),
.A3(net10622),
.ZN(net2100)
);

INV_X1 c1992(
.A(net2181),
.ZN(net2101)
);

INV_X2 c1993(
.A(net2007),
.ZN(net2102)
);

INV_X8 c1994(
.A(net1142),
.ZN(net2103)
);

INV_X16 c1995(
.A(net2186),
.ZN(net2104)
);

DFFR_X2 c1996(
.D(net2176),
.RN(net1144),
.CK(clk),
.Q(net2106),
.QN(net2105)
);

INV_X32 c1997(
.A(net1161),
.ZN(net2107)
);

INV_X4 c1998(
.A(net10474),
.ZN(net2108)
);

AND2_X4 c1999(
.A1(net2105),
.A2(net10821),
.ZN(net2109)
);

INV_X1 c2000(
.A(net1189),
.ZN(net2110)
);

NOR3_X2 c2001(
.A1(net2110),
.A2(net2102),
.A3(net1961),
.ZN(net2111)
);

AND2_X1 c2002(
.A1(net2108),
.A2(net2169),
.ZN(net2112)
);

NAND2_X1 c2003(
.A1(net2111),
.A2(net214),
.ZN(net2113)
);

INV_X2 c2004(
.A(net9673),
.ZN(net2114)
);

INV_X8 c2005(
.A(net9673),
.ZN(net2115)
);

OAI221_X4 c2006(
.A(net1128),
.B1(net1162),
.B2(net2107),
.C1(net2161),
.C2(net191),
.ZN(net2116)
);

NAND2_X2 c2007(
.A1(net2186),
.A2(net2181),
.ZN(net2117)
);

INV_X16 c2008(
.A(net2101),
.ZN(net2118)
);

INV_X32 c2009(
.A(net9831),
.ZN(net2119)
);

NAND2_X4 c2010(
.A1(net2112),
.A2(net2119),
.ZN(net2120)
);

OAI221_X2 c2011(
.A(net2118),
.B1(net118),
.B2(net236),
.C1(net1100),
.C2(net2161),
.ZN(net2121)
);

AND2_X2 c2012(
.A1(net2115),
.A2(net1996),
.ZN(net2122)
);

AND3_X4 c2013(
.A1(net2102),
.A2(net1141),
.A3(net1951),
.ZN(net2123)
);

XOR2_X1 c2014(
.A(net2117),
.B(net2109),
.Z(net2124)
);

NOR2_X1 c2015(
.A1(net2166),
.A2(net2119),
.ZN(net2125)
);

NAND3_X2 c2016(
.A1(net2091),
.A2(net2117),
.A3(net1165),
.ZN(net2126)
);

INV_X4 c2017(
.A(net10176),
.ZN(net2127)
);

OR2_X2 c2018(
.A1(net2173),
.A2(net1993),
.ZN(net2128)
);

OR3_X1 c2019(
.A1(net2124),
.A2(net2112),
.A3(net1101),
.ZN(net2129)
);

NOR2_X4 c2020(
.A1(net2119),
.A2(net2186),
.ZN(net2130)
);

NOR2_X2 c2021(
.A1(net1177),
.A2(net2110),
.ZN(net2131)
);

XOR2_X2 c2022(
.A(net2128),
.B(net2174),
.Z(net2132)
);

INV_X1 c2023(
.A(net2120),
.ZN(net2133)
);

INV_X2 c2024(
.A(net2133),
.ZN(net2134)
);

XNOR2_X1 c2025(
.A(net2121),
.B(net2127),
.ZN(net2135)
);

MUX2_X1 c2026(
.A(net2123),
.B(net2128),
.S(net11047),
.Z(net2136)
);

OR2_X4 c2027(
.A1(net2057),
.A2(net1185),
.ZN(net2137)
);

OAI21_X4 c2028(
.A(net1144),
.B1(net2128),
.B2(net2174),
.ZN(net2138)
);

INV_X8 c2029(
.A(net2131),
.ZN(net2139)
);

INV_X16 c2030(
.A(net2106),
.ZN(net2140)
);

OR2_X1 c2031(
.A1(net2182),
.A2(net2112),
.ZN(net2141)
);

INV_X32 c2032(
.A(net10083),
.ZN(net2142)
);

MUX2_X2 c2033(
.A(net2123),
.B(net2120),
.S(net1047),
.Z(net2143)
);

INV_X4 c2034(
.A(net9910),
.ZN(net2144)
);

DFFRS_X1 c2035(
.D(net2137),
.RN(net2139),
.SN(net1177),
.CK(clk),
.Q(net2146),
.QN(net2145)
);

NAND3_X4 c2036(
.A1(net2109),
.A2(net2141),
.A3(net2179),
.ZN(net2147)
);

OAI22_X4 c2037(
.A1(net1135),
.A2(net2146),
.B1(net2129),
.B2(net2179),
.ZN(net2148)
);

XNOR2_X2 c2038(
.A(net2132),
.B(net2146),
.ZN(net2149)
);

OR3_X4 c2039(
.A1(net2138),
.A2(net2106),
.A3(net2040),
.ZN(net2150)
);

AND2_X4 c2040(
.A1(net214),
.A2(net2141),
.ZN(net2151)
);

AND3_X2 c2041(
.A1(net1101),
.A2(net2101),
.A3(net11398),
.ZN(net2152)
);

NOR3_X1 c2042(
.A1(net2130),
.A2(net57),
.A3(net11271),
.ZN(net2153)
);

OR3_X2 c2043(
.A1(net2136),
.A2(net2152),
.A3(net11271),
.ZN(net2154)
);

SDFFRS_X2 c2044(
.D(net2114),
.RN(net2143),
.SE(net1959),
.SI(net1190),
.SN(net1107),
.CK(clk),
.Q(net2156),
.QN(net2155)
);

AOI22_X2 c2045(
.A1(net2140),
.A2(net2178),
.B1(net2155),
.B2(net2153),
.ZN(net2157)
);

AND2_X1 c2046(
.A1(net2134),
.A2(net2156),
.ZN(net2158)
);

AOI221_X4 c2047(
.A(net2156),
.B1(net2121),
.B2(net1204),
.C1(net2158),
.C2(net124),
.ZN(net2159)
);

AOI221_X2 c2048(
.A(net2129),
.B1(net1202),
.B2(net2155),
.C1(net2158),
.C2(net2016),
.ZN(net2160)
);

INV_X1 c2049(
.A(net1150),
.ZN(net2161)
);

OAI21_X2 c2050(
.A(net2097),
.B1(net1169),
.B2(net1915),
.ZN(net2162)
);

INV_X2 c2051(
.A(net9992),
.ZN(net2163)
);

NAND2_X1 c2052(
.A1(net1127),
.A2(net213),
.ZN(net2164)
);

INV_X8 c2053(
.A(net9951),
.ZN(net2165)
);

INV_X16 c2054(
.A(net1205),
.ZN(net2166)
);

INV_X32 c2055(
.A(net11418),
.ZN(net2167)
);

OAI21_X1 c2056(
.A(net1162),
.B1(net1206),
.B2(net1144),
.ZN(net2168)
);

INV_X4 c2057(
.A(net1159),
.ZN(net2169)
);

AOI221_X1 c2058(
.A(net212),
.B1(net1961),
.B2(net2078),
.C1(net1160),
.C2(net2169),
.ZN(net2170)
);

INV_X1 c2059(
.A(net2169),
.ZN(net2171)
);

NAND2_X2 c2060(
.A1(net1107),
.A2(net1128),
.ZN(net2172)
);

NAND2_X4 c2061(
.A1(net1067),
.A2(net2169),
.ZN(net2173)
);

AND2_X2 c2062(
.A1(net1191),
.A2(net2161),
.ZN(net2174)
);

AOI21_X2 c2063(
.A(net87),
.B1(net1188),
.B2(net2171),
.ZN(net2175)
);

XOR2_X1 c2064(
.A(net2174),
.B(net2061),
.Z(net2176)
);

INV_X2 c2065(
.A(net2175),
.ZN(net2177)
);

NOR2_X1 c2066(
.A1(net2175),
.A2(net1142),
.ZN(net2178)
);

OR2_X2 c2067(
.A1(net2165),
.A2(net1993),
.ZN(net2179)
);

NOR2_X4 c2068(
.A1(net1164),
.A2(net2177),
.ZN(net2180)
);

INV_X8 c2069(
.A(net9816),
.ZN(net2181)
);

INV_X16 c2070(
.A(net2177),
.ZN(net2182)
);

NOR2_X2 c2071(
.A1(net2161),
.A2(net2164),
.ZN(net2183)
);

AOI21_X1 c2072(
.A(net1165),
.B1(net1993),
.B2(net2007),
.ZN(net2184)
);

INV_X32 c2073(
.A(net10257),
.ZN(net2185)
);

INV_X4 c2074(
.A(net10175),
.ZN(net2186)
);

INV_X1 c2075(
.A(net10959),
.ZN(net2187)
);

INV_X2 c2076(
.A(net237),
.ZN(net2188)
);

INV_X8 c2077(
.A(net11207),
.ZN(net2189)
);

XOR2_X2 c2078(
.A(net1264),
.B(net1151),
.Z(net2190)
);

XNOR2_X1 c2079(
.A(net2190),
.B(net2144),
.ZN(net2191)
);

INV_X16 c2080(
.A(net314),
.ZN(net2192)
);

OR2_X4 c2081(
.A1(net1065),
.A2(net1288),
.ZN(net2193)
);

INV_X32 c2082(
.A(net2110),
.ZN(net2194)
);

INV_X4 c2083(
.A(net1236),
.ZN(net2195)
);

INV_X1 c2084(
.A(net1259),
.ZN(net2196)
);

AOI21_X4 c2085(
.A(net2104),
.B1(net2041),
.B2(net2139),
.ZN(net2197)
);

OR2_X1 c2086(
.A1(net1153),
.A2(net1922),
.ZN(net2198)
);

INV_X2 c2087(
.A(net2194),
.ZN(net2199)
);

INV_X8 c2088(
.A(net2190),
.ZN(net2200)
);

INV_X16 c2089(
.A(net2152),
.ZN(net2201)
);

INV_X32 c2090(
.A(net1186),
.ZN(net2202)
);

INV_X4 c2091(
.A(net1291),
.ZN(net2203)
);

XNOR2_X2 c2092(
.A(net1262),
.B(net2187),
.ZN(net2204)
);

INV_X1 c2093(
.A(net2192),
.ZN(net2205)
);

INV_X2 c2094(
.A(net2041),
.ZN(net2206)
);

INV_X8 c2095(
.A(net10302),
.ZN(net2207)
);

INV_X16 c2096(
.A(net11207),
.ZN(net2208)
);

DFFRS_X2 c2097(
.D(net1272),
.RN(net2158),
.SN(net317),
.CK(clk),
.Q(net2210),
.QN(net2209)
);

AND2_X4 c2098(
.A1(net2103),
.A2(net70),
.ZN(net2211)
);

DFFS_X1 c2099(
.D(net1206),
.SN(net2169),
.CK(clk),
.Q(net2213),
.QN(net2212)
);

AND2_X1 c2100(
.A1(net2205),
.A2(net2028),
.ZN(net2214)
);

INV_X32 c2101(
.A(net2107),
.ZN(net2215)
);

INV_X4 c2102(
.A(net2195),
.ZN(net2216)
);

NAND2_X1 c2103(
.A1(net1293),
.A2(net2201),
.ZN(net2217)
);

INV_X1 c2104(
.A(net2211),
.ZN(net2218)
);

AOI222_X1 c2105(
.A1(net2218),
.A2(net2205),
.B1(net2199),
.B2(net2107),
.C1(net1225),
.C2(net1217),
.ZN(net2219)
);

INV_X2 c2106(
.A(net1279),
.ZN(net2220)
);

NAND2_X2 c2107(
.A1(net2217),
.A2(net10959),
.ZN(net2221)
);

NAND2_X4 c2108(
.A1(net1230),
.A2(net1086),
.ZN(net2222)
);

AND2_X2 c2109(
.A1(net1915),
.A2(net2188),
.ZN(net2223)
);

XOR2_X1 c2110(
.A(net2215),
.B(net2202),
.Z(net2224)
);

NOR2_X1 c2111(
.A1(net2201),
.A2(net2047),
.ZN(net2225)
);

OR2_X2 c2112(
.A1(net2225),
.A2(net2212),
.ZN(net2226)
);

INV_X8 c2113(
.A(net11157),
.ZN(net2227)
);

AND3_X1 c2114(
.A1(net2216),
.A2(net2206),
.A3(net2158),
.ZN(net2228)
);

INV_X16 c2115(
.A(net9850),
.ZN(net2229)
);

INV_X32 c2116(
.A(net11093),
.ZN(net2230)
);

NOR2_X4 c2117(
.A1(net2163),
.A2(net314),
.ZN(net2231)
);

NOR2_X2 c2118(
.A1(net2229),
.A2(net2223),
.ZN(net2232)
);

NAND3_X1 c2119(
.A1(net2047),
.A2(net1959),
.A3(net10827),
.ZN(net2233)
);

INV_X4 c2120(
.A(net2207),
.ZN(net2234)
);

INV_X1 c2121(
.A(net2200),
.ZN(net2235)
);

INV_X2 c2122(
.A(net2188),
.ZN(net2236)
);

XOR2_X2 c2123(
.A(net1240),
.B(net2235),
.Z(net2237)
);

NOR3_X4 c2124(
.A1(net254),
.A2(net1240),
.A3(net314),
.ZN(net2238)
);

NAND4_X4 c2125(
.A1(net2219),
.A2(net2208),
.A3(net1264),
.A4(net2016),
.ZN(net2239)
);

XNOR2_X1 c2126(
.A(net2238),
.B(net10960),
.ZN(net2240)
);

OAI211_X2 c2127(
.A(net315),
.B(net2235),
.C1(net2208),
.C2(net2192),
.ZN(net2241)
);

OR2_X4 c2128(
.A1(net2232),
.A2(net2192),
.ZN(net2242)
);

SDFF_X1 c2129(
.D(net1241),
.SE(net2219),
.SI(net2238),
.CK(clk),
.Q(net2244),
.QN(net2243)
);

INV_X8 c2130(
.A(net11270),
.ZN(net2245)
);

INV_X16 c2131(
.A(net10858),
.ZN(net2246)
);

DFFS_X2 c2132(
.D(net2244),
.SN(net1195),
.CK(clk),
.Q(net2248),
.QN(net2247)
);

OR2_X1 c2133(
.A1(net2245),
.A2(net2195),
.ZN(net2249)
);

XNOR2_X2 c2134(
.A(net2226),
.B(net2240),
.ZN(net2250)
);

OR4_X2 c2135(
.A1(net2210),
.A2(net2237),
.A3(net1263),
.A4(net2240),
.ZN(net2251)
);

AND2_X4 c2136(
.A1(net2214),
.A2(net2248),
.ZN(net2252)
);

AND2_X1 c2137(
.A1(net2222),
.A2(net2252),
.ZN(net2253)
);

NOR3_X2 c2138(
.A1(net2202),
.A2(net2243),
.A3(net2179),
.ZN(net2254)
);

AND3_X4 c2139(
.A1(net2250),
.A2(net2240),
.A3(net2229),
.ZN(net2255)
);

SDFF_X2 c2140(
.D(net2246),
.SE(net2252),
.SI(net1206),
.CK(clk),
.Q(net2257),
.QN(net2256)
);

NAND3_X2 c2141(
.A1(net2230),
.A2(net2220),
.A3(net2145),
.ZN(net2258)
);

NAND2_X1 c2142(
.A1(net2223),
.A2(net2250),
.ZN(net2259)
);

NAND2_X2 c2143(
.A1(net1255),
.A2(net2157),
.ZN(net2260)
);

NAND2_X4 c2144(
.A1(net2242),
.A2(net2259),
.ZN(net2261)
);

OR3_X1 c2145(
.A1(net290),
.A2(net2249),
.A3(net2241),
.ZN(net2262)
);

MUX2_X1 c2146(
.A(net2206),
.B(net2251),
.S(net2257),
.Z(net2263)
);

OAI21_X4 c2147(
.A(net2249),
.B1(net1959),
.B2(net11335),
.ZN(net2264)
);

AND2_X2 c2148(
.A1(net2253),
.A2(net2104),
.ZN(net2265)
);

XOR2_X1 c2149(
.A(net2208),
.B(net11101),
.Z(net2266)
);

MUX2_X2 c2150(
.A(net2249),
.B(net2237),
.S(net2188),
.Z(net2267)
);

NOR2_X1 c2151(
.A1(net2251),
.A2(net2210),
.ZN(net2268)
);

OR2_X2 c2152(
.A1(net2231),
.A2(net2107),
.ZN(net2269)
);

NOR2_X4 c2153(
.A1(net2268),
.A2(net2232),
.ZN(net2270)
);

DFFRS_X1 c2154(
.D(net2269),
.RN(net2266),
.SN(net2270),
.CK(clk),
.Q(net2272),
.QN(net2271)
);

NOR2_X2 c2155(
.A1(net1263),
.A2(net2218),
.ZN(net2273)
);

XOR2_X2 c2156(
.A(net1185),
.B(net2188),
.Z(net2274)
);

XNOR2_X1 c2157(
.A(net2273),
.B(net2209),
.ZN(net2275)
);

INV_X32 c2158(
.A(net2090),
.ZN(net2276)
);

INV_X4 c2159(
.A(net199),
.ZN(net2277)
);

OR2_X4 c2160(
.A1(net1358),
.A2(net334),
.ZN(net2278)
);

INV_X1 c2161(
.A(net33),
.ZN(net2279)
);

INV_X2 c2162(
.A(net2148),
.ZN(net2280)
);

INV_X8 c2163(
.A(net9699),
.ZN(net2281)
);

OR2_X1 c2164(
.A1(net1227),
.A2(net2236),
.ZN(net2282)
);

NAND3_X4 c2165(
.A1(net1280),
.A2(net2139),
.A3(net2279),
.ZN(net2283)
);

INV_X16 c2166(
.A(net2278),
.ZN(net2284)
);

XNOR2_X2 c2167(
.A(net2281),
.B(net1341),
.ZN(net2285)
);

DFFR_X1 c2168(
.D(net1375),
.RN(net2260),
.CK(clk),
.Q(net2287),
.QN(net2286)
);

AND2_X4 c2169(
.A1(net2277),
.A2(net11138),
.ZN(net2288)
);

AND2_X1 c2170(
.A1(net2275),
.A2(net290),
.ZN(net2289)
);

NAND2_X1 c2171(
.A1(net2248),
.A2(net377),
.ZN(net2290)
);

INV_X32 c2172(
.A(net11072),
.ZN(net2291)
);

NAND2_X2 c2173(
.A1(net2291),
.A2(net1316),
.ZN(net2292)
);

NAND2_X4 c2174(
.A1(net2280),
.A2(net1203),
.ZN(net2293)
);

AND2_X2 c2175(
.A1(net1350),
.A2(net1374),
.ZN(net2294)
);

INV_X4 c2176(
.A(net318),
.ZN(net2295)
);

XOR2_X1 c2177(
.A(net317),
.B(net10943),
.Z(net2296)
);

INV_X1 c2178(
.A(net9699),
.ZN(net2297)
);

NOR2_X1 c2179(
.A1(net2297),
.A2(net2296),
.ZN(net2298)
);

INV_X2 c2180(
.A(net1359),
.ZN(net2299)
);

OR2_X2 c2181(
.A1(net351),
.A2(net2276),
.ZN(net2300)
);

INV_X8 c2182(
.A(net10382),
.ZN(net2301)
);

OR3_X4 c2183(
.A1(net1214),
.A2(net1351),
.A3(net1190),
.ZN(net2302)
);

NOR2_X4 c2184(
.A1(net2187),
.A2(net1318),
.ZN(net2303)
);

NOR2_X2 c2185(
.A1(net2282),
.A2(net1350),
.ZN(net2304)
);

XOR2_X2 c2186(
.A(net2139),
.B(net2300),
.Z(net2305)
);

XNOR2_X1 c2187(
.A(net1307),
.B(net1318),
.ZN(net2306)
);

OR2_X4 c2188(
.A1(net2284),
.A2(net2304),
.ZN(net2307)
);

INV_X16 c2189(
.A(net10068),
.ZN(net2308)
);

INV_X32 c2190(
.A(net1254),
.ZN(net2309)
);

OR2_X1 c2191(
.A1(net1100),
.A2(net2301),
.ZN(net2310)
);

XNOR2_X2 c2192(
.A(net1318),
.B(net334),
.ZN(net2311)
);

INV_X4 c2193(
.A(net384),
.ZN(net2312)
);

AND2_X4 c2194(
.A1(net2307),
.A2(net1343),
.ZN(net2313)
);

INV_X1 c2195(
.A(net2289),
.ZN(net2314)
);

AND2_X1 c2196(
.A1(net2303),
.A2(net2280),
.ZN(net2315)
);

NAND2_X1 c2197(
.A1(net1369),
.A2(net2282),
.ZN(net2316)
);

NAND2_X2 c2198(
.A1(net2285),
.A2(net2236),
.ZN(net2317)
);

NAND2_X4 c2199(
.A1(net2298),
.A2(net2259),
.ZN(net2318)
);

AND2_X2 c2200(
.A1(net2315),
.A2(net2282),
.ZN(net2319)
);

XOR2_X1 c2201(
.A(net10943),
.B(net11110),
.Z(net2320)
);

AND3_X2 c2202(
.A1(net2303),
.A2(net2316),
.A3(net11068),
.ZN(net2321)
);

NOR2_X1 c2203(
.A1(net409),
.A2(net2320),
.ZN(net2322)
);

INV_X2 c2204(
.A(net10186),
.ZN(net2323)
);

NOR3_X1 c2205(
.A1(net2293),
.A2(net2314),
.A3(net2304),
.ZN(net2324)
);

OR2_X2 c2206(
.A1(net1333),
.A2(net2287),
.ZN(net2325)
);

SDFFRS_X1 c2207(
.D(net2204),
.RN(net2247),
.SE(net1310),
.SI(net2256),
.SN(net1379),
.CK(clk),
.Q(net2327),
.QN(net2326)
);

NOR2_X4 c2208(
.A1(net2295),
.A2(net2323),
.ZN(net2328)
);

AOI222_X4 c2209(
.A1(net1190),
.A2(net1361),
.B1(net2292),
.B2(net2301),
.C1(net2276),
.C2(net2280),
.ZN(net2329)
);

NOR2_X2 c2210(
.A1(net2321),
.A2(net11110),
.ZN(net2330)
);

XOR2_X2 c2211(
.A(net2047),
.B(net2304),
.Z(net2331)
);

XNOR2_X1 c2212(
.A(net1354),
.B(net2306),
.ZN(net2332)
);

OR2_X4 c2213(
.A1(net2213),
.A2(net2317),
.ZN(net2333)
);

OR2_X1 c2214(
.A1(net2325),
.A2(net2320),
.ZN(net2334)
);

SDFFRS_X2 c2215(
.D(net2331),
.RN(net2308),
.SE(net1348),
.SI(net408),
.SN(net11504),
.CK(clk),
.Q(net2336),
.QN(net2335)
);

OR3_X2 c2216(
.A1(net2309),
.A2(net1224),
.A3(net11468),
.ZN(net2337)
);

XNOR2_X2 c2217(
.A(net2303),
.B(net11344),
.ZN(net2338)
);

AND2_X4 c2218(
.A1(net334),
.A2(net1338),
.ZN(net2339)
);

AND2_X1 c2219(
.A1(net2322),
.A2(net2338),
.ZN(net2340)
);

OAI21_X2 c2220(
.A(net2301),
.B1(net2303),
.B2(net2276),
.ZN(net2341)
);

DFFRS_X2 c2221(
.D(net2305),
.RN(net2301),
.SN(net11060),
.CK(clk),
.Q(net2343),
.QN(net2342)
);

NAND2_X1 c2222(
.A1(net1224),
.A2(net2240),
.ZN(net2344)
);

NAND2_X2 c2223(
.A1(net377),
.A2(net2325),
.ZN(net2345)
);

NAND2_X4 c2224(
.A1(net1327),
.A2(net1247),
.ZN(net2346)
);

AND2_X2 c2225(
.A1(net2320),
.A2(net2287),
.ZN(net2347)
);

DFFR_X2 c2226(
.D(net2305),
.RN(net2325),
.CK(clk),
.Q(net2349),
.QN(net2348)
);

XOR2_X1 c2227(
.A(net2344),
.B(net2342),
.Z(net2350)
);

OAI21_X1 c2228(
.A(net2279),
.B1(net283),
.B2(net2334),
.ZN(net2351)
);

OAI33_X1 c2229(
.A1(net2343),
.A2(net1270),
.A3(net2320),
.B1(net1247),
.B2(net2280),
.B3(net1227),
.ZN(net2352)
);

AOI21_X2 c2230(
.A(net2292),
.B1(net1227),
.B2(net1375),
.ZN(net2353)
);

NOR2_X1 c2231(
.A1(net2353),
.A2(net2334),
.ZN(net2354)
);

AOI222_X2 c2232(
.A1(net2353),
.A2(net2335),
.B1(net2286),
.B2(net1086),
.C1(net2351),
.C2(net11047),
.ZN(net2355)
);

SDFF_X1 c2233(
.D(net2199),
.SE(net2321),
.SI(net2300),
.CK(clk),
.Q(net2357),
.QN(net2356)
);

SDFF_X2 c2234(
.D(net2158),
.SE(net2357),
.SI(net2354),
.CK(clk),
.Q(net2359),
.QN(net2358)
);

AOI21_X1 c2235(
.A(net2350),
.B1(net2359),
.B2(net2148),
.ZN(net2360)
);

AOI21_X4 c2236(
.A(net1348),
.B1(net2336),
.B2(net11357),
.ZN(net2361)
);

DFFRS_X1 c2237(
.D(net2352),
.RN(net2354),
.SN(net2090),
.CK(clk),
.Q(net2363),
.QN(net2362)
);

OAI222_X1 c2238(
.A1(net2360),
.A2(net2334),
.B1(net1369),
.B2(net2354),
.C1(net2335),
.C2(net2256),
.ZN(net2364)
);

AOI211_X1 c2239(
.A(net2167),
.B(net2328),
.C1(net2334),
.C2(net1310),
.ZN(net2365)
);

AND3_X1 c2240(
.A1(net1100),
.A2(net2354),
.A3(net11295),
.ZN(net2366)
);

INV_X8 c2241(
.A(net2300),
.ZN(net2367)
);

INV_X16 c2242(
.A(net11322),
.ZN(net2368)
);

INV_X32 c2243(
.A(net11043),
.ZN(net2369)
);

INV_X4 c2244(
.A(net2361),
.ZN(net2370)
);

OR2_X2 c2245(
.A1(net2310),
.A2(net2370),
.ZN(net2371)
);

NAND3_X1 c2246(
.A1(net2260),
.A2(net2310),
.A3(net2356),
.ZN(net2372)
);

INV_X1 c2247(
.A(net2334),
.ZN(net2373)
);

NOR3_X4 c2248(
.A1(net1423),
.A2(net1379),
.A3(net357),
.ZN(net2374)
);

OAI221_X1 c2249(
.A(net2339),
.B1(net2373),
.B2(net2257),
.C1(net1401),
.C2(net1428),
.ZN(net2375)
);

NOR2_X4 c2250(
.A1(net2349),
.A2(net432),
.ZN(net2376)
);

INV_X2 c2251(
.A(net11286),
.ZN(net2377)
);

NOR3_X2 c2252(
.A1(net2259),
.A2(net1428),
.A3(net1466),
.ZN(net2378)
);

NOR2_X2 c2253(
.A1(net1403),
.A2(net11060),
.ZN(net2379)
);

INV_X8 c2254(
.A(net1152),
.ZN(net2380)
);

INV_X16 c2255(
.A(net2357),
.ZN(net2381)
);

INV_X32 c2256(
.A(net2381),
.ZN(net2382)
);

XOR2_X2 c2257(
.A(net464),
.B(net1464),
.Z(net2383)
);

AND3_X4 c2258(
.A1(net1460),
.A2(net449),
.A3(net1374),
.ZN(net2384)
);

INV_X4 c2259(
.A(net9741),
.ZN(net2385)
);

INV_X1 c2260(
.A(net2375),
.ZN(net2386)
);

INV_X2 c2261(
.A(net9741),
.ZN(net2387)
);

INV_X8 c2262(
.A(net2316),
.ZN(net2388)
);

XNOR2_X1 c2263(
.A(net2236),
.B(net2380),
.ZN(net2389)
);

OR2_X4 c2264(
.A1(net2369),
.A2(net2373),
.ZN(net2390)
);

OR2_X1 c2265(
.A1(net2252),
.A2(net425),
.ZN(net2391)
);

XNOR2_X2 c2266(
.A(net2374),
.B(net2383),
.ZN(net2392)
);

DFFS_X1 c2267(
.D(net2386),
.SN(net2260),
.CK(clk),
.Q(net2394),
.QN(net2393)
);

AND2_X4 c2268(
.A1(net2391),
.A2(net2280),
.ZN(net2395)
);

INV_X16 c2269(
.A(net1467),
.ZN(net2396)
);

NAND3_X2 c2270(
.A1(net449),
.A2(net1443),
.A3(net2345),
.ZN(net2397)
);

AND2_X1 c2271(
.A1(net2377),
.A2(net2382),
.ZN(net2398)
);

NAND2_X1 c2272(
.A1(net1444),
.A2(net2257),
.ZN(net2399)
);

NAND2_X2 c2273(
.A1(net2398),
.A2(net2288),
.ZN(net2400)
);

NAND2_X4 c2274(
.A1(net1379),
.A2(net10663),
.ZN(net2401)
);

AND2_X2 c2275(
.A1(net2387),
.A2(net2390),
.ZN(net2402)
);

XOR2_X1 c2276(
.A(net2402),
.B(net2390),
.Z(net2403)
);

NOR2_X1 c2277(
.A1(net2400),
.A2(net2341),
.ZN(net2404)
);

OR2_X2 c2278(
.A1(net2288),
.A2(net1227),
.ZN(net2405)
);

NOR2_X4 c2279(
.A1(net1379),
.A2(net1434),
.ZN(net2406)
);

NOR2_X2 c2280(
.A1(net1343),
.A2(net2400),
.ZN(net2407)
);

DFFRS_X2 c2281(
.D(net2404),
.RN(net2376),
.SN(net1225),
.CK(clk),
.Q(net2409),
.QN(net2408)
);

INV_X32 c2282(
.A(net432),
.ZN(net2410)
);

INV_X4 c2283(
.A(net11410),
.ZN(net2411)
);

XOR2_X2 c2284(
.A(net2394),
.B(net2383),
.Z(net2412)
);

XNOR2_X1 c2285(
.A(net2157),
.B(net2353),
.ZN(net2413)
);

OR2_X4 c2286(
.A1(net2406),
.A2(net1464),
.ZN(net2414)
);

OR3_X1 c2287(
.A1(net1446),
.A2(net2393),
.A3(net2411),
.ZN(net2415)
);

OR2_X1 c2288(
.A1(net2376),
.A2(net2415),
.ZN(net2416)
);

XNOR2_X2 c2289(
.A(net2416),
.B(net2390),
.ZN(net2417)
);

AND2_X4 c2290(
.A1(net1394),
.A2(net1343),
.ZN(net2418)
);

OAI221_X4 c2291(
.A(net2403),
.B1(net449),
.B2(net2241),
.C1(net2390),
.C2(net11322),
.ZN(net2419)
);

AND2_X1 c2292(
.A1(net2370),
.A2(net2336),
.ZN(net2420)
);

NAND2_X1 c2293(
.A1(net2410),
.A2(net10662),
.ZN(net2421)
);

NAND2_X2 c2294(
.A1(net2396),
.A2(net1297),
.ZN(net2422)
);

DFFS_X2 c2295(
.D(net2413),
.SN(net2367),
.CK(clk),
.Q(net2424),
.QN(net2423)
);

INV_X1 c2296(
.A(net2422),
.ZN(net2425)
);

NAND2_X4 c2297(
.A1(net1086),
.A2(net2392),
.ZN(net2426)
);

INV_X2 c2298(
.A(net11482),
.ZN(net2427)
);

INV_X8 c2299(
.A(net11115),
.ZN(net2428)
);

AND2_X2 c2300(
.A1(net2426),
.A2(net2411),
.ZN(net2429)
);

XOR2_X1 c2301(
.A(net2392),
.B(net432),
.Z(net2430)
);

SDFF_X1 c2302(
.D(net1430),
.SE(net428),
.SI(net2348),
.CK(clk),
.Q(net2432),
.QN(net2431)
);

INV_X16 c2303(
.A(net2424),
.ZN(net2433)
);

MUX2_X1 c2304(
.A(net2430),
.B(net2423),
.S(net2403),
.Z(net2434)
);

NOR2_X1 c2305(
.A1(net2407),
.A2(net2374),
.ZN(net2435)
);

OR2_X2 c2306(
.A1(net1411),
.A2(net2427),
.ZN(net2436)
);

NOR2_X4 c2307(
.A1(net2418),
.A2(net2412),
.ZN(net2437)
);

NOR2_X2 c2308(
.A1(net2373),
.A2(net2392),
.ZN(net2438)
);

SDFF_X2 c2309(
.D(net2378),
.SE(net2437),
.SI(net2438),
.CK(clk),
.Q(net2440),
.QN(net2439)
);

INV_X32 c2310(
.A(net10483),
.ZN(net2441)
);

XOR2_X2 c2311(
.A(net2385),
.B(net2432),
.Z(net2442)
);

NAND4_X2 c2312(
.A1(net2432),
.A2(net1431),
.A3(net2439),
.A4(net2438),
.ZN(net2443)
);

OAI222_X4 c2313(
.A1(net2257),
.A2(net2408),
.B1(net2442),
.B2(net2351),
.C1(net2437),
.C2(net2367),
.ZN(net2444)
);

XNOR2_X1 c2314(
.A(net1431),
.B(net2425),
.ZN(net2445)
);

SDFFR_X2 c2315(
.D(net2443),
.RN(net2353),
.SE(net2437),
.SI(net10874),
.CK(clk),
.Q(net2447),
.QN(net2446)
);

OAI21_X4 c2316(
.A(net2429),
.B1(net2435),
.B2(net2439),
.ZN(net2448)
);

OAI222_X2 c2317(
.A1(net2428),
.A2(net2440),
.B1(net2448),
.B2(net2431),
.C1(net2437),
.C2(net1086),
.ZN(net2449)
);

OAI221_X2 c2318(
.A(net2437),
.B1(net2432),
.B2(net2436),
.C1(net2390),
.C2(net2438),
.ZN(net2450)
);

MUX2_X2 c2319(
.A(net1443),
.B(net2437),
.S(net1309),
.Z(net2451)
);

OR4_X4 c2320(
.A1(net2448),
.A2(net2427),
.A3(net2437),
.A4(net11516),
.ZN(net2452)
);

AOI221_X4 c2321(
.A(net2341),
.B1(net2443),
.B2(net2448),
.C1(net2437),
.C2(net2235),
.ZN(net2453)
);

AOI222_X1 c2322(
.A1(net2349),
.A2(net2438),
.B1(net2448),
.B2(net2431),
.C1(net2446),
.C2(net10857),
.ZN(net2454)
);

DFFRS_X1 c2323(
.D(net2441),
.RN(net2448),
.SN(net10727),
.CK(clk),
.Q(net2456),
.QN(net2455)
);

INV_X4 c2324(
.A(net1508),
.ZN(net2457)
);

INV_X1 c2325(
.A(net11407),
.ZN(net2458)
);

OR2_X4 c2326(
.A1(net2451),
.A2(net2421),
.ZN(net2459)
);

INV_X2 c2327(
.A(net535),
.ZN(net2460)
);

INV_X8 c2328(
.A(net2458),
.ZN(net2461)
);

AOI222_X4 c2329(
.A1(net2368),
.A2(net1399),
.B1(net1526),
.B2(net1428),
.C1(net1513),
.C2(net11074),
.ZN(net2462)
);

NAND3_X4 c2330(
.A1(net2353),
.A2(net2363),
.A3(net1374),
.ZN(net2463)
);

INV_X16 c2331(
.A(net11369),
.ZN(net2464)
);

INV_X32 c2332(
.A(net10590),
.ZN(net2465)
);

INV_X4 c2333(
.A(net2442),
.ZN(net2466)
);

OR2_X1 c2334(
.A1(net1530),
.A2(net11308),
.ZN(net2467)
);

XNOR2_X2 c2335(
.A(net2465),
.B(net2451),
.ZN(net2468)
);

INV_X1 c2336(
.A(net10590),
.ZN(net2469)
);

AND2_X4 c2337(
.A1(net1500),
.A2(net2462),
.ZN(net2470)
);

AND2_X1 c2338(
.A1(net2467),
.A2(net496),
.ZN(net2471)
);

NAND2_X1 c2339(
.A1(net1212),
.A2(net1479),
.ZN(net2472)
);

INV_X2 c2340(
.A(net2401),
.ZN(net2473)
);

INV_X8 c2341(
.A(net2469),
.ZN(net2474)
);

NAND2_X2 c2342(
.A1(net2473),
.A2(net2142),
.ZN(net2475)
);

NAND2_X4 c2343(
.A1(net2345),
.A2(net11514),
.ZN(net2476)
);

INV_X16 c2344(
.A(net2475),
.ZN(net2477)
);

AND2_X2 c2345(
.A1(net2427),
.A2(net2471),
.ZN(net2478)
);

INV_X32 c2346(
.A(net10471),
.ZN(net2479)
);

XOR2_X1 c2347(
.A(net2421),
.B(net2415),
.Z(net2480)
);

DFFR_X1 c2348(
.D(net2459),
.RN(net1525),
.CK(clk),
.Q(net2482),
.QN(net2481)
);

NOR2_X1 c2349(
.A1(net2464),
.A2(net2481),
.ZN(net2483)
);

DFFR_X2 c2350(
.D(net1557),
.RN(net2470),
.CK(clk),
.Q(net2485),
.QN(net2484)
);

OR2_X2 c2351(
.A1(net2460),
.A2(net2464),
.ZN(net2486)
);

NOR2_X4 c2352(
.A1(net2486),
.A2(net2476),
.ZN(net2487)
);

OR3_X4 c2353(
.A1(net2482),
.A2(net2312),
.A3(net1526),
.ZN(net2488)
);

INV_X4 c2354(
.A(net1519),
.ZN(net2489)
);

NOR2_X2 c2355(
.A1(net2466),
.A2(net2486),
.ZN(net2490)
);

INV_X1 c2356(
.A(net2476),
.ZN(net2491)
);

INV_X2 c2357(
.A(net1532),
.ZN(net2492)
);

DFFRS_X2 c2358(
.D(net1552),
.RN(net2475),
.SN(net1418),
.CK(clk),
.Q(net2494),
.QN(net2493)
);

AOI221_X2 c2359(
.A(net2359),
.B1(net2466),
.B2(net2487),
.C1(net2476),
.C2(net1513),
.ZN(net2495)
);

INV_X8 c2360(
.A(net11193),
.ZN(net2496)
);

XOR2_X2 c2361(
.A(net2462),
.B(net2479),
.Z(net2497)
);

DFFS_X1 c2362(
.D(net2479),
.SN(net2371),
.CK(clk),
.Q(net2499),
.QN(net2498)
);

XNOR2_X1 c2363(
.A(net2415),
.B(net2451),
.ZN(net2500)
);

OR2_X4 c2364(
.A1(net2472),
.A2(net2493),
.ZN(net2501)
);

INV_X16 c2365(
.A(net10589),
.ZN(net2502)
);

OR2_X1 c2366(
.A1(net2323),
.A2(net2457),
.ZN(net2503)
);

INV_X32 c2367(
.A(net2414),
.ZN(net2504)
);

XNOR2_X2 c2368(
.A(net2362),
.B(net11357),
.ZN(net2505)
);

AND2_X4 c2369(
.A1(net2483),
.A2(net11507),
.ZN(net2506)
);

AND3_X2 c2370(
.A1(net1468),
.A2(net2482),
.A3(net2368),
.ZN(net2507)
);

AND2_X1 c2371(
.A1(net2479),
.A2(net346),
.ZN(net2508)
);

NAND2_X1 c2372(
.A1(net2495),
.A2(net2415),
.ZN(net2509)
);

INV_X4 c2373(
.A(net2499),
.ZN(net2510)
);

NAND2_X2 c2374(
.A1(net1489),
.A2(net2500),
.ZN(net2511)
);

NAND2_X4 c2375(
.A1(net2405),
.A2(net2485),
.ZN(net2512)
);

INV_X1 c2376(
.A(net1541),
.ZN(net2513)
);

AND2_X2 c2377(
.A1(net524),
.A2(net11506),
.ZN(net2514)
);

XOR2_X1 c2378(
.A(net1470),
.B(net2379),
.Z(net2515)
);

INV_X2 c2379(
.A(net2507),
.ZN(net2516)
);

NOR2_X1 c2380(
.A1(net1548),
.A2(net2476),
.ZN(net2517)
);

INV_X8 c2381(
.A(net10131),
.ZN(net2518)
);

OR2_X2 c2382(
.A1(net2502),
.A2(net2499),
.ZN(net2519)
);

OAI33_X1 c2383(
.A1(net2492),
.A2(net2488),
.A3(net2405),
.B1(net2479),
.B2(net1399),
.B3(net2483),
.ZN(net2520)
);

NOR3_X1 c2384(
.A1(net522),
.A2(net2477),
.A3(net1513),
.ZN(net2521)
);

NOR2_X4 c2385(
.A1(net2515),
.A2(net2514),
.ZN(net2522)
);

INV_X16 c2386(
.A(net11054),
.ZN(net2523)
);

OR3_X2 c2387(
.A1(net2504),
.A2(net2473),
.A3(net2490),
.ZN(net2524)
);

NOR2_X2 c2388(
.A1(net2518),
.A2(net2483),
.ZN(net2525)
);

XOR2_X2 c2389(
.A(net2525),
.B(net2481),
.Z(net2526)
);

SDFF_X1 c2390(
.D(net2524),
.SE(net2501),
.SI(net1541),
.CK(clk),
.Q(net2528),
.QN(net2527)
);

OAI21_X2 c2391(
.A(net2464),
.B1(net2479),
.B2(net2526),
.ZN(net2529)
);

XNOR2_X1 c2392(
.A(net2475),
.B(net2526),
.ZN(net2530)
);

OR2_X4 c2393(
.A1(net2516),
.A2(net2523),
.ZN(net2531)
);

OR2_X1 c2394(
.A1(net2487),
.A2(net466),
.ZN(net2532)
);

XNOR2_X2 c2395(
.A(net2488),
.B(net2530),
.ZN(net2533)
);

SDFFRS_X1 c2396(
.D(net2480),
.RN(net2528),
.SE(net2529),
.SI(net1541),
.SN(net2461),
.CK(clk),
.Q(net2535),
.QN(net2534)
);

AND2_X4 c2397(
.A1(net2478),
.A2(net2533),
.ZN(net2536)
);

AOI222_X2 c2398(
.A1(net2512),
.A2(net2498),
.B1(net2526),
.B2(net1513),
.C1(net1374),
.C2(net11517),
.ZN(net2537)
);

INV_X32 c2399(
.A(net11369),
.ZN(net2538)
);

AND2_X1 c2400(
.A1(net2538),
.A2(net2479),
.ZN(net2539)
);

OAI21_X1 c2401(
.A(net2531),
.B1(net2304),
.B2(net2461),
.ZN(net2540)
);

AOI21_X2 c2402(
.A(net2539),
.B1(net2494),
.B2(net2500),
.ZN(net2541)
);

INV_X4 c2403(
.A(net11017),
.ZN(net2542)
);

INV_X1 c2404(
.A(net10371),
.ZN(net2543)
);

SDFF_X2 c2405(
.D(net2543),
.SE(net2522),
.SI(net2540),
.CK(clk),
.Q(net2545),
.QN(net2544)
);

AOI221_X1 c2406(
.A(net2500),
.B1(net2521),
.B2(net1513),
.C1(net2544),
.C2(net2527),
.ZN(net2546)
);

INV_X2 c2407(
.A(net10075),
.ZN(net2547)
);

INV_X8 c2408(
.A(net1644),
.ZN(net2548)
);

NAND2_X1 c2409(
.A1(net1504),
.A2(net2530),
.ZN(net2549)
);

INV_X16 c2410(
.A(net9713),
.ZN(net2550)
);

INV_X32 c2411(
.A(net1447),
.ZN(net2551)
);

INV_X4 c2412(
.A(net2549),
.ZN(net2552)
);

INV_X1 c2413(
.A(net9854),
.ZN(net2553)
);

AOI21_X1 c2414(
.A(net2142),
.B1(net2553),
.B2(net1513),
.ZN(net2554)
);

INV_X2 c2415(
.A(net10228),
.ZN(net2555)
);

INV_X8 c2416(
.A(net1631),
.ZN(net2556)
);

AOI21_X4 c2417(
.A(net2547),
.B1(net2555),
.B2(net10873),
.ZN(net2557)
);

INV_X16 c2418(
.A(net596),
.ZN(net2558)
);

INV_X32 c2419(
.A(net1580),
.ZN(net2559)
);

NAND2_X2 c2420(
.A1(net2557),
.A2(net1619),
.ZN(net2560)
);

NAND2_X4 c2421(
.A1(net1584),
.A2(net2554),
.ZN(net2561)
);

AND2_X2 c2422(
.A1(net2503),
.A2(net11515),
.ZN(net2562)
);

XOR2_X1 c2423(
.A(net2304),
.B(net2557),
.Z(net2563)
);

INV_X4 c2424(
.A(net9848),
.ZN(net2564)
);

INV_X1 c2425(
.A(net2558),
.ZN(net2565)
);

OAI22_X2 c2426(
.A1(net2548),
.A2(net1607),
.B1(net1632),
.B2(net2461),
.ZN(net2566)
);

NOR2_X1 c2427(
.A1(net2565),
.A2(net2555),
.ZN(net2567)
);

OR2_X2 c2428(
.A1(net2559),
.A2(net1646),
.ZN(net2568)
);

NOR2_X4 c2429(
.A1(net2529),
.A2(net2510),
.ZN(net2569)
);

NOR2_X2 c2430(
.A1(net605),
.A2(net2471),
.ZN(net2570)
);

INV_X2 c2431(
.A(net656),
.ZN(net2571)
);

INV_X8 c2432(
.A(net10272),
.ZN(net2572)
);

AND3_X1 c2433(
.A1(net2483),
.A2(net2563),
.A3(net2457),
.ZN(net2573)
);

INV_X16 c2434(
.A(net11420),
.ZN(net2574)
);

XOR2_X2 c2435(
.A(net2471),
.B(net2570),
.Z(net2575)
);

DFFRS_X1 c2436(
.D(net2563),
.RN(net2566),
.SN(net2567),
.CK(clk),
.Q(net2577),
.QN(net2576)
);

XNOR2_X1 c2437(
.A(net616),
.B(net2553),
.ZN(net2578)
);

OR2_X4 c2438(
.A1(net2572),
.A2(net1594),
.ZN(net2579)
);

INV_X32 c2439(
.A(net10278),
.ZN(net2580)
);

OR2_X1 c2440(
.A1(net2562),
.A2(net2577),
.ZN(net2581)
);

XNOR2_X2 c2441(
.A(net2578),
.B(net2457),
.ZN(net2582)
);

NAND3_X1 c2442(
.A1(net2579),
.A2(net2565),
.A3(net2581),
.ZN(net2583)
);

AND2_X4 c2443(
.A1(net2474),
.A2(net10525),
.ZN(net2584)
);

AND2_X1 c2444(
.A1(net2574),
.A2(net2304),
.ZN(net2585)
);

INV_X4 c2445(
.A(net9713),
.ZN(net2586)
);

INV_X1 c2446(
.A(net10494),
.ZN(net2587)
);

NOR3_X4 c2447(
.A1(net2553),
.A2(net2547),
.A3(net1604),
.ZN(net2588)
);

INV_X2 c2448(
.A(net10427),
.ZN(net2589)
);

OAI211_X4 c2449(
.A(net1428),
.B(net2587),
.C1(net2581),
.C2(net2380),
.ZN(net2590)
);

NAND2_X1 c2450(
.A1(net2503),
.A2(net1607),
.ZN(net2591)
);

NOR3_X2 c2451(
.A1(net2489),
.A2(net2511),
.A3(net11119),
.ZN(net2592)
);

DFFS_X2 c2452(
.D(net2501),
.SN(net11018),
.CK(clk),
.Q(net2594),
.QN(net2593)
);

NAND2_X2 c2453(
.A1(net2571),
.A2(net466),
.ZN(net2595)
);

NAND2_X4 c2454(
.A1(net2577),
.A2(net2529),
.ZN(net2596)
);

AND2_X2 c2455(
.A1(net2587),
.A2(net2508),
.ZN(net2597)
);

XOR2_X1 c2456(
.A(net2581),
.B(net1647),
.Z(net2598)
);

NOR2_X1 c2457(
.A1(net2596),
.A2(net2553),
.ZN(net2599)
);

INV_X8 c2458(
.A(net2468),
.ZN(net2600)
);

AND3_X4 c2459(
.A1(net2591),
.A2(net2580),
.A3(net2555),
.ZN(net2601)
);

NAND3_X2 c2460(
.A1(net2564),
.A2(net2581),
.A3(net1609),
.ZN(net2602)
);

OR2_X2 c2461(
.A1(net1633),
.A2(net1646),
.ZN(net2603)
);

NOR2_X4 c2462(
.A1(net2436),
.A2(net1644),
.ZN(net2604)
);

NOR2_X2 c2463(
.A1(net1632),
.A2(net1428),
.ZN(net2605)
);

INV_X16 c2464(
.A(net2604),
.ZN(net2606)
);

XOR2_X2 c2465(
.A(net1618),
.B(net11086),
.Z(net2607)
);

XNOR2_X1 c2466(
.A(net2599),
.B(net1635),
.ZN(net2608)
);

INV_X32 c2467(
.A(net2584),
.ZN(net2609)
);

OR2_X4 c2468(
.A1(net2547),
.A2(net2581),
.ZN(net2610)
);

INV_X4 c2469(
.A(net10524),
.ZN(net2611)
);

OR2_X1 c2470(
.A1(net2611),
.A2(net638),
.ZN(net2612)
);

XNOR2_X2 c2471(
.A(net2457),
.B(net1580),
.ZN(net2613)
);

AND2_X4 c2472(
.A1(net2612),
.A2(net2610),
.ZN(net2614)
);

AND2_X1 c2473(
.A1(net357),
.A2(net2380),
.ZN(net2615)
);

NAND2_X1 c2474(
.A1(net2510),
.A2(net2576),
.ZN(net2616)
);

NAND2_X2 c2475(
.A1(net2607),
.A2(net2604),
.ZN(net2617)
);

NAND2_X4 c2476(
.A1(net1618),
.A2(net2580),
.ZN(net2618)
);

AND2_X2 c2477(
.A1(net2616),
.A2(net2604),
.ZN(net2619)
);

SDFFS_X1 c2478(
.D(net652),
.SE(net2619),
.SI(net2529),
.SN(net1635),
.CK(clk),
.Q(net2621),
.QN(net2620)
);

OAI211_X1 c2479(
.A(net2613),
.B(net1643),
.C1(net1635),
.C2(net11517),
.ZN(net2622)
);

XOR2_X1 c2480(
.A(net2595),
.B(net2608),
.Z(net2623)
);

INV_X1 c2481(
.A(net9940),
.ZN(net2624)
);

OR3_X1 c2482(
.A1(net2555),
.A2(net2616),
.A3(net2571),
.ZN(net2625)
);

NOR4_X4 c2483(
.A1(net2622),
.A2(net2620),
.A3(net2625),
.A4(net2593),
.ZN(net2626)
);

NOR2_X1 c2484(
.A1(net2598),
.A2(net2608),
.ZN(net2627)
);

NOR4_X2 c2485(
.A1(net2624),
.A2(net2610),
.A3(net2503),
.A4(net656),
.ZN(net2628)
);

MUX2_X1 c2486(
.A(net2234),
.B(net2572),
.S(net2557),
.Z(net2629)
);

AOI211_X4 c2487(
.A(net2624),
.B(net2618),
.C1(net2629),
.C2(net10807),
.ZN(net2630)
);

OAI21_X4 c2488(
.A(net2615),
.B1(net2623),
.B2(net11086),
.ZN(net2631)
);

MUX2_X2 c2489(
.A(net2628),
.B(net2609),
.S(net11005),
.Z(net2632)
);

DFFR_X1 c2490(
.D(net752),
.RN(net2546),
.CK(clk),
.Q(net2634),
.QN(net2633)
);

OR2_X2 c2491(
.A1(net1651),
.A2(net1642),
.ZN(net2635)
);

NOR2_X4 c2492(
.A1(net2560),
.A2(net2554),
.ZN(net2636)
);

INV_X2 c2493(
.A(net2462),
.ZN(net2637)
);

INV_X8 c2494(
.A(net1693),
.ZN(net2638)
);

NOR2_X2 c2495(
.A1(net2608),
.A2(net2556),
.ZN(net2639)
);

XOR2_X2 c2496(
.A(net2496),
.B(net2519),
.Z(net2640)
);

INV_X16 c2497(
.A(net9797),
.ZN(net2641)
);

NAND3_X4 c2498(
.A1(net2639),
.A2(net1599),
.A3(net707),
.ZN(net2642)
);

XNOR2_X1 c2499(
.A(net2640),
.B(net1693),
.ZN(net2643)
);

OR2_X4 c2500(
.A1(net1644),
.A2(net2643),
.ZN(net2644)
);

OR2_X1 c2501(
.A1(net2550),
.A2(net2637),
.ZN(net2645)
);

INV_X32 c2502(
.A(net11393),
.ZN(net2646)
);

XNOR2_X2 c2503(
.A(net2644),
.B(net2312),
.ZN(net2647)
);

INV_X4 c2504(
.A(net1373),
.ZN(net2648)
);

INV_X1 c2505(
.A(net1666),
.ZN(net2649)
);

AND2_X4 c2506(
.A1(net1642),
.A2(net707),
.ZN(net2650)
);

AND2_X1 c2507(
.A1(net2312),
.A2(net2608),
.ZN(net2651)
);

NAND2_X1 c2508(
.A1(net1702),
.A2(net1730),
.ZN(net2652)
);

OR3_X4 c2509(
.A1(net1523),
.A2(net1635),
.A3(net2477),
.ZN(net2653)
);

INV_X2 c2510(
.A(net10178),
.ZN(net2654)
);

NAND2_X2 c2511(
.A1(net2625),
.A2(net11120),
.ZN(net2655)
);

NAND2_X4 c2512(
.A1(net2568),
.A2(net2550),
.ZN(net2656)
);

AND2_X2 c2513(
.A1(net686),
.A2(net2625),
.ZN(net2657)
);

XOR2_X1 c2514(
.A(net1685),
.B(net2483),
.Z(net2658)
);

NOR2_X1 c2515(
.A1(net2474),
.A2(net2570),
.ZN(net2659)
);

INV_X8 c2516(
.A(net11151),
.ZN(net2660)
);

INV_X16 c2517(
.A(net11367),
.ZN(net2661)
);

OR2_X2 c2518(
.A1(net1695),
.A2(net2649),
.ZN(net2662)
);

NOR2_X4 c2519(
.A1(net1692),
.A2(net1718),
.ZN(net2663)
);

INV_X32 c2520(
.A(net10226),
.ZN(net2664)
);

AND3_X2 c2521(
.A1(net2556),
.A2(net2638),
.A3(net2647),
.ZN(net2665)
);

NOR2_X2 c2522(
.A1(net2654),
.A2(net1696),
.ZN(net2666)
);

XOR2_X2 c2523(
.A(net2656),
.B(net2568),
.Z(net2667)
);

INV_X4 c2524(
.A(net9797),
.ZN(net2668)
);

INV_X1 c2525(
.A(net9971),
.ZN(net2669)
);

INV_X2 c2526(
.A(net2505),
.ZN(net2670)
);

XNOR2_X1 c2527(
.A(net1732),
.B(net2666),
.ZN(net2671)
);

NOR4_X1 c2528(
.A1(net2648),
.A2(net1692),
.A3(net2669),
.A4(net2649),
.ZN(net2672)
);

INV_X8 c2529(
.A(net1689),
.ZN(net2673)
);

OR2_X4 c2530(
.A1(net2673),
.A2(net1734),
.ZN(net2674)
);

OR2_X1 c2531(
.A1(net2666),
.A2(net10584),
.ZN(net2675)
);

INV_X16 c2532(
.A(net10399),
.ZN(net2676)
);

XNOR2_X2 c2533(
.A(net2675),
.B(net2461),
.ZN(net2677)
);

OAI221_X1 c2534(
.A(net2477),
.B1(net2670),
.B2(net2660),
.C1(net1731),
.C2(net1399),
.ZN(net2678)
);

AND2_X4 c2535(
.A1(net1619),
.A2(net2554),
.ZN(net2679)
);

NOR3_X1 c2536(
.A1(net2636),
.A2(net2653),
.A3(net686),
.ZN(net2680)
);

AND2_X1 c2537(
.A1(net705),
.A2(net2640),
.ZN(net2681)
);

NAND2_X1 c2538(
.A1(net2677),
.A2(net2670),
.ZN(net2682)
);

NAND2_X2 c2539(
.A1(net2519),
.A2(net2670),
.ZN(net2683)
);

NAND2_X4 c2540(
.A1(net2664),
.A2(net2658),
.ZN(net2684)
);

DFFR_X2 c2541(
.D(net2660),
.RN(net1703),
.CK(clk),
.Q(net2686),
.QN(net2685)
);

OR3_X2 c2542(
.A1(net2570),
.A2(net1689),
.A3(net2685),
.ZN(net2687)
);

DFFS_X1 c2543(
.D(net2647),
.SN(net705),
.CK(clk),
.Q(net2689),
.QN(net2688)
);

AND2_X2 c2544(
.A1(net2409),
.A2(net2679),
.ZN(net2690)
);

XOR2_X1 c2545(
.A(net1660),
.B(net2686),
.Z(net2691)
);

INV_X32 c2546(
.A(net11134),
.ZN(net2692)
);

NOR2_X1 c2547(
.A1(net2554),
.A2(net2686),
.ZN(net2693)
);

OAI21_X2 c2548(
.A(net2693),
.B1(net2664),
.B2(net2679),
.ZN(net2694)
);

OR2_X2 c2549(
.A1(net1662),
.A2(net2644),
.ZN(net2695)
);

INV_X4 c2550(
.A(net11255),
.ZN(net2696)
);

NOR2_X4 c2551(
.A1(net2659),
.A2(net2687),
.ZN(net2697)
);

NOR2_X2 c2552(
.A1(net991),
.A2(net2685),
.ZN(net2698)
);

XOR2_X2 c2553(
.A(net1706),
.B(net2679),
.Z(net2699)
);

XNOR2_X1 c2554(
.A(net1712),
.B(net2671),
.ZN(net2700)
);

OR2_X4 c2555(
.A1(net2689),
.A2(net11149),
.ZN(net2701)
);

OR2_X1 c2556(
.A1(net2646),
.A2(net1701),
.ZN(net2702)
);

DFFRS_X2 c2557(
.D(net2672),
.RN(net2654),
.SN(net11359),
.CK(clk),
.Q(net2704),
.QN(net2703)
);

INV_X1 c2558(
.A(net10415),
.ZN(net2705)
);

XNOR2_X2 c2559(
.A(net2668),
.B(net2691),
.ZN(net2706)
);

OAI221_X4 c2560(
.A(net2705),
.B1(net2706),
.B2(net2483),
.C1(net699),
.C2(net2670),
.ZN(net2707)
);

INV_X2 c2561(
.A(net10225),
.ZN(net2708)
);

OAI21_X1 c2562(
.A(net2708),
.B1(net626),
.B2(net11212),
.ZN(net2709)
);

AND2_X4 c2563(
.A1(net2697),
.A2(net2696),
.ZN(net2710)
);

AOI21_X2 c2564(
.A(net2710),
.B1(net2709),
.B2(net2692),
.ZN(net2711)
);

OAI222_X1 c2565(
.A1(net2658),
.A2(net2706),
.B1(net758),
.B2(net1599),
.C1(net2697),
.C2(net2709),
.ZN(net2712)
);

AOI21_X1 c2566(
.A(net2575),
.B1(net2703),
.B2(net11212),
.ZN(net2713)
);

AOI21_X4 c2567(
.A(net2682),
.B1(net2712),
.B2(net11470),
.ZN(net2714)
);

AND2_X1 c2568(
.A1(net2686),
.A2(net2654),
.ZN(net2715)
);

AND3_X1 c2569(
.A1(net2708),
.A2(net2709),
.A3(net1729),
.ZN(net2716)
);

OAI221_X2 c2570(
.A(net2709),
.B1(net2692),
.B2(net2649),
.C1(net10853),
.C2(net11470),
.ZN(net2717)
);

NAND2_X1 c2571(
.A1(net2712),
.A2(net2683),
.ZN(net2718)
);

INV_X8 c2572(
.A(net10466),
.ZN(net2719)
);

INV_X16 c2573(
.A(net11340),
.ZN(net2720)
);

NAND2_X2 c2574(
.A1(net1800),
.A2(net2638),
.ZN(net2721)
);

INV_X32 c2575(
.A(net11452),
.ZN(net2722)
);

INV_X4 c2576(
.A(net812),
.ZN(net2723)
);

INV_X1 c2577(
.A(net2678),
.ZN(net2724)
);

INV_X2 c2578(
.A(net2652),
.ZN(net2725)
);

AOI211_X2 c2579(
.A(net1801),
.B(net1810),
.C1(net2580),
.C2(net2692),
.ZN(net2726)
);

NAND2_X4 c2580(
.A1(net1820),
.A2(net2671),
.ZN(net2727)
);

AND2_X2 c2581(
.A1(net2707),
.A2(net1800),
.ZN(net2728)
);

INV_X8 c2582(
.A(net1809),
.ZN(net2729)
);

NAND3_X1 c2583(
.A1(net2721),
.A2(net1701),
.A3(net1810),
.ZN(net2730)
);

INV_X16 c2584(
.A(net10458),
.ZN(net2731)
);

INV_X32 c2585(
.A(net9745),
.ZN(net2732)
);

INV_X4 c2586(
.A(net2641),
.ZN(net2733)
);

INV_X1 c2587(
.A(net10329),
.ZN(net2734)
);

XOR2_X1 c2588(
.A(net1499),
.B(net2534),
.Z(net2735)
);

NOR2_X1 c2589(
.A1(net2692),
.A2(net1752),
.ZN(net2736)
);

INV_X2 c2590(
.A(net2727),
.ZN(net2737)
);

INV_X8 c2591(
.A(net2691),
.ZN(net2738)
);

INV_X16 c2592(
.A(net2701),
.ZN(net2739)
);

NOR3_X4 c2593(
.A1(net2723),
.A2(net2725),
.A3(net2739),
.ZN(net2740)
);

INV_X32 c2594(
.A(net2638),
.ZN(net2741)
);

INV_X4 c2595(
.A(net11380),
.ZN(net2742)
);

OR2_X2 c2596(
.A1(net2579),
.A2(net1760),
.ZN(net2743)
);

NOR2_X4 c2597(
.A1(net2742),
.A2(net2692),
.ZN(net2744)
);

INV_X1 c2598(
.A(net11318),
.ZN(net2745)
);

INV_X2 c2599(
.A(net10585),
.ZN(net2746)
);

NOR2_X2 c2600(
.A1(net2736),
.A2(net1800),
.ZN(net2747)
);

NOR3_X2 c2601(
.A1(net2546),
.A2(net2688),
.A3(net2724),
.ZN(net2748)
);

XOR2_X2 c2602(
.A(net2731),
.B(net1595),
.Z(net2749)
);

XNOR2_X1 c2603(
.A(net1737),
.B(net810),
.ZN(net2750)
);

OR2_X4 c2604(
.A1(net834),
.A2(net2579),
.ZN(net2751)
);

OR2_X1 c2605(
.A1(net1803),
.A2(net2751),
.ZN(net2752)
);

INV_X8 c2606(
.A(net1792),
.ZN(net2753)
);

XNOR2_X2 c2607(
.A(net2746),
.B(net1776),
.ZN(net2754)
);

AND2_X4 c2608(
.A1(net1752),
.A2(net2709),
.ZN(net2755)
);

AND2_X1 c2609(
.A1(net2721),
.A2(net11349),
.ZN(net2756)
);

NAND2_X1 c2610(
.A1(net2715),
.A2(net1686),
.ZN(net2757)
);

INV_X16 c2611(
.A(net9745),
.ZN(net2758)
);

NAND2_X2 c2612(
.A1(net2757),
.A2(net699),
.ZN(net2759)
);

INV_X32 c2613(
.A(net11051),
.ZN(net2760)
);

NAND2_X4 c2614(
.A1(net2745),
.A2(net2580),
.ZN(net2761)
);

AND2_X2 c2615(
.A1(net2637),
.A2(net1737),
.ZN(net2762)
);

XOR2_X1 c2616(
.A(net2758),
.B(net11355),
.Z(net2763)
);

DFFS_X2 c2617(
.D(net1818),
.SN(net2758),
.CK(clk),
.Q(net2765),
.QN(net2764)
);

NOR2_X1 c2618(
.A1(net2722),
.A2(net2758),
.ZN(net2766)
);

OR2_X2 c2619(
.A1(net2666),
.A2(net2766),
.ZN(net2767)
);

NOR2_X4 c2620(
.A1(net1815),
.A2(net626),
.ZN(net2768)
);

NOR2_X2 c2621(
.A1(net2737),
.A2(net2752),
.ZN(net2769)
);

XOR2_X2 c2622(
.A(net2752),
.B(net2671),
.Z(net2770)
);

AOI22_X1 c2623(
.A1(net2738),
.A2(net2751),
.B1(net2763),
.B2(net2753),
.ZN(net2771)
);

XNOR2_X1 c2624(
.A(net2770),
.B(net2769),
.ZN(net2772)
);

OR2_X4 c2625(
.A1(net2655),
.A2(net1809),
.ZN(net2773)
);

AOI221_X4 c2626(
.A(net2768),
.B1(net2728),
.B2(net1800),
.C1(net1743),
.C2(net2749),
.ZN(net2774)
);

AND3_X4 c2627(
.A1(net2728),
.A2(net2758),
.A3(net11189),
.ZN(net2775)
);

OR2_X1 c2628(
.A1(net2761),
.A2(net2769),
.ZN(net2776)
);

XNOR2_X2 c2629(
.A(net1794),
.B(net2692),
.ZN(net2777)
);

AND2_X4 c2630(
.A1(net2743),
.A2(net2741),
.ZN(net2778)
);

NAND3_X2 c2631(
.A1(net2775),
.A2(net2758),
.A3(net2723),
.ZN(net2779)
);

SDFF_X1 c2632(
.D(net2776),
.SE(net2772),
.SI(net2778),
.CK(clk),
.Q(net2781),
.QN(net2780)
);

AND2_X1 c2633(
.A1(net2740),
.A2(net2739),
.ZN(net2782)
);

NAND2_X1 c2634(
.A1(net2782),
.A2(net2780),
.ZN(net2783)
);

NAND2_X2 c2635(
.A1(net2741),
.A2(net2759),
.ZN(net2784)
);

INV_X4 c2636(
.A(net11052),
.ZN(net2785)
);

NAND2_X4 c2637(
.A1(net2756),
.A2(net11355),
.ZN(net2786)
);

SDFFS_X2 c2638(
.D(net2786),
.SE(net2764),
.SI(net2773),
.SN(net2758),
.CK(clk),
.Q(net2788),
.QN(net2787)
);

OR3_X1 c2639(
.A1(net2783),
.A2(net2508),
.A3(net2579),
.ZN(net2789)
);

AND2_X2 c2640(
.A1(net2363),
.A2(net2787),
.ZN(net2790)
);

AND4_X4 c2641(
.A1(net2698),
.A2(net2671),
.A3(net2787),
.A4(net2754),
.ZN(net2791)
);

XOR2_X1 c2642(
.A(net2756),
.B(net2791),
.Z(net2792)
);

AOI221_X2 c2643(
.A(net707),
.B1(net2594),
.B2(net2753),
.C1(net2749),
.C2(net11349),
.ZN(net2793)
);

NOR2_X1 c2644(
.A1(net2728),
.A2(net2786),
.ZN(net2794)
);

OR2_X2 c2645(
.A1(net2793),
.A2(net1667),
.ZN(net2795)
);

DFFR_X1 c2646(
.D(net2766),
.RN(net2794),
.CK(clk),
.Q(net2797),
.QN(net2796)
);

INV_X1 c2647(
.A(net11350),
.ZN(net2798)
);

NOR2_X4 c2648(
.A1(net2798),
.A2(net2788),
.ZN(net2799)
);

AOI221_X1 c2649(
.A(net2789),
.B1(net2786),
.B2(net2782),
.C1(net2799),
.C2(net2749),
.ZN(net2800)
);

NOR2_X2 c2650(
.A1(net2784),
.A2(net2752),
.ZN(net2801)
);

XOR2_X2 c2651(
.A(net2792),
.B(net2794),
.Z(net2802)
);

XNOR2_X1 c2652(
.A(net2774),
.B(net2796),
.ZN(net2803)
);

OR2_X4 c2653(
.A1(net2759),
.A2(net2797),
.ZN(net2804)
);

OR2_X1 c2654(
.A1(net1562),
.A2(net10946),
.ZN(net2805)
);

XNOR2_X2 c2655(
.A(net2796),
.B(net11356),
.ZN(net2806)
);

AND2_X4 c2656(
.A1(net1901),
.A2(net1860),
.ZN(net2807)
);

AND2_X1 c2657(
.A1(net1762),
.A2(net1838),
.ZN(net2808)
);

NAND2_X1 c2658(
.A1(net1831),
.A2(net2769),
.ZN(net2809)
);

MUX2_X1 c2659(
.A(net2734),
.B(net1887),
.S(net1750),
.Z(net2810)
);

OAI221_X1 c2660(
.A(net1718),
.B1(net939),
.B2(net863),
.C1(net2751),
.C2(net784),
.ZN(net2811)
);

DFFR_X2 c2661(
.D(net2623),
.RN(net10757),
.CK(clk),
.Q(net2813),
.QN(net2812)
);

NAND2_X2 c2662(
.A1(net934),
.A2(net2808),
.ZN(net2814)
);

INV_X2 c2663(
.A(net9756),
.ZN(net2815)
);

NAND2_X4 c2664(
.A1(net1871),
.A2(net2813),
.ZN(net2816)
);

AND2_X2 c2665(
.A1(net2814),
.A2(net1870),
.ZN(net2817)
);

XOR2_X1 c2666(
.A(net1613),
.B(net900),
.Z(net2818)
);

DFFS_X1 c2667(
.D(net779),
.SN(net2623),
.CK(clk),
.Q(net2820),
.QN(net2819)
);

DFFS_X2 c2668(
.D(net2818),
.SN(net1845),
.CK(clk),
.Q(net2822),
.QN(net2821)
);

NOR2_X1 c2669(
.A1(net882),
.A2(net889),
.ZN(net2823)
);

OR2_X2 c2670(
.A1(net2380),
.A2(net900),
.ZN(net2824)
);

NOR2_X4 c2671(
.A1(net939),
.A2(net1857),
.ZN(net2825)
);

NOR2_X2 c2672(
.A1(net2797),
.A2(net1807),
.ZN(net2826)
);

XOR2_X2 c2673(
.A(net933),
.B(net900),
.Z(net2827)
);

XNOR2_X1 c2674(
.A(net800),
.B(net1860),
.ZN(net2828)
);

OAI21_X4 c2675(
.A(net699),
.B1(net2785),
.B2(net914),
.ZN(net2829)
);

OR2_X4 c2676(
.A1(net901),
.A2(net2818),
.ZN(net2830)
);

OR2_X1 c2677(
.A1(net912),
.A2(net2812),
.ZN(net2831)
);

XNOR2_X2 c2678(
.A(net2813),
.B(net2826),
.ZN(net2832)
);

AND2_X4 c2679(
.A1(net1667),
.A2(net2814),
.ZN(net2833)
);

AND2_X1 c2680(
.A1(net2767),
.A2(net934),
.ZN(net2834)
);

NAND2_X1 c2681(
.A1(net1880),
.A2(net2811),
.ZN(net2835)
);

INV_X8 c2682(
.A(net2755),
.ZN(net2836)
);

NAND2_X2 c2683(
.A1(net2653),
.A2(net2811),
.ZN(net2837)
);

INV_X16 c2684(
.A(net10407),
.ZN(net2838)
);

NAND2_X4 c2685(
.A1(net1863),
.A2(net2829),
.ZN(net2839)
);

AND2_X2 c2686(
.A1(net1760),
.A2(net2824),
.ZN(net2840)
);

XOR2_X1 c2687(
.A(net2788),
.B(net2815),
.Z(net2841)
);

NOR2_X1 c2688(
.A1(net877),
.A2(net10537),
.ZN(net2842)
);

SDFF_X2 c2689(
.D(net2825),
.SE(net1868),
.SI(net1871),
.CK(clk),
.Q(net2844),
.QN(net2843)
);

OR2_X2 c2690(
.A1(net932),
.A2(net1807),
.ZN(net2845)
);

MUX2_X2 c2691(
.A(net1844),
.B(net2790),
.S(net1840),
.Z(net2846)
);

NOR2_X4 c2692(
.A1(net1888),
.A2(net2846),
.ZN(net2847)
);

NOR2_X2 c2693(
.A1(net900),
.A2(net2838),
.ZN(net2848)
);

XOR2_X2 c2694(
.A(net2841),
.B(net2839),
.Z(net2849)
);

XNOR2_X1 c2695(
.A(net926),
.B(net2846),
.ZN(net2850)
);

OAI221_X4 c2696(
.A(net2790),
.B1(net1867),
.B2(net1750),
.C1(net2839),
.C2(net2848),
.ZN(net2851)
);

DFFRS_X1 c2697(
.D(net2851),
.RN(net2827),
.SN(net926),
.CK(clk),
.Q(net2853),
.QN(net2852)
);

OR2_X4 c2698(
.A1(net1841),
.A2(net2852),
.ZN(net2854)
);

OR2_X1 c2699(
.A1(net823),
.A2(net1870),
.ZN(net2855)
);

XNOR2_X2 c2700(
.A(net2847),
.B(net882),
.ZN(net2856)
);

NAND3_X4 c2701(
.A1(net2769),
.A2(net2836),
.A3(net1759),
.ZN(net2857)
);

AND2_X4 c2702(
.A1(net909),
.A2(net1762),
.ZN(net2858)
);

SDFFRS_X2 c2703(
.D(net922),
.RN(net2623),
.SE(net2780),
.SI(net2814),
.SN(net1870),
.CK(clk),
.Q(net2860),
.QN(net2859)
);

DFFR_X1 c2704(
.D(net2689),
.RN(net2857),
.CK(clk),
.Q(net2862),
.QN(net2861)
);

OR3_X4 c2705(
.A1(net2834),
.A2(net2862),
.A3(net863),
.ZN(net2863)
);

NAND4_X1 c2706(
.A1(net2858),
.A2(net1893),
.A3(net933),
.A4(net2849),
.ZN(net2864)
);

AND2_X1 c2707(
.A1(net2838),
.A2(net10991),
.ZN(net2865)
);

INV_X32 c2708(
.A(net9919),
.ZN(net2866)
);

INV_X4 c2709(
.A(net10400),
.ZN(net2867)
);

DFFR_X2 c2710(
.D(net2830),
.RN(net2850),
.CK(clk),
.Q(net2869),
.QN(net2868)
);

NAND2_X1 c2711(
.A1(net2804),
.A2(net2865),
.ZN(net2870)
);

OR4_X1 c2712(
.A1(net2868),
.A2(net2846),
.A3(net1892),
.A4(net11517),
.ZN(net2871)
);

NAND2_X2 c2713(
.A1(net2758),
.A2(net2870),
.ZN(net2872)
);

DFFS_X1 c2714(
.D(net1845),
.SN(net2871),
.CK(clk),
.Q(net2874),
.QN(net2873)
);

AND3_X2 c2715(
.A1(net849),
.A2(net1910),
.A3(net2847),
.ZN(net2875)
);

NOR3_X1 c2716(
.A1(net784),
.A2(net2865),
.A3(net914),
.ZN(net2876)
);

NAND2_X4 c2717(
.A1(net1697),
.A2(net2855),
.ZN(net2877)
);

OR3_X2 c2718(
.A1(net2832),
.A2(net1909),
.A3(net2734),
.ZN(net2878)
);

INV_X1 c2719(
.A(net10267),
.ZN(net2879)
);

AND2_X2 c2720(
.A1(net2785),
.A2(net2867),
.ZN(net2880)
);

XOR2_X1 c2721(
.A(net1594),
.B(net2816),
.Z(net2881)
);

SDFFR_X1 c2722(
.D(net2875),
.RN(net2877),
.SE(net2861),
.SI(net889),
.CK(clk),
.Q(net2883),
.QN(net2882)
);

NOR2_X1 c2723(
.A1(net2580),
.A2(net2823),
.ZN(net2884)
);

OR2_X2 c2724(
.A1(net2884),
.A2(net2594),
.ZN(net2885)
);

DFFRS_X2 c2725(
.D(net2885),
.RN(net2877),
.SN(net2882),
.CK(clk),
.Q(net2887),
.QN(net2886)
);

OAI221_X2 c2726(
.A(net2837),
.B1(net926),
.B2(net2880),
.C1(net2886),
.C2(net2861),
.ZN(net2888)
);

INV_X2 c2727(
.A(net9755),
.ZN(net2889)
);

OAI21_X2 c2728(
.A(net2856),
.B1(net2842),
.B2(net1697),
.ZN(net2890)
);

NOR2_X4 c2729(
.A1(net2886),
.A2(net10788),
.ZN(net2891)
);

NOR2_X2 c2730(
.A1(net2828),
.A2(net2890),
.ZN(net2892)
);

OAI21_X1 c2731(
.A(net1750),
.B1(net2887),
.B2(net2878),
.ZN(net2893)
);

XOR2_X2 c2732(
.A(net1647),
.B(net10787),
.Z(net2894)
);

SDFF_X1 c2733(
.D(net2871),
.SE(net1881),
.SI(net2894),
.CK(clk),
.Q(net2896),
.QN(net2895)
);

OAI22_X1 c2734(
.A1(net1838),
.A2(net2859),
.B1(net2877),
.B2(net2894),
.ZN(net2897)
);

AOI21_X2 c2735(
.A(net2865),
.B1(net2880),
.B2(net2891),
.ZN(net2898)
);

AOI21_X1 c2736(
.A(net2898),
.B1(net2889),
.B2(net2895),
.ZN(net2899)
);

AOI21_X4 c2737(
.A(net2899),
.B1(net2893),
.B2(net2755),
.ZN(net2900)
);

OAI222_X4 c2738(
.A1(net1807),
.A2(net2899),
.B1(net2894),
.B2(net863),
.C1(net2877),
.C2(net10536),
.ZN(net2901)
);

INV_X8 c2739(
.A(net1999),
.ZN(net2902)
);

INV_X16 c2740(
.A(net1972),
.ZN(net2903)
);

INV_X32 c2741(
.A(net963),
.ZN(net2904)
);

DFFS_X2 c2742(
.D(in24),
.SN(net1023),
.CK(clk),
.Q(net2906),
.QN(net2905)
);

INV_X4 c2743(
.A(net2904),
.ZN(net2907)
);

INV_X1 c2744(
.A(net1930),
.ZN(net2908)
);

INV_X2 c2745(
.A(net2903),
.ZN(net2909)
);

INV_X8 c2746(
.A(net2902),
.ZN(net2910)
);

XNOR2_X1 c2747(
.A(net960),
.B(net11510),
.ZN(net2911)
);

OR2_X4 c2748(
.A1(net968),
.A2(net2904),
.ZN(net2912)
);

OR2_X1 c2749(
.A1(net1924),
.A2(in7),
.ZN(net2913)
);

XNOR2_X2 c2750(
.A(net1957),
.B(net1994),
.ZN(net2914)
);

INV_X16 c2751(
.A(net14),
.ZN(net2915)
);

INV_X32 c2752(
.A(net969),
.ZN(net2916)
);

AND2_X4 c2753(
.A1(net963),
.A2(net1982),
.ZN(net2917)
);

AND3_X1 c2754(
.A1(net2910),
.A2(net2911),
.A3(net2916),
.ZN(net2918)
);

AND2_X1 c2755(
.A1(net2913),
.A2(net1933),
.ZN(net2919)
);

INV_X4 c2756(
.A(net2913),
.ZN(net2920)
);

INV_X1 c2757(
.A(net1946),
.ZN(net2921)
);

NAND2_X1 c2758(
.A1(net2916),
.A2(net11511),
.ZN(net2922)
);

NAND2_X2 c2759(
.A1(net2922),
.A2(net2903),
.ZN(net2923)
);

INV_X2 c2760(
.A(net1005),
.ZN(net2924)
);

NAND3_X1 c2761(
.A1(net2921),
.A2(net1930),
.A3(net1000),
.ZN(net2925)
);

INV_X8 c2762(
.A(net1982),
.ZN(net2926)
);

INV_X16 c2763(
.A(net1980),
.ZN(net2927)
);

NOR3_X4 c2764(
.A1(net2917),
.A2(net2924),
.A3(net33),
.ZN(net2928)
);

NAND2_X4 c2765(
.A1(net1999),
.A2(net2922),
.ZN(net2929)
);

INV_X32 c2766(
.A(net9661),
.ZN(net2930)
);

DFFR_X1 c2767(
.D(net2925),
.RN(net1936),
.CK(clk),
.Q(net2932),
.QN(net2931)
);

INV_X4 c2768(
.A(net9662),
.ZN(net2933)
);

NOR3_X2 c2769(
.A1(net2933),
.A2(net2919),
.A3(in24),
.ZN(net2934)
);

INV_X1 c2770(
.A(net1930),
.ZN(net2935)
);

AND2_X2 c2771(
.A1(net2916),
.A2(net1968),
.ZN(net2936)
);

AND3_X4 c2772(
.A1(net2934),
.A2(net2920),
.A3(net2926),
.ZN(net2937)
);

XOR2_X1 c2773(
.A(net2912),
.B(net2905),
.Z(net2938)
);

INV_X2 c2774(
.A(net2911),
.ZN(net2939)
);

NOR2_X1 c2775(
.A1(net1930),
.A2(net10692),
.ZN(net2940)
);

OR2_X2 c2776(
.A1(net2938),
.A2(net988),
.ZN(net2941)
);

INV_X8 c2777(
.A(net2930),
.ZN(net2942)
);

NOR2_X4 c2778(
.A1(net1995),
.A2(net1946),
.ZN(net2943)
);

INV_X16 c2779(
.A(net1005),
.ZN(net2944)
);

NOR2_X2 c2780(
.A1(net2920),
.A2(net2909),
.ZN(net2945)
);

XOR2_X2 c2781(
.A(net2908),
.B(net2919),
.Z(net2946)
);

INV_X32 c2782(
.A(net2914),
.ZN(net2947)
);

INV_X4 c2783(
.A(net2922),
.ZN(net2948)
);

XNOR2_X1 c2784(
.A(net2927),
.B(net2930),
.ZN(net2949)
);

OR2_X4 c2785(
.A1(net2945),
.A2(net2933),
.ZN(net2950)
);

OR2_X1 c2786(
.A1(net2950),
.A2(net10649),
.ZN(net2951)
);

XNOR2_X2 c2787(
.A(net1933),
.B(net10648),
.ZN(net2952)
);

INV_X1 c2788(
.A(net2918),
.ZN(net2953)
);

AND2_X4 c2789(
.A1(net2952),
.A2(net2946),
.ZN(net2954)
);

INV_X2 c2790(
.A(net2951),
.ZN(net2955)
);

SDFF_X2 c2791(
.D(net2939),
.SE(net2929),
.SI(net2931),
.CK(clk),
.Q(net2957),
.QN(net2956)
);

AND2_X1 c2792(
.A1(net2947),
.A2(net2936),
.ZN(net2958)
);

NAND3_X2 c2793(
.A1(net2940),
.A2(net2930),
.A3(net2933),
.ZN(net2959)
);

DFFR_X2 c2794(
.D(net2948),
.RN(net2932),
.CK(clk),
.Q(net2961),
.QN(net2960)
);

DFFRS_X1 c2795(
.D(net2957),
.RN(net2947),
.SN(net2958),
.CK(clk),
.Q(net2963),
.QN(net2962)
);

NAND2_X1 c2796(
.A1(net1920),
.A2(net2955),
.ZN(net2964)
);

DFFRS_X2 c2797(
.D(net2919),
.RN(net2953),
.SN(net2912),
.CK(clk),
.Q(net2966),
.QN(net2965)
);

NAND2_X2 c2798(
.A1(net2936),
.A2(net2925),
.ZN(net2967)
);

SDFF_X1 c2799(
.D(net2950),
.SE(net2963),
.SI(net2958),
.CK(clk),
.Q(net2969),
.QN(net2968)
);

DFFS_X1 c2800(
.D(net2959),
.SN(net2967),
.CK(clk),
.Q(net2971),
.QN(net2970)
);

NAND2_X4 c2801(
.A1(net2946),
.A2(net960),
.ZN(net2972)
);

SDFF_X2 c2802(
.D(net2932),
.SE(net2953),
.SI(net2956),
.CK(clk),
.Q(net2974),
.QN(net2973)
);

OR3_X1 c2803(
.A1(net2943),
.A2(net2970),
.A3(net2930),
.ZN(net2975)
);

MUX2_X1 c2804(
.A(net2955),
.B(net2910),
.S(net2968),
.Z(net2976)
);

OAI21_X4 c2805(
.A(net2937),
.B1(net2944),
.B2(net2917),
.ZN(net2977)
);

MUX2_X2 c2806(
.A(net2924),
.B(net2969),
.S(net2973),
.Z(net2978)
);

AND2_X2 c2807(
.A1(net2921),
.A2(net2914),
.ZN(net2979)
);

AND4_X2 c2808(
.A1(net2969),
.A2(net2975),
.A3(net2915),
.A4(net1915),
.ZN(net2980)
);

DFFRS_X1 c2809(
.D(net2953),
.RN(net2975),
.SN(net2977),
.CK(clk),
.Q(net2982),
.QN(net2981)
);

XOR2_X1 c2810(
.A(net2935),
.B(net2977),
.Z(net2983)
);

NOR2_X1 c2811(
.A1(net2975),
.A2(net1982),
.ZN(net2984)
);

NAND3_X4 c2812(
.A1(net2974),
.A2(net2981),
.A3(net2978),
.ZN(net2985)
);

OR2_X2 c2813(
.A1(net2977),
.A2(net2979),
.ZN(net2986)
);

NOR2_X4 c2814(
.A1(net2934),
.A2(net2978),
.ZN(net2987)
);

DFFS_X2 c2815(
.D(net1023),
.SN(net1978),
.CK(clk),
.Q(net2989),
.QN(net2988)
);

NOR2_X2 c2816(
.A1(net2978),
.A2(net2984),
.ZN(net2990)
);

DFFRS_X2 c2817(
.D(net1973),
.RN(net2959),
.SN(net2958),
.CK(clk),
.Q(net2992),
.QN(net2991)
);

XOR2_X2 c2818(
.A(net2982),
.B(net2984),
.Z(net2993)
);

AOI221_X4 c2819(
.A(net2939),
.B1(net2930),
.B2(net2977),
.C1(net2964),
.C2(net2987),
.ZN(net2994)
);

SDFFRS_X1 c2820(
.D(net2993),
.RN(net2977),
.SE(net2988),
.SI(net2987),
.SN(net2980),
.CK(clk),
.Q(net2996),
.QN(net2995)
);

XNOR2_X1 c2821(
.A(net2993),
.B(net10649),
.ZN(net2997)
);

OR2_X4 c2822(
.A1(net2915),
.A2(net2078),
.ZN(net2998)
);

INV_X8 c2823(
.A(net1038),
.ZN(net2999)
);

INV_X16 c2824(
.A(net2972),
.ZN(net3000)
);

DFFR_X1 c2825(
.D(net1109),
.RN(net2016),
.CK(clk),
.Q(net3002),
.QN(net3001)
);

INV_X32 c2826(
.A(net1067),
.ZN(net3003)
);

INV_X4 c2827(
.A(net2989),
.ZN(net3004)
);

OR2_X1 c2828(
.A1(net1968),
.A2(net2941),
.ZN(net3005)
);

INV_X1 c2829(
.A(net2027),
.ZN(net3006)
);

INV_X2 c2830(
.A(net1051),
.ZN(net3007)
);

INV_X8 c2831(
.A(net9680),
.ZN(net3008)
);

INV_X16 c2832(
.A(net2996),
.ZN(net3009)
);

INV_X32 c2833(
.A(net10932),
.ZN(net3010)
);

INV_X4 c2834(
.A(net2961),
.ZN(net3011)
);

INV_X1 c2835(
.A(net10623),
.ZN(net3012)
);

INV_X2 c2836(
.A(net2020),
.ZN(net3013)
);

INV_X8 c2837(
.A(net2944),
.ZN(net3014)
);

INV_X16 c2838(
.A(net3003),
.ZN(net3015)
);

INV_X32 c2839(
.A(net3013),
.ZN(net3016)
);

INV_X4 c2840(
.A(net3012),
.ZN(net3017)
);

XNOR2_X2 c2841(
.A(net2985),
.B(net3000),
.ZN(net3018)
);

INV_X1 c2842(
.A(net2992),
.ZN(net3019)
);

INV_X2 c2843(
.A(net9679),
.ZN(net3020)
);

INV_X8 c2844(
.A(net29),
.ZN(net3021)
);

INV_X16 c2845(
.A(net3015),
.ZN(net3022)
);

AND2_X4 c2846(
.A1(net2941),
.A2(net3015),
.ZN(net3023)
);

AND2_X1 c2847(
.A1(net3006),
.A2(net991),
.ZN(net3024)
);

INV_X32 c2848(
.A(net2971),
.ZN(net3025)
);

NAND2_X1 c2849(
.A1(net2072),
.A2(net3015),
.ZN(net3026)
);

OR3_X4 c2850(
.A1(net2056),
.A2(net3021),
.A3(net2991),
.ZN(net3027)
);

AND3_X2 c2851(
.A1(net2909),
.A2(net3001),
.A3(net3021),
.ZN(net3028)
);

NOR3_X1 c2852(
.A1(net3016),
.A2(net2096),
.A3(net2013),
.ZN(net3029)
);

NAND2_X2 c2853(
.A1(net3025),
.A2(net1951),
.ZN(net3030)
);

NAND2_X4 c2854(
.A1(net3012),
.A2(net2069),
.ZN(net3031)
);

INV_X4 c2855(
.A(net3021),
.ZN(net3032)
);

AND2_X2 c2856(
.A1(net2094),
.A2(net2964),
.ZN(net3033)
);

INV_X1 c2857(
.A(net2089),
.ZN(net3034)
);

INV_X2 c2858(
.A(net3014),
.ZN(net3035)
);

INV_X8 c2859(
.A(net9896),
.ZN(net3036)
);

INV_X16 c2860(
.A(net3007),
.ZN(net3037)
);

OR3_X2 c2861(
.A1(net3032),
.A2(net3015),
.A3(net1932),
.ZN(net3038)
);

INV_X32 c2862(
.A(net9878),
.ZN(net3039)
);

XOR2_X1 c2863(
.A(net3037),
.B(net78),
.Z(net3040)
);

INV_X4 c2864(
.A(net3024),
.ZN(net3041)
);

INV_X1 c2865(
.A(net3040),
.ZN(net3042)
);

INV_X2 c2866(
.A(net3020),
.ZN(net3043)
);

DFFR_X2 c2867(
.D(net3030),
.RN(net2958),
.CK(clk),
.Q(net3045),
.QN(net3044)
);

DFFS_X1 c2868(
.D(net3026),
.SN(net2077),
.CK(clk),
.Q(net3047),
.QN(net3046)
);

NOR2_X1 c2869(
.A1(net3041),
.A2(net3036),
.ZN(net3048)
);

OR2_X2 c2870(
.A1(net3019),
.A2(net10660),
.ZN(net3049)
);

NOR2_X4 c2871(
.A1(net2999),
.A2(net3036),
.ZN(net3050)
);

NOR2_X2 c2872(
.A1(net3034),
.A2(net3046),
.ZN(net3051)
);

INV_X8 c2873(
.A(net3042),
.ZN(net3052)
);

INV_X16 c2874(
.A(net9869),
.ZN(net3053)
);

XOR2_X2 c2875(
.A(net3029),
.B(net3019),
.Z(net3054)
);

INV_X32 c2876(
.A(net1957),
.ZN(net3055)
);

INV_X4 c2877(
.A(net3052),
.ZN(net3056)
);

XNOR2_X1 c2878(
.A(net3011),
.B(net3041),
.ZN(net3057)
);

SDFFR_X2 c2879(
.D(net3049),
.RN(net1118),
.SE(net2044),
.SI(net3038),
.CK(clk),
.Q(net3059),
.QN(net3058)
);

OR2_X4 c2880(
.A1(net3008),
.A2(net2960),
.ZN(net3060)
);

OR2_X1 c2881(
.A1(net3051),
.A2(net3036),
.ZN(net3061)
);

XNOR2_X2 c2882(
.A(net986),
.B(net2066),
.ZN(net3062)
);

INV_X1 c2883(
.A(net10100),
.ZN(net3063)
);

AND2_X4 c2884(
.A1(net3055),
.A2(net3059),
.ZN(net3064)
);

AND2_X1 c2885(
.A1(net3000),
.A2(net3064),
.ZN(net3065)
);

OAI21_X2 c2886(
.A(net3065),
.B1(net3053),
.B2(net2078),
.ZN(net3066)
);

NAND2_X1 c2887(
.A1(net3039),
.A2(net3064),
.ZN(net3067)
);

OAI21_X1 c2888(
.A(net2998),
.B1(net3031),
.B2(net3036),
.ZN(net3068)
);

NAND2_X2 c2889(
.A1(net1979),
.A2(net3067),
.ZN(net3069)
);

AOI21_X2 c2890(
.A(net3068),
.B1(net3035),
.B2(net2905),
.ZN(net3070)
);

NAND2_X4 c2891(
.A1(net3053),
.A2(net3069),
.ZN(net3071)
);

DFFS_X2 c2892(
.D(net3002),
.SN(net2083),
.CK(clk),
.Q(net3073),
.QN(net3072)
);

AND2_X2 c2893(
.A1(net2044),
.A2(net3061),
.ZN(net3074)
);

AOI21_X1 c2894(
.A(net3066),
.B1(net2029),
.B2(net3067),
.ZN(net3075)
);

XOR2_X1 c2895(
.A(net3036),
.B(net10820),
.Z(net3076)
);

SDFF_X1 c2896(
.D(net2038),
.SE(net3071),
.SI(net2962),
.CK(clk),
.Q(net3078),
.QN(net3077)
);

NOR2_X1 c2897(
.A1(net3075),
.A2(net3028),
.ZN(net3079)
);

OR2_X2 c2898(
.A1(net3078),
.A2(net3073),
.ZN(net3080)
);

AOI21_X4 c2899(
.A(net2033),
.B1(net3072),
.B2(net3080),
.ZN(net3081)
);

AND4_X1 c2900(
.A1(net3081),
.A2(net3022),
.A3(net3072),
.A4(net3080),
.ZN(net3082)
);

NOR2_X4 c2901(
.A1(net3077),
.A2(net10710),
.ZN(net3083)
);

OAI222_X2 c2902(
.A1(net3080),
.A2(net3073),
.B1(net3047),
.B2(net3071),
.C1(net3063),
.C2(net3004),
.ZN(net3084)
);

AOI222_X1 c2903(
.A1(net3076),
.A2(net3058),
.B1(net3017),
.B2(net3074),
.C1(net1996),
.C2(net3084),
.ZN(net3085)
);

AND3_X1 c2904(
.A1(net3057),
.A2(net3080),
.A3(net3084),
.ZN(net3086)
);

NOR2_X2 c2905(
.A1(net3045),
.A2(net3084),
.ZN(net3087)
);

AOI22_X4 c2906(
.A1(net2170),
.A2(net2997),
.B1(net2179),
.B2(net33),
.ZN(net3088)
);

INV_X2 c2907(
.A(net2101),
.ZN(net3089)
);

INV_X8 c2908(
.A(net2114),
.ZN(net3090)
);

INV_X16 c2909(
.A(net9776),
.ZN(net3091)
);

XOR2_X2 c2910(
.A(net3056),
.B(net2903),
.Z(net3092)
);

INV_X32 c2911(
.A(net9776),
.ZN(net3093)
);

INV_X4 c2912(
.A(net3090),
.ZN(net3094)
);

XNOR2_X1 c2913(
.A(net3089),
.B(net2122),
.ZN(net3095)
);

NAND3_X1 c2914(
.A1(net2164),
.A2(net1155),
.A3(net3019),
.ZN(net3096)
);

INV_X1 c2915(
.A(net2126),
.ZN(net3097)
);

INV_X2 c2916(
.A(net2051),
.ZN(net3098)
);

OR2_X4 c2917(
.A1(net3098),
.A2(net1193),
.ZN(net3099)
);

OR2_X1 c2918(
.A1(net3097),
.A2(net2051),
.ZN(net3100)
);

XNOR2_X2 c2919(
.A(net3094),
.B(net3067),
.ZN(net3101)
);

INV_X8 c2920(
.A(net10964),
.ZN(net3102)
);

INV_X16 c2921(
.A(net11285),
.ZN(net3103)
);

INV_X32 c2922(
.A(net3101),
.ZN(net3104)
);

AND2_X4 c2923(
.A1(net2171),
.A2(net2088),
.ZN(net3105)
);

INV_X4 c2924(
.A(net2078),
.ZN(net3106)
);

INV_X1 c2925(
.A(net2183),
.ZN(net3107)
);

INV_X2 c2926(
.A(net11361),
.ZN(net3108)
);

AND2_X1 c2927(
.A1(net3095),
.A2(net3104),
.ZN(net3109)
);

NAND2_X1 c2928(
.A1(net3071),
.A2(net2171),
.ZN(net3110)
);

INV_X8 c2929(
.A(net11170),
.ZN(net3111)
);

INV_X16 c2930(
.A(net3100),
.ZN(net3112)
);

INV_X32 c2931(
.A(net3110),
.ZN(net3113)
);

INV_X4 c2932(
.A(net3103),
.ZN(net3114)
);

INV_X1 c2933(
.A(net3111),
.ZN(net3115)
);

NAND2_X2 c2934(
.A1(net3115),
.A2(net3074),
.ZN(net3116)
);

INV_X2 c2935(
.A(net3109),
.ZN(net3117)
);

NAND2_X4 c2936(
.A1(net1155),
.A2(net2183),
.ZN(net3118)
);

INV_X8 c2937(
.A(net11418),
.ZN(net3119)
);

AND2_X2 c2938(
.A1(net2048),
.A2(net1996),
.ZN(net3120)
);

INV_X16 c2939(
.A(net10705),
.ZN(net3121)
);

XOR2_X1 c2940(
.A(net1169),
.B(net3112),
.Z(net3122)
);

INV_X32 c2941(
.A(net3102),
.ZN(net3123)
);

NOR2_X1 c2942(
.A1(net2907),
.A2(net11238),
.ZN(net3124)
);

OR2_X2 c2943(
.A1(net3121),
.A2(net3044),
.ZN(net3125)
);

INV_X4 c2944(
.A(net1996),
.ZN(net3126)
);

INV_X1 c2945(
.A(net9816),
.ZN(net3127)
);

NOR2_X4 c2946(
.A1(net3123),
.A2(net3120),
.ZN(net3128)
);

NOR2_X2 c2947(
.A1(net3091),
.A2(net2179),
.ZN(net3129)
);

XOR2_X2 c2948(
.A(net3067),
.B(net3128),
.Z(net3130)
);

XNOR2_X1 c2949(
.A(net2997),
.B(net3129),
.ZN(net3131)
);

INV_X2 c2950(
.A(net3130),
.ZN(net3132)
);

INV_X8 c2951(
.A(net3050),
.ZN(net3133)
);

OR2_X4 c2952(
.A1(net2958),
.A2(net191),
.ZN(net3134)
);

INV_X16 c2953(
.A(net11130),
.ZN(net3135)
);

INV_X32 c2954(
.A(net11048),
.ZN(net3136)
);

INV_X4 c2955(
.A(net11002),
.ZN(net3137)
);

NOR3_X4 c2956(
.A1(net3127),
.A2(net3126),
.A3(net3128),
.ZN(net3138)
);

OR2_X1 c2957(
.A1(net3138),
.A2(net3137),
.ZN(net3139)
);

XNOR2_X2 c2958(
.A(net3128),
.B(net3121),
.ZN(net3140)
);

NOR3_X2 c2959(
.A1(net3135),
.A2(net3113),
.A3(net3074),
.ZN(net3141)
);

AND2_X4 c2960(
.A1(net3137),
.A2(net3104),
.ZN(net3142)
);

INV_X1 c2961(
.A(net1101),
.ZN(net3143)
);

AND2_X1 c2962(
.A1(net3136),
.A2(net3127),
.ZN(net3144)
);

NAND2_X1 c2963(
.A1(net3106),
.A2(net3113),
.ZN(net3145)
);

NAND2_X2 c2964(
.A1(net3125),
.A2(net3129),
.ZN(net3146)
);

NAND2_X4 c2965(
.A1(net1047),
.A2(net3129),
.ZN(net3147)
);

AND2_X2 c2966(
.A1(net3131),
.A2(net3125),
.ZN(net3148)
);

INV_X2 c2967(
.A(net11107),
.ZN(net3149)
);

INV_X8 c2968(
.A(net10099),
.ZN(net3150)
);

AND3_X4 c2969(
.A1(net3105),
.A2(net3071),
.A3(net3108),
.ZN(net3151)
);

NAND3_X2 c2970(
.A1(net3019),
.A2(net3150),
.A3(net3023),
.ZN(net3152)
);

XOR2_X1 c2971(
.A(net1145),
.B(net2161),
.Z(net3153)
);

AOI221_X2 c2972(
.A(net3153),
.B1(net2183),
.B2(net2997),
.C1(net2144),
.C2(net3129),
.ZN(net3154)
);

NOR2_X1 c2973(
.A1(net3113),
.A2(net3154),
.ZN(net3155)
);

INV_X16 c2974(
.A(net3148),
.ZN(net3156)
);

OR2_X2 c2975(
.A1(net3140),
.A2(net3150),
.ZN(net3157)
);

OAI22_X4 c2976(
.A1(net189),
.A2(net3154),
.B1(net3156),
.B2(net2179),
.ZN(net3158)
);

NOR2_X4 c2977(
.A1(net3147),
.A2(net3120),
.ZN(net3159)
);

NOR2_X2 c2978(
.A1(net3141),
.A2(net3155),
.ZN(net3160)
);

INV_X32 c2979(
.A(net11272),
.ZN(net3161)
);

SDFF_X2 c2980(
.D(net3074),
.SE(net3139),
.SI(net3156),
.CK(clk),
.Q(net3163),
.QN(net3162)
);

OR3_X1 c2981(
.A1(net3145),
.A2(net3149),
.A3(net3162),
.ZN(net3164)
);

MUX2_X1 c2982(
.A(net3151),
.B(net1915),
.S(net3145),
.Z(net3165)
);

AOI221_X1 c2983(
.A(net3116),
.B1(net3133),
.B2(net3142),
.C1(net3128),
.C2(net3108),
.ZN(net3166)
);

OAI221_X1 c2984(
.A(net3107),
.B1(net3133),
.B2(net3161),
.C1(net3083),
.C2(net3108),
.ZN(net3167)
);

OAI21_X4 c2985(
.A(net3143),
.B1(net3150),
.B2(net3137),
.ZN(net3168)
);

DFFRS_X1 c2986(
.D(net3160),
.RN(net3128),
.SN(net10661),
.CK(clk),
.Q(net3170),
.QN(net3169)
);

MUX2_X2 c2987(
.A(net3159),
.B(net3148),
.S(net3170),
.Z(net3171)
);

XOR2_X2 c2988(
.A(net2263),
.B(net2169),
.Z(net3172)
);

XNOR2_X1 c2989(
.A(net3114),
.B(net2227),
.ZN(net3173)
);

INV_X4 c2990(
.A(net3069),
.ZN(net3174)
);

INV_X1 c2991(
.A(net2197),
.ZN(net3175)
);

OR2_X4 c2992(
.A1(net2092),
.A2(net2238),
.ZN(net3176)
);

OR2_X1 c2993(
.A1(net272),
.A2(net1229),
.ZN(net3177)
);

XNOR2_X2 c2994(
.A(net3175),
.B(net2189),
.ZN(net3178)
);

INV_X2 c2995(
.A(net3144),
.ZN(net3179)
);

INV_X8 c2996(
.A(net3142),
.ZN(net3180)
);

AND2_X4 c2997(
.A1(net1288),
.A2(net11237),
.ZN(net3181)
);

INV_X16 c2998(
.A(net10265),
.ZN(net3182)
);

INV_X32 c2999(
.A(net11309),
.ZN(net3183)
);

NAND3_X4 c3000(
.A1(net3180),
.A2(net3142),
.A3(net3169),
.ZN(net3184)
);

AND2_X1 c3001(
.A1(net2169),
.A2(net3069),
.ZN(net3185)
);

OR3_X4 c3002(
.A1(net3172),
.A2(net1229),
.A3(net11321),
.ZN(net3186)
);

NAND2_X1 c3003(
.A1(net1922),
.A2(net3163),
.ZN(net3187)
);

NAND2_X2 c3004(
.A1(net2192),
.A2(net78),
.ZN(net3188)
);

NAND2_X4 c3005(
.A1(net1035),
.A2(net3171),
.ZN(net3189)
);

AND2_X2 c3006(
.A1(net3185),
.A2(net3182),
.ZN(net3190)
);

INV_X4 c3007(
.A(net11309),
.ZN(net3191)
);

XOR2_X1 c3008(
.A(net2196),
.B(net1220),
.Z(net3192)
);

INV_X1 c3009(
.A(net3176),
.ZN(net3193)
);

NOR2_X1 c3010(
.A1(net3146),
.A2(net2023),
.ZN(net3194)
);

OR2_X2 c3011(
.A1(net2238),
.A2(net11269),
.ZN(net3195)
);

NOR2_X4 c3012(
.A1(net2255),
.A2(net2197),
.ZN(net3196)
);

NOR2_X2 c3013(
.A1(net3196),
.A2(net1288),
.ZN(net3197)
);

INV_X2 c3014(
.A(net10330),
.ZN(net3198)
);

DFFR_X1 c3015(
.D(net3157),
.RN(net3198),
.CK(clk),
.Q(net3200),
.QN(net3199)
);

INV_X8 c3016(
.A(net10488),
.ZN(net3201)
);

XOR2_X2 c3017(
.A(net2238),
.B(net3162),
.Z(net3202)
);

INV_X16 c3018(
.A(net3183),
.ZN(net3203)
);

INV_X32 c3019(
.A(net11327),
.ZN(net3204)
);

AND3_X2 c3020(
.A1(net999),
.A2(net3158),
.A3(net3167),
.ZN(net3205)
);

DFFRS_X2 c3021(
.D(net3154),
.RN(net2241),
.SN(net11139),
.CK(clk),
.Q(net3207),
.QN(net3206)
);

XNOR2_X1 c3022(
.A(net1195),
.B(net285),
.ZN(net3208)
);

INV_X4 c3023(
.A(net9991),
.ZN(net3209)
);

INV_X1 c3024(
.A(net11092),
.ZN(net3210)
);

OR2_X4 c3025(
.A1(net3181),
.A2(net11269),
.ZN(net3211)
);

INV_X2 c3026(
.A(net11270),
.ZN(net3212)
);

OAI221_X4 c3027(
.A(net3203),
.B1(net3202),
.B2(net3162),
.C1(net3004),
.C2(net2192),
.ZN(net3213)
);

OR2_X1 c3028(
.A1(net2189),
.A2(net3213),
.ZN(net3214)
);

XNOR2_X2 c3029(
.A(net3188),
.B(net3210),
.ZN(net3215)
);

AND2_X4 c3030(
.A1(net3204),
.A2(net3083),
.ZN(net3216)
);

AND2_X1 c3031(
.A1(net2903),
.A2(net3156),
.ZN(net3217)
);

SDFFRS_X2 c3032(
.D(net3190),
.RN(net283),
.SE(net3217),
.SI(net3201),
.SN(net11321),
.CK(clk),
.Q(net3219),
.QN(net3218)
);

INV_X8 c3033(
.A(net191),
.ZN(net3220)
);

NAND2_X1 c3034(
.A1(net2274),
.A2(net3216),
.ZN(net3221)
);

NAND2_X2 c3035(
.A1(net3202),
.A2(net3198),
.ZN(net3222)
);

NAND2_X4 c3036(
.A1(net3083),
.A2(net3218),
.ZN(net3223)
);

NOR3_X1 c3037(
.A1(net3212),
.A2(net2144),
.A3(net2016),
.ZN(net3224)
);

AND2_X2 c3038(
.A1(net3213),
.A2(net3206),
.ZN(net3225)
);

OR3_X2 c3039(
.A1(net3221),
.A2(net2238),
.A3(net3223),
.ZN(net3226)
);

XOR2_X1 c3040(
.A(net3220),
.B(net3219),
.Z(net3227)
);

NOR2_X1 c3041(
.A1(net3194),
.A2(net3200),
.ZN(net3228)
);

OAI21_X2 c3042(
.A(net3224),
.B1(net3217),
.B2(net3201),
.ZN(net3229)
);

OR2_X2 c3043(
.A1(net3173),
.A2(net1253),
.ZN(net3230)
);

NOR2_X4 c3044(
.A1(net3126),
.A2(net3220),
.ZN(net3231)
);

NOR2_X2 c3045(
.A1(net3215),
.A2(net3171),
.ZN(net3232)
);

XOR2_X2 c3046(
.A(net3222),
.B(net3212),
.Z(net3233)
);

OAI21_X1 c3047(
.A(net3230),
.B1(net3206),
.B2(net11200),
.ZN(net3234)
);

AOI21_X2 c3048(
.A(net2029),
.B1(net3213),
.B2(net3146),
.ZN(net3235)
);

AOI21_X1 c3049(
.A(net1253),
.B1(net3231),
.B2(net3201),
.ZN(net3236)
);

XNOR2_X1 c3050(
.A(net3195),
.B(net3235),
.ZN(net3237)
);

INV_X16 c3051(
.A(net11069),
.ZN(net3238)
);

AOI21_X4 c3052(
.A(net3234),
.B1(net2069),
.B2(net3238),
.ZN(net3239)
);

SDFFRS_X1 c3053(
.D(net3210),
.RN(net3217),
.SE(net3069),
.SI(net2192),
.SN(net3129),
.CK(clk),
.Q(net3241),
.QN(net3240)
);

SDFF_X1 c3054(
.D(net3227),
.SE(net3241),
.SI(net3237),
.CK(clk),
.Q(net3243),
.QN(net3242)
);

AND3_X1 c3055(
.A1(net3187),
.A2(net3220),
.A3(net3173),
.ZN(net3244)
);

OR2_X4 c3056(
.A1(net3233),
.A2(net3216),
.ZN(net3245)
);

OAI221_X2 c3057(
.A(net3244),
.B1(net3230),
.B2(net3228),
.C1(net3182),
.C2(net3242),
.ZN(net3246)
);

OR2_X1 c3058(
.A1(net3228),
.A2(net11200),
.ZN(net3247)
);

NAND3_X1 c3059(
.A1(net3239),
.A2(net3177),
.A3(net3083),
.ZN(net3248)
);

SDFF_X2 c3060(
.D(net3236),
.SE(net3247),
.SI(net2903),
.CK(clk),
.Q(net3250),
.QN(net3249)
);

SDFFRS_X2 c3061(
.D(net3198),
.RN(net3204),
.SE(net1253),
.SI(net3240),
.SN(net3217),
.CK(clk),
.Q(net3252),
.QN(net3251)
);

NOR3_X4 c3062(
.A1(net3231),
.A2(net3170),
.A3(net3223),
.ZN(net3253)
);

AOI222_X4 c3063(
.A1(net3250),
.A2(net3238),
.B1(net3236),
.B2(net3242),
.C1(net3054),
.C2(net3201),
.ZN(net3254)
);

NOR3_X2 c3064(
.A1(net3219),
.A2(net3250),
.A3(net3237),
.ZN(net3255)
);

AND3_X4 c3065(
.A1(net3225),
.A2(net3142),
.A3(net3231),
.ZN(net3256)
);

DFFR_X2 c3066(
.D(net3254),
.RN(net3237),
.CK(clk),
.Q(net3258),
.QN(net3257)
);

INV_X32 c3067(
.A(net11277),
.ZN(net3259)
);

OAI33_X1 c3068(
.A1(net3214),
.A2(net3252),
.A3(net1915),
.B1(net3256),
.B2(net3259),
.B3(net3249),
.ZN(net3260)
);

XNOR2_X2 c3069(
.A(net3179),
.B(net3259),
.ZN(net3261)
);

AOI222_X2 c3070(
.A1(net3246),
.A2(net3168),
.B1(net3257),
.B2(net3259),
.C1(net3198),
.C2(net11344),
.ZN(net3262)
);

INV_X4 c3071(
.A(net2332),
.ZN(net3263)
);

INV_X1 c3072(
.A(net11473),
.ZN(net3264)
);

INV_X2 c3073(
.A(net11069),
.ZN(net3265)
);

INV_X8 c3074(
.A(net2240),
.ZN(net3266)
);

INV_X16 c3075(
.A(net3124),
.ZN(net3267)
);

AND2_X4 c3076(
.A1(net2306),
.A2(net3240),
.ZN(net3268)
);

INV_X32 c3077(
.A(net2179),
.ZN(net3269)
);

NAND3_X2 c3078(
.A1(net372),
.A2(net2023),
.A3(net2235),
.ZN(net3270)
);

AND2_X1 c3079(
.A1(net352),
.A2(net2326),
.ZN(net3271)
);

INV_X4 c3080(
.A(net2327),
.ZN(net3272)
);

NAND2_X1 c3081(
.A1(net2354),
.A2(net2254),
.ZN(net3273)
);

NAND2_X2 c3082(
.A1(net2346),
.A2(net2023),
.ZN(net3274)
);

INV_X1 c3083(
.A(net1351),
.ZN(net3275)
);

INV_X2 c3084(
.A(net9664),
.ZN(net3276)
);

NAND2_X4 c3085(
.A1(net2338),
.A2(net3242),
.ZN(net3277)
);

AND2_X2 c3086(
.A1(net3241),
.A2(net3177),
.ZN(net3278)
);

XOR2_X1 c3087(
.A(net3271),
.B(net2235),
.Z(net3279)
);

INV_X8 c3088(
.A(net3266),
.ZN(net3280)
);

INV_X16 c3089(
.A(net3272),
.ZN(net3281)
);

INV_X32 c3090(
.A(net9663),
.ZN(net3282)
);

INV_X4 c3091(
.A(net3267),
.ZN(net3283)
);

OR3_X1 c3092(
.A1(net3243),
.A2(net3276),
.A3(net11279),
.ZN(net3284)
);

INV_X1 c3093(
.A(net2069),
.ZN(net3285)
);

NOR2_X1 c3094(
.A1(net2335),
.A2(net11468),
.ZN(net3286)
);

INV_X2 c3095(
.A(net11233),
.ZN(net3287)
);

INV_X8 c3096(
.A(net3213),
.ZN(net3288)
);

OR2_X2 c3097(
.A1(net2191),
.A2(net3265),
.ZN(net3289)
);

MUX2_X1 c3098(
.A(net3275),
.B(net3126),
.S(net2069),
.Z(net3290)
);

INV_X16 c3099(
.A(net10424),
.ZN(net3291)
);

NOR2_X4 c3100(
.A1(net3178),
.A2(net2235),
.ZN(net3292)
);

INV_X32 c3101(
.A(net3287),
.ZN(net3293)
);

OAI21_X4 c3102(
.A(net3274),
.B1(net2323),
.B2(net3192),
.ZN(net3294)
);

SDFFS_X1 c3103(
.D(net3285),
.SE(net2327),
.SI(net3192),
.SN(net11513),
.CK(clk),
.Q(net3296),
.QN(net3295)
);

INV_X4 c3104(
.A(net9850),
.ZN(net3297)
);

MUX2_X2 c3105(
.A(net3269),
.B(net2191),
.S(net2332),
.Z(net3298)
);

NAND3_X4 c3106(
.A1(net2928),
.A2(net2276),
.A3(net11303),
.ZN(net3299)
);

OR3_X4 c3107(
.A1(net1270),
.A2(net3286),
.A3(net3291),
.ZN(net3300)
);

AND3_X2 c3108(
.A1(net3300),
.A2(net2332),
.A3(net3287),
.ZN(net3301)
);

NOR2_X2 c3109(
.A1(net2346),
.A2(net11168),
.ZN(net3302)
);

INV_X1 c3110(
.A(net3171),
.ZN(net3303)
);

INV_X2 c3111(
.A(net9828),
.ZN(net3304)
);

DFFS_X1 c3112(
.D(net3245),
.SN(net3267),
.CK(clk),
.Q(net3306),
.QN(net3305)
);

INV_X8 c3113(
.A(net2023),
.ZN(net3307)
);

INV_X16 c3114(
.A(net3282),
.ZN(net3308)
);

XOR2_X2 c3115(
.A(net3304),
.B(net2277),
.Z(net3309)
);

XNOR2_X1 c3116(
.A(net3288),
.B(net3291),
.ZN(net3310)
);

DFFS_X2 c3117(
.D(net3298),
.SN(net3237),
.CK(clk),
.Q(net3312),
.QN(net3311)
);

INV_X32 c3118(
.A(net3279),
.ZN(net3313)
);

OR2_X4 c3119(
.A1(net3313),
.A2(net3307),
.ZN(net3314)
);

OR2_X1 c3120(
.A1(net3286),
.A2(net3314),
.ZN(net3315)
);

NOR3_X1 c3121(
.A1(net2340),
.A2(net1217),
.A3(net3279),
.ZN(net3316)
);

AOI22_X2 c3122(
.A1(net3315),
.A2(net3228),
.B1(net3266),
.B2(net3308),
.ZN(net3317)
);

XNOR2_X2 c3123(
.A(net3283),
.B(net1297),
.ZN(net3318)
);

DFFR_X1 c3124(
.D(net3289),
.RN(net3317),
.CK(clk),
.Q(net3320),
.QN(net3319)
);

INV_X4 c3125(
.A(net2290),
.ZN(net3321)
);

OR3_X2 c3126(
.A1(net3284),
.A2(net2333),
.A3(net3313),
.ZN(net3322)
);

OAI21_X2 c3127(
.A(net1338),
.B1(net3287),
.B2(net3308),
.ZN(net3323)
);

INV_X1 c3128(
.A(net11109),
.ZN(net3324)
);

OAI21_X1 c3129(
.A(net3318),
.B1(net3201),
.B2(net3282),
.ZN(net3325)
);

DFFRS_X1 c3130(
.D(net3299),
.RN(net1247),
.SN(net2338),
.CK(clk),
.Q(net3327),
.QN(net3326)
);

AND2_X4 c3131(
.A1(net3265),
.A2(net3307),
.ZN(net3328)
);

AND2_X1 c3132(
.A1(net3278),
.A2(net3279),
.ZN(net3329)
);

AOI21_X2 c3133(
.A(net3290),
.B1(net3201),
.B2(net3319),
.ZN(net3330)
);

AOI21_X1 c3134(
.A(net3307),
.B1(net3324),
.B2(net3299),
.ZN(net3331)
);

NAND2_X1 c3135(
.A1(net3324),
.A2(net1270),
.ZN(net3332)
);

NAND2_X2 c3136(
.A1(net3301),
.A2(net3297),
.ZN(net3333)
);

NAND2_X4 c3137(
.A1(net2308),
.A2(net11168),
.ZN(net3334)
);

AOI21_X4 c3138(
.A(net3332),
.B1(net3328),
.B2(net2351),
.ZN(net3335)
);

DFFRS_X2 c3139(
.D(net3303),
.RN(net2280),
.SN(net3271),
.CK(clk),
.Q(net3337),
.QN(net3336)
);

AND2_X2 c3140(
.A1(net3316),
.A2(net3297),
.ZN(net3338)
);

XOR2_X1 c3141(
.A(net3321),
.B(net11246),
.Z(net3339)
);

NOR2_X1 c3142(
.A1(net3323),
.A2(net3171),
.ZN(net3340)
);

OR2_X2 c3143(
.A1(net3308),
.A2(net3329),
.ZN(net3341)
);

AND3_X1 c3144(
.A1(net3339),
.A2(net3336),
.A3(net3323),
.ZN(net3342)
);

NAND3_X1 c3145(
.A1(net3342),
.A2(net3311),
.A3(net3295),
.ZN(net3343)
);

NOR2_X4 c3146(
.A1(net3302),
.A2(net3228),
.ZN(net3344)
);

SDFF_X1 c3147(
.D(net3344),
.SE(net3343),
.SI(net3251),
.CK(clk),
.Q(net3346),
.QN(net3345)
);

NOR3_X4 c3148(
.A1(net3343),
.A2(net3320),
.A3(net3271),
.ZN(net3347)
);

NOR3_X2 c3149(
.A1(net3281),
.A2(net3266),
.A3(net3341),
.ZN(net3348)
);

AND3_X4 c3150(
.A1(net3337),
.A2(net3346),
.A3(net3302),
.ZN(net3349)
);

NOR2_X2 c3151(
.A1(net3329),
.A2(net3348),
.ZN(net3350)
);

OAI222_X1 c3152(
.A1(net3350),
.A2(net3330),
.B1(net3349),
.B2(net3308),
.C1(net3319),
.C2(net3341),
.ZN(net3351)
);

NAND4_X4 c3153(
.A1(net3348),
.A2(net3337),
.A3(net3332),
.A4(net3341),
.ZN(net3352)
);

INV_X2 c3154(
.A(net11486),
.ZN(net3353)
);

INV_X8 c3155(
.A(net2235),
.ZN(net3354)
);

XOR2_X2 c3156(
.A(net1225),
.B(net3129),
.Z(net3355)
);

INV_X16 c3157(
.A(net11214),
.ZN(net3356)
);

INV_X32 c3158(
.A(net11068),
.ZN(net3357)
);

XNOR2_X1 c3159(
.A(net344),
.B(net3319),
.ZN(net3358)
);

INV_X4 c3160(
.A(net11206),
.ZN(net3359)
);

NAND3_X2 c3161(
.A1(net2410),
.A2(net3332),
.A3(net3358),
.ZN(net3360)
);

INV_X1 c3162(
.A(net10362),
.ZN(net3361)
);

INV_X2 c3163(
.A(net3360),
.ZN(net3362)
);

OR2_X4 c3164(
.A1(net2389),
.A2(net2438),
.ZN(net3363)
);

OR2_X1 c3165(
.A1(net428),
.A2(net2347),
.ZN(net3364)
);

INV_X8 c3166(
.A(net2347),
.ZN(net3365)
);

XNOR2_X2 c3167(
.A(net2412),
.B(net3356),
.ZN(net3366)
);

AND2_X4 c3168(
.A1(net2443),
.A2(net3356),
.ZN(net3367)
);

AND2_X1 c3169(
.A1(net3363),
.A2(net1361),
.ZN(net3368)
);

INV_X16 c3170(
.A(net3366),
.ZN(net3369)
);

INV_X32 c3171(
.A(net3357),
.ZN(net3370)
);

OR3_X1 c3172(
.A1(net1464),
.A2(net3363),
.A3(net3177),
.ZN(net3371)
);

INV_X4 c3173(
.A(net9719),
.ZN(net3372)
);

INV_X1 c3174(
.A(net3293),
.ZN(net3373)
);

INV_X2 c3175(
.A(net3370),
.ZN(net3374)
);

INV_X8 c3176(
.A(net2441),
.ZN(net3375)
);

MUX2_X1 c3177(
.A(net3177),
.B(net2447),
.S(net2420),
.Z(net3376)
);

NAND2_X1 c3178(
.A1(net3338),
.A2(net3322),
.ZN(net3377)
);

INV_X16 c3179(
.A(net3358),
.ZN(net3378)
);

INV_X32 c3180(
.A(net2434),
.ZN(net3379)
);

INV_X4 c3181(
.A(net3369),
.ZN(net3380)
);

OAI21_X4 c3182(
.A(net2433),
.B1(net3334),
.B2(net2410),
.ZN(net3381)
);

INV_X1 c3183(
.A(net10235),
.ZN(net3382)
);

INV_X2 c3184(
.A(net11513),
.ZN(net3383)
);

NAND2_X2 c3185(
.A1(net3353),
.A2(net3322),
.ZN(net3384)
);

OAI222_X4 c3186(
.A1(net2345),
.A2(net3354),
.B1(net3345),
.B2(net3383),
.C1(net2351),
.C2(net2386),
.ZN(net3385)
);

MUX2_X2 c3187(
.A(net369),
.B(net2379),
.S(net11289),
.Z(net3386)
);

INV_X8 c3188(
.A(net10014),
.ZN(net3387)
);

INV_X16 c3189(
.A(net10086),
.ZN(net3388)
);

NAND2_X4 c3190(
.A1(net2317),
.A2(net3375),
.ZN(net3389)
);

AND2_X2 c3191(
.A1(net3380),
.A2(net3370),
.ZN(net3390)
);

XOR2_X1 c3192(
.A(net3377),
.B(net2434),
.Z(net3391)
);

INV_X32 c3193(
.A(net9828),
.ZN(net3392)
);

NOR2_X1 c3194(
.A1(net3375),
.A2(net2434),
.ZN(net3393)
);

INV_X4 c3195(
.A(net11274),
.ZN(net3394)
);

OR2_X2 c3196(
.A1(net3384),
.A2(net3383),
.ZN(net3395)
);

NOR2_X4 c3197(
.A1(net3394),
.A2(net3376),
.ZN(net3396)
);

NOR2_X2 c3198(
.A1(net3396),
.A2(net3384),
.ZN(net3397)
);

XOR2_X2 c3199(
.A(net3392),
.B(net2390),
.Z(net3398)
);

INV_X1 c3200(
.A(net3383),
.ZN(net3399)
);

XNOR2_X1 c3201(
.A(net3387),
.B(net428),
.ZN(net3400)
);

OR2_X4 c3202(
.A1(net3376),
.A2(net3383),
.ZN(net3401)
);

OR2_X1 c3203(
.A1(net3389),
.A2(net3382),
.ZN(net3402)
);

INV_X2 c3204(
.A(net10965),
.ZN(net3403)
);

OAI211_X2 c3205(
.A(net3401),
.B(net3359),
.C1(net2388),
.C2(net3397),
.ZN(net3404)
);

INV_X8 c3206(
.A(net10767),
.ZN(net3405)
);

INV_X16 c3207(
.A(net3386),
.ZN(net3406)
);

XNOR2_X2 c3208(
.A(net3388),
.B(net2440),
.ZN(net3407)
);

AND2_X4 c3209(
.A1(net3395),
.A2(net1353),
.ZN(net3408)
);

OR4_X2 c3210(
.A1(net3192),
.A2(net3401),
.A3(net3226),
.A4(net3308),
.ZN(net3409)
);

INV_X32 c3211(
.A(net3402),
.ZN(net3410)
);

AND2_X1 c3212(
.A1(net1401),
.A2(net3389),
.ZN(net3411)
);

INV_X4 c3213(
.A(net3398),
.ZN(net3412)
);

AOI221_X4 c3214(
.A(net3403),
.B1(net3408),
.B2(net3360),
.C1(net3346),
.C2(net3369),
.ZN(net3413)
);

INV_X1 c3215(
.A(net11272),
.ZN(net3414)
);

OAI222_X2 c3216(
.A1(net3412),
.A2(net3414),
.B1(net2434),
.B2(net1401),
.C1(net2241),
.C2(net3341),
.ZN(net3415)
);

NAND3_X4 c3217(
.A1(net2450),
.A2(net10725),
.A3(net11274),
.ZN(net3416)
);

NAND2_X1 c3218(
.A1(net428),
.A2(net11289),
.ZN(net3417)
);

INV_X2 c3219(
.A(net3381),
.ZN(net3418)
);

INV_X8 c3220(
.A(net10236),
.ZN(net3419)
);

INV_X16 c3221(
.A(net3322),
.ZN(net3420)
);

OR3_X4 c3222(
.A1(net3419),
.A2(net3377),
.A3(net3370),
.ZN(net3421)
);

NAND2_X2 c3223(
.A1(net3421),
.A2(net11139),
.ZN(net3422)
);

NAND2_X4 c3224(
.A1(net3406),
.A2(net11476),
.ZN(net3423)
);

INV_X32 c3225(
.A(net9719),
.ZN(net3424)
);

AND2_X2 c3226(
.A1(net3347),
.A2(net3386),
.ZN(net3425)
);

XOR2_X1 c3227(
.A(net3421),
.B(net3420),
.Z(net3426)
);

INV_X4 c3228(
.A(net3361),
.ZN(net3427)
);

NOR2_X1 c3229(
.A1(net3420),
.A2(net3177),
.ZN(net3428)
);

AND3_X2 c3230(
.A1(net3427),
.A2(net2390),
.A3(net344),
.ZN(net3429)
);

INV_X1 c3231(
.A(net11214),
.ZN(net3430)
);

NOR3_X1 c3232(
.A1(net2447),
.A2(net3429),
.A3(net3308),
.ZN(net3431)
);

INV_X2 c3233(
.A(net11222),
.ZN(net3432)
);

OR3_X2 c3234(
.A1(net3399),
.A2(net3432),
.A3(net3405),
.ZN(net3433)
);

OR2_X2 c3235(
.A1(net3430),
.A2(net3432),
.ZN(net3434)
);

NOR2_X4 c3236(
.A1(net3434),
.A2(net11303),
.ZN(net3435)
);

INV_X8 c3237(
.A(net3374),
.ZN(net3436)
);

INV_X16 c3238(
.A(net3173),
.ZN(net3437)
);

NOR2_X2 c3239(
.A1(net3320),
.A2(net2438),
.ZN(net3438)
);

XOR2_X2 c3240(
.A(net2515),
.B(net2491),
.Z(net3439)
);

XNOR2_X1 c3241(
.A(net1374),
.B(net3437),
.ZN(net3440)
);

INV_X32 c3242(
.A(net1514),
.ZN(net3441)
);

INV_X4 c3243(
.A(net1386),
.ZN(net3442)
);

OR2_X4 c3244(
.A1(net3438),
.A2(net1475),
.ZN(net3443)
);

INV_X1 c3245(
.A(net3436),
.ZN(net3444)
);

OR2_X1 c3246(
.A1(net3280),
.A2(net2379),
.ZN(net3445)
);

INV_X2 c3247(
.A(net10340),
.ZN(net3446)
);

OAI21_X2 c3248(
.A(net3362),
.B1(net2533),
.B2(net3340),
.ZN(net3447)
);

XNOR2_X2 c3249(
.A(net3346),
.B(net3405),
.ZN(net3448)
);

AND2_X4 c3250(
.A1(net3444),
.A2(net3264),
.ZN(net3449)
);

INV_X8 c3251(
.A(net2506),
.ZN(net3450)
);

SDFF_X2 c3252(
.D(net3375),
.SE(net3423),
.SI(net3354),
.CK(clk),
.Q(net3452),
.QN(net3451)
);

AND2_X1 c3253(
.A1(net2390),
.A2(net1491),
.ZN(net3453)
);

INV_X16 c3254(
.A(net2272),
.ZN(net3454)
);

INV_X32 c3255(
.A(net11058),
.ZN(net3455)
);

INV_X4 c3256(
.A(net9752),
.ZN(net3456)
);

INV_X1 c3257(
.A(net11246),
.ZN(net3457)
);

NAND2_X1 c3258(
.A1(net3372),
.A2(net11519),
.ZN(net3458)
);

NAND2_X2 c3259(
.A1(net3449),
.A2(net3448),
.ZN(net3459)
);

INV_X2 c3260(
.A(net11192),
.ZN(net3460)
);

INV_X8 c3261(
.A(net10589),
.ZN(net3461)
);

NAND2_X4 c3262(
.A1(net3461),
.A2(net3454),
.ZN(net3462)
);

INV_X16 c3263(
.A(net3438),
.ZN(net3463)
);

AND2_X2 c3264(
.A1(net3378),
.A2(net11518),
.ZN(net3464)
);

INV_X32 c3265(
.A(net3462),
.ZN(net3465)
);

XOR2_X1 c3266(
.A(net2545),
.B(net1527),
.Z(net3466)
);

NOR2_X1 c3267(
.A1(net2323),
.A2(net3428),
.ZN(net3467)
);

OR2_X2 c3268(
.A1(net3320),
.A2(net3454),
.ZN(net3468)
);

INV_X4 c3269(
.A(net2494),
.ZN(net3469)
);

NOR2_X4 c3270(
.A1(net3439),
.A2(net1412),
.ZN(net3470)
);

INV_X1 c3271(
.A(net10464),
.ZN(net3471)
);

NOR2_X2 c3272(
.A1(net3465),
.A2(net3464),
.ZN(net3472)
);

XOR2_X2 c3273(
.A(net3437),
.B(net2542),
.Z(net3473)
);

XNOR2_X1 c3274(
.A(net346),
.B(net3438),
.ZN(net3474)
);

OR2_X4 c3275(
.A1(net3325),
.A2(net3448),
.ZN(net3475)
);

OR2_X1 c3276(
.A1(net3456),
.A2(net2517),
.ZN(net3476)
);

XNOR2_X2 c3277(
.A(net3472),
.B(net2534),
.ZN(net3477)
);

INV_X2 c3278(
.A(net10130),
.ZN(net3478)
);

OAI21_X1 c3279(
.A(net3467),
.B1(net2490),
.B2(net3393),
.ZN(net3479)
);

AND2_X4 c3280(
.A1(net3441),
.A2(net10728),
.ZN(net3480)
);

INV_X8 c3281(
.A(net2438),
.ZN(net3481)
);

AOI21_X2 c3282(
.A(net3468),
.B1(net2271),
.B2(net3470),
.ZN(net3482)
);

AND2_X1 c3283(
.A1(net3481),
.A2(net2545),
.ZN(net3483)
);

INV_X16 c3284(
.A(net9751),
.ZN(net3484)
);

AOI21_X1 c3285(
.A(net3428),
.B1(net2506),
.B2(net3477),
.ZN(net3485)
);

AOI21_X4 c3286(
.A(net3475),
.B1(net3448),
.B2(net538),
.ZN(net3486)
);

AND3_X1 c3287(
.A1(net3485),
.A2(net1475),
.A3(net1386),
.ZN(net3487)
);

SDFFS_X2 c3288(
.D(net3486),
.SE(net3453),
.SI(net3418),
.SN(net3345),
.CK(clk),
.Q(net3489),
.QN(net3488)
);

NAND3_X1 c3289(
.A1(net538),
.A2(net3489),
.A3(net3477),
.ZN(net3490)
);

NAND2_X1 c3290(
.A1(net1475),
.A2(net3437),
.ZN(net3491)
);

NAND2_X2 c3291(
.A1(net2526),
.A2(net11370),
.ZN(net3492)
);

INV_X32 c3292(
.A(net10470),
.ZN(net3493)
);

INV_X4 c3293(
.A(net10320),
.ZN(net3494)
);

NOR3_X4 c3294(
.A1(net3483),
.A2(net3453),
.A3(net3460),
.ZN(net3495)
);

NAND2_X4 c3295(
.A1(net3450),
.A2(net1514),
.ZN(net3496)
);

INV_X1 c3296(
.A(net3480),
.ZN(net3497)
);

AND2_X2 c3297(
.A1(net3459),
.A2(net1504),
.ZN(net3498)
);

XOR2_X1 c3298(
.A(net2506),
.B(net11251),
.Z(net3499)
);

INV_X2 c3299(
.A(net10350),
.ZN(net3500)
);

NOR2_X1 c3300(
.A1(net3500),
.A2(net3498),
.ZN(net3501)
);

AOI211_X1 c3301(
.A(net1479),
.B(net3418),
.C1(net3454),
.C2(net3498),
.ZN(net3502)
);

OR2_X2 c3302(
.A1(net3484),
.A2(net3501),
.ZN(net3503)
);

DFFRS_X1 c3303(
.D(net3405),
.RN(net3487),
.SN(net3470),
.CK(clk),
.Q(net3505),
.QN(net3504)
);

NOR2_X4 c3304(
.A1(net3472),
.A2(net10984),
.ZN(net3506)
);

NOR3_X2 c3305(
.A1(net3489),
.A2(net3484),
.A3(net3264),
.ZN(net3507)
);

NOR2_X2 c3306(
.A1(net2379),
.A2(net3477),
.ZN(net3508)
);

INV_X8 c3307(
.A(net11302),
.ZN(net3509)
);

AOI222_X1 c3308(
.A1(net3487),
.A2(net3414),
.B1(net3508),
.B2(net3471),
.C1(net3373),
.C2(net2153),
.ZN(net3510)
);

AND3_X4 c3309(
.A1(net3473),
.A2(net3485),
.A3(net2469),
.ZN(net3511)
);

NAND3_X2 c3310(
.A1(net3501),
.A2(net3449),
.A3(net3509),
.ZN(net3512)
);

OR3_X1 c3311(
.A1(net3506),
.A2(net2379),
.A3(net11519),
.ZN(net3513)
);

XOR2_X2 c3312(
.A(net3463),
.B(net3488),
.Z(net3514)
);

NAND4_X2 c3313(
.A1(net3494),
.A2(net3373),
.A3(net3512),
.A4(net3509),
.ZN(net3515)
);

MUX2_X1 c3314(
.A(net3504),
.B(net3498),
.S(net11295),
.Z(net3516)
);

INV_X16 c3315(
.A(net10098),
.ZN(net3517)
);

OAI21_X4 c3316(
.A(net3517),
.B1(net3501),
.B2(net11522),
.ZN(net3518)
);

AOI222_X4 c3317(
.A1(net3513),
.A2(net3512),
.B1(net3516),
.B2(net1353),
.C1(net3418),
.C2(net3470),
.ZN(net3519)
);

MUX2_X2 c3318(
.A(net3471),
.B(net3464),
.S(net10726),
.Z(net3520)
);

NAND3_X4 c3319(
.A1(net2440),
.A2(net2438),
.A3(net3517),
.ZN(net3521)
);

INV_X32 c3320(
.A(net9645),
.ZN(net3522)
);

INV_X4 c3321(
.A(net2601),
.ZN(net3523)
);

XNOR2_X1 c3322(
.A(net2609),
.B(net2380),
.ZN(net3524)
);

INV_X1 c3323(
.A(net2533),
.ZN(net3525)
);

OR2_X4 c3324(
.A1(net2333),
.A2(net3516),
.ZN(net3526)
);

OR2_X1 c3325(
.A1(net2523),
.A2(net3373),
.ZN(net3527)
);

INV_X2 c3326(
.A(net2603),
.ZN(net3528)
);

INV_X8 c3327(
.A(net11346),
.ZN(net3529)
);

INV_X16 c3328(
.A(net626),
.ZN(net3530)
);

INV_X32 c3329(
.A(net10079),
.ZN(net3531)
);

XNOR2_X2 c3330(
.A(net2456),
.B(net2377),
.ZN(net3532)
);

INV_X4 c3331(
.A(net10025),
.ZN(net3533)
);

INV_X1 c3332(
.A(net2569),
.ZN(net3534)
);

INV_X2 c3333(
.A(net3532),
.ZN(net3535)
);

DFFR_X2 c3334(
.D(net2602),
.RN(net3373),
.CK(clk),
.Q(net3537),
.QN(net3536)
);

AND2_X4 c3335(
.A1(net3469),
.A2(net2601),
.ZN(net3538)
);

INV_X8 c3336(
.A(net3523),
.ZN(net3539)
);

INV_X16 c3337(
.A(net3539),
.ZN(net3540)
);

AND2_X1 c3338(
.A1(net3538),
.A2(net3471),
.ZN(net3541)
);

NAND2_X1 c3339(
.A1(net2153),
.A2(net1607),
.ZN(net3542)
);

INV_X32 c3340(
.A(net9890),
.ZN(net3543)
);

OR3_X4 c3341(
.A1(net3522),
.A2(net3530),
.A3(net3527),
.ZN(net3544)
);

INV_X4 c3342(
.A(net3508),
.ZN(net3545)
);

NAND2_X2 c3343(
.A1(net3464),
.A2(net3509),
.ZN(net3546)
);

DFFRS_X2 c3344(
.D(net2610),
.RN(net2455),
.SN(net3340),
.CK(clk),
.Q(net3548),
.QN(net3547)
);

NAND2_X4 c3345(
.A1(net3537),
.A2(net3543),
.ZN(net3549)
);

INV_X1 c3346(
.A(net9890),
.ZN(net3550)
);

AND2_X2 c3347(
.A1(net3530),
.A2(net3472),
.ZN(net3551)
);

AND3_X2 c3348(
.A1(net2614),
.A2(net3530),
.A3(net2532),
.ZN(net3552)
);

XOR2_X1 c3349(
.A(net3449),
.B(net3536),
.Z(net3553)
);

INV_X2 c3350(
.A(net3546),
.ZN(net3554)
);

INV_X8 c3351(
.A(net9957),
.ZN(net3555)
);

NOR2_X1 c3352(
.A1(net2590),
.A2(net2609),
.ZN(net3556)
);

OR2_X2 c3353(
.A1(net1607),
.A2(net3554),
.ZN(net3557)
);

INV_X16 c3354(
.A(net10124),
.ZN(net3558)
);

INV_X32 c3355(
.A(net2586),
.ZN(net3559)
);

INV_X4 c3356(
.A(net3556),
.ZN(net3560)
);

INV_X1 c3357(
.A(net10283),
.ZN(net3561)
);

NOR2_X4 c3358(
.A1(net3559),
.A2(net3472),
.ZN(net3562)
);

NOR2_X2 c3359(
.A1(net3550),
.A2(net3561),
.ZN(net3563)
);

INV_X2 c3360(
.A(net3505),
.ZN(net3564)
);

XOR2_X2 c3361(
.A(net1403),
.B(net3535),
.Z(net3565)
);

XNOR2_X1 c3362(
.A(net2597),
.B(net3561),
.ZN(net3566)
);

OR2_X4 c3363(
.A1(net3554),
.A2(net3435),
.ZN(net3567)
);

OR2_X1 c3364(
.A1(net3552),
.A2(net3564),
.ZN(net3568)
);

XNOR2_X2 c3365(
.A(net3525),
.B(net3557),
.ZN(net3569)
);

AND2_X4 c3366(
.A1(net3560),
.A2(net3527),
.ZN(net3570)
);

INV_X8 c3367(
.A(net3561),
.ZN(net3571)
);

AND2_X1 c3368(
.A1(net3533),
.A2(net2557),
.ZN(net3572)
);

OAI33_X1 c3369(
.A1(net3431),
.A2(net3564),
.A3(net2629),
.B1(net3453),
.B2(net2557),
.B3(net1513),
.ZN(net3573)
);

INV_X16 c3370(
.A(net11449),
.ZN(net3574)
);

NOR3_X1 c3371(
.A1(net3537),
.A2(net1637),
.A3(net3561),
.ZN(net3575)
);

INV_X32 c3372(
.A(net11441),
.ZN(net3576)
);

NAND2_X1 c3373(
.A1(net3570),
.A2(net3561),
.ZN(net3577)
);

INV_X4 c3374(
.A(net10145),
.ZN(net3578)
);

INV_X1 c3375(
.A(net3553),
.ZN(net3579)
);

INV_X2 c3376(
.A(net3562),
.ZN(net3580)
);

AOI221_X2 c3377(
.A(net1504),
.B1(net3564),
.B2(net3574),
.C1(net2589),
.C2(net2629),
.ZN(net3581)
);

OR3_X2 c3378(
.A1(net3527),
.A2(net3580),
.A3(net2928),
.ZN(net3582)
);

OAI21_X2 c3379(
.A(net2459),
.B1(net3452),
.B2(net3580),
.ZN(net3583)
);

NAND2_X2 c3380(
.A1(net3578),
.A2(net3561),
.ZN(net3584)
);

NAND2_X4 c3381(
.A1(net3558),
.A2(net3564),
.ZN(net3585)
);

OAI21_X1 c3382(
.A(net3472),
.B1(net3568),
.B2(net3564),
.ZN(net3586)
);

INV_X8 c3383(
.A(net11296),
.ZN(net3587)
);

AND2_X2 c3384(
.A1(net3442),
.A2(net2601),
.ZN(net3588)
);

XOR2_X1 c3385(
.A(net3581),
.B(net3580),
.Z(net3589)
);

NOR2_X1 c3386(
.A1(net3564),
.A2(net3578),
.ZN(net3590)
);

AOI21_X2 c3387(
.A(net3574),
.B1(net3544),
.B2(net2532),
.ZN(net3591)
);

OR2_X2 c3388(
.A1(net3587),
.A2(net3523),
.ZN(net3592)
);

AOI21_X1 c3389(
.A(net3576),
.B1(net3545),
.B2(net3554),
.ZN(net3593)
);

INV_X16 c3390(
.A(net9645),
.ZN(net3594)
);

NOR2_X4 c3391(
.A1(net3584),
.A2(net3594),
.ZN(net3595)
);

NOR2_X2 c3392(
.A1(net3557),
.A2(net3584),
.ZN(net3596)
);

AOI21_X4 c3393(
.A(net3566),
.B1(net3595),
.B2(net3596),
.ZN(net3597)
);

XOR2_X2 c3394(
.A(net3589),
.B(net3596),
.Z(net3598)
);

AND3_X1 c3395(
.A1(net3579),
.A2(net3580),
.A3(net3594),
.ZN(net3599)
);

SDFF_X1 c3396(
.D(net3580),
.SE(net3577),
.SI(net3599),
.CK(clk),
.Q(net3601),
.QN(net3600)
);

XNOR2_X1 c3397(
.A(net3591),
.B(net10506),
.ZN(net3602)
);

NAND3_X1 c3398(
.A1(net2632),
.A2(net1309),
.A3(net3600),
.ZN(net3603)
);

NOR3_X4 c3399(
.A1(net3603),
.A2(net3595),
.A3(net3580),
.ZN(net3604)
);

NOR3_X2 c3400(
.A1(net2530),
.A2(net3590),
.A3(net3604),
.ZN(net3605)
);

OR2_X4 c3401(
.A1(net3601),
.A2(net10507),
.ZN(net3606)
);

AND3_X4 c3402(
.A1(net3606),
.A2(net3594),
.A3(net10875),
.ZN(net3607)
);

OR2_X1 c3403(
.A1(net2649),
.A2(net696),
.ZN(net3608)
);

XNOR2_X2 c3404(
.A(net3529),
.B(net3575),
.ZN(net3609)
);

AND2_X4 c3405(
.A1(net1353),
.A2(net2621),
.ZN(net3610)
);

AND2_X1 c3406(
.A1(net1609),
.A2(net2589),
.ZN(net3611)
);

NAND2_X1 c3407(
.A1(net507),
.A2(net3568),
.ZN(net3612)
);

INV_X32 c3408(
.A(net11133),
.ZN(net3613)
);

INV_X4 c3409(
.A(net10947),
.ZN(net3614)
);

INV_X1 c3410(
.A(net3534),
.ZN(net3615)
);

INV_X2 c3411(
.A(net3492),
.ZN(net3616)
);

DFFS_X1 c3412(
.D(net3498),
.SN(net2605),
.CK(clk),
.Q(net3618),
.QN(net3617)
);

INV_X8 c3413(
.A(net11133),
.ZN(net3619)
);

INV_X16 c3414(
.A(net3597),
.ZN(net3620)
);

NAND2_X2 c3415(
.A1(net3540),
.A2(net2649),
.ZN(net3621)
);

NAND2_X4 c3416(
.A1(net3599),
.A2(net3544),
.ZN(net3622)
);

INV_X32 c3417(
.A(net3441),
.ZN(net3623)
);

NAND3_X2 c3418(
.A1(net3354),
.A2(net3565),
.A3(net2649),
.ZN(net3624)
);

INV_X4 c3419(
.A(net10297),
.ZN(net3625)
);

AND2_X2 c3420(
.A1(net3551),
.A2(net3592),
.ZN(net3626)
);

INV_X1 c3421(
.A(net11359),
.ZN(net3627)
);

INV_X2 c3422(
.A(net3535),
.ZN(net3628)
);

XOR2_X1 c3423(
.A(net3618),
.B(net3535),
.Z(net3629)
);

SDFF_X2 c3424(
.D(net1525),
.SE(net3498),
.SI(net654),
.CK(clk),
.Q(net3631),
.QN(net3630)
);

NOR2_X1 c3425(
.A1(net3493),
.A2(net3630),
.ZN(net3632)
);

OR2_X2 c3426(
.A1(net2483),
.A2(net2713),
.ZN(net3633)
);

NOR2_X4 c3427(
.A1(net758),
.A2(net2589),
.ZN(net3634)
);

NOR2_X2 c3428(
.A1(net3592),
.A2(net3599),
.ZN(net3635)
);

XOR2_X2 c3429(
.A(net1645),
.B(net3498),
.Z(net3636)
);

XNOR2_X1 c3430(
.A(net2621),
.B(net3626),
.ZN(net3637)
);

INV_X8 c3431(
.A(net11134),
.ZN(net3638)
);

OR3_X1 c3432(
.A1(net3624),
.A2(net3634),
.A3(net1729),
.ZN(net3639)
);

OR2_X4 c3433(
.A1(net3531),
.A2(net2557),
.ZN(net3640)
);

OR2_X1 c3434(
.A1(net2336),
.A2(net3631),
.ZN(net3641)
);

INV_X16 c3435(
.A(net11298),
.ZN(net3642)
);

INV_X32 c3436(
.A(net11152),
.ZN(net3643)
);

XNOR2_X2 c3437(
.A(net3636),
.B(net2621),
.ZN(net3644)
);

INV_X4 c3438(
.A(net3623),
.ZN(net3645)
);

AND2_X4 c3439(
.A1(net1522),
.A2(net3627),
.ZN(net3646)
);

INV_X1 c3440(
.A(net10366),
.ZN(net3647)
);

AND2_X1 c3441(
.A1(net3614),
.A2(net2649),
.ZN(net3648)
);

INV_X2 c3442(
.A(net11003),
.ZN(net3649)
);

NAND2_X1 c3443(
.A1(net3628),
.A2(net2661),
.ZN(net3650)
);

NAND2_X2 c3444(
.A1(net3632),
.A2(net3637),
.ZN(net3651)
);

INV_X8 c3445(
.A(net9928),
.ZN(net3652)
);

NAND2_X4 c3446(
.A1(net2676),
.A2(net3633),
.ZN(net3653)
);

INV_X16 c3447(
.A(net11255),
.ZN(net3654)
);

MUX2_X1 c3448(
.A(net3647),
.B(net2153),
.S(net3638),
.Z(net3655)
);

AND2_X2 c3449(
.A1(net3625),
.A2(net3644),
.ZN(net3656)
);

XOR2_X1 c3450(
.A(net3613),
.B(net3544),
.Z(net3657)
);

NOR2_X1 c3451(
.A1(net3645),
.A2(net11174),
.ZN(net3658)
);

INV_X32 c3452(
.A(net11465),
.ZN(net3659)
);

OR2_X2 c3453(
.A1(net3650),
.A2(net11174),
.ZN(net3660)
);

NOR2_X4 c3454(
.A1(net3575),
.A2(net3610),
.ZN(net3661)
);

NOR2_X2 c3455(
.A1(net3638),
.A2(net3658),
.ZN(net3662)
);

XOR2_X2 c3456(
.A(net3568),
.B(net2634),
.Z(net3663)
);

XNOR2_X1 c3457(
.A(net2368),
.B(net3612),
.ZN(net3664)
);

OR2_X4 c3458(
.A1(net3630),
.A2(net11117),
.ZN(net3665)
);

OAI21_X4 c3459(
.A(net3549),
.B1(net3665),
.B2(net3638),
.ZN(net3666)
);

OR2_X1 c3460(
.A1(net3655),
.A2(net3535),
.ZN(net3667)
);

XNOR2_X2 c3461(
.A(net3658),
.B(net3629),
.ZN(net3668)
);

AND2_X4 c3462(
.A1(net3659),
.A2(net3629),
.ZN(net3669)
);

AND2_X1 c3463(
.A1(net3609),
.A2(net3669),
.ZN(net3670)
);

NAND2_X1 c3464(
.A1(net3573),
.A2(net3670),
.ZN(net3671)
);

MUX2_X2 c3465(
.A(net3657),
.B(net2704),
.S(net3666),
.Z(net3672)
);

AOI222_X2 c3466(
.A1(net3641),
.A2(net3524),
.B1(net3612),
.B2(net3666),
.C1(net2649),
.C2(net3615),
.ZN(net3673)
);

AOI221_X1 c3467(
.A(net3672),
.B1(net1701),
.B2(net3634),
.C1(net3632),
.C2(net3666),
.ZN(net3674)
);

NAND2_X2 c3468(
.A1(net3643),
.A2(net1687),
.ZN(net3675)
);

INV_X4 c3469(
.A(net11152),
.ZN(net3676)
);

INV_X1 c3470(
.A(net11062),
.ZN(net3677)
);

NAND3_X4 c3471(
.A1(net3372),
.A2(net3668),
.A3(net3617),
.ZN(net3678)
);

INV_X2 c3472(
.A(net10010),
.ZN(net3679)
);

NAND2_X4 c3473(
.A1(net3679),
.A2(net694),
.ZN(net3680)
);

AND2_X2 c3474(
.A1(net3680),
.A2(net11150),
.ZN(net3681)
);

XOR2_X1 c3475(
.A(net3596),
.B(net3615),
.Z(net3682)
);

NOR2_X1 c3476(
.A1(net3658),
.A2(net11150),
.ZN(net3683)
);

OR2_X2 c3477(
.A1(net2657),
.A2(net3683),
.ZN(net3684)
);

OR3_X4 c3478(
.A1(net3684),
.A2(net3632),
.A3(net3670),
.ZN(net3685)
);

AND3_X2 c3479(
.A1(net3684),
.A2(net3618),
.A3(net11117),
.ZN(net3686)
);

OAI221_X1 c3480(
.A(net3683),
.B1(net3597),
.B2(net3666),
.C1(net3615),
.C2(net1599),
.ZN(net3687)
);

NOR2_X4 c3481(
.A1(net3682),
.A2(net3610),
.ZN(net3688)
);

NOR2_X2 c3482(
.A1(net3678),
.A2(net3682),
.ZN(net3689)
);

XOR2_X2 c3483(
.A(net2514),
.B(net3678),
.Z(net3690)
);

SDFFRS_X1 c3484(
.D(net3689),
.RN(net3678),
.SE(net3684),
.SI(net3451),
.SN(net3666),
.CK(clk),
.Q(net3692),
.QN(net3691)
);

OR4_X4 c3485(
.A1(net2663),
.A2(net3684),
.A3(net3692),
.A4(net3666),
.ZN(net3693)
);

INV_X8 c3486(
.A(net843),
.ZN(net3694)
);

INV_X16 c3487(
.A(net11188),
.ZN(net3695)
);

XNOR2_X1 c3488(
.A(net2768),
.B(net2749),
.ZN(net3696)
);

INV_X32 c3489(
.A(net11525),
.ZN(net3697)
);

OR2_X4 c3490(
.A1(net2744),
.A2(net2806),
.ZN(net3698)
);

OR2_X1 c3491(
.A1(net496),
.A2(net2781),
.ZN(net3699)
);

INV_X4 c3492(
.A(net9646),
.ZN(net3700)
);

XNOR2_X2 c3493(
.A(net3633),
.B(net2805),
.ZN(net3701)
);

AND2_X4 c3494(
.A1(net1782),
.A2(net774),
.ZN(net3702)
);

INV_X1 c3495(
.A(net11317),
.ZN(net3703)
);

NOR3_X1 c3496(
.A1(net1675),
.A2(net3675),
.A3(net3666),
.ZN(net3704)
);

AND2_X1 c3497(
.A1(net2732),
.A2(net3704),
.ZN(net3705)
);

INV_X2 c3498(
.A(net10547),
.ZN(net3706)
);

NAND2_X1 c3499(
.A1(net2750),
.A2(net3542),
.ZN(net3707)
);

INV_X8 c3500(
.A(net1691),
.ZN(net3708)
);

OAI22_X2 c3501(
.A1(net789),
.A2(net2716),
.B1(net3704),
.B2(net11030),
.ZN(net3709)
);

INV_X16 c3502(
.A(net2795),
.ZN(net3710)
);

OR3_X2 c3503(
.A1(net2801),
.A2(net3708),
.A3(net2754),
.ZN(net3711)
);

INV_X32 c3504(
.A(net9647),
.ZN(net3712)
);

OAI21_X2 c3505(
.A(net467),
.B1(net3541),
.B2(net2754),
.ZN(net3713)
);

DFFRS_X1 c3506(
.D(net3642),
.RN(net2801),
.SN(net3708),
.CK(clk),
.Q(net3715),
.QN(net3714)
);

NAND2_X2 c3507(
.A1(net3703),
.A2(net3629),
.ZN(net3716)
);

OAI211_X4 c3508(
.A(net3694),
.B(net2725),
.C1(net3714),
.C2(net3666),
.ZN(net3717)
);

OAI21_X1 c3509(
.A(net2753),
.B1(net3695),
.B2(net10529),
.ZN(net3718)
);

NAND2_X4 c3510(
.A1(net3373),
.A2(net1743),
.ZN(net3719)
);

AND2_X2 c3511(
.A1(net3631),
.A2(net840),
.ZN(net3720)
);

INV_X4 c3512(
.A(net11364),
.ZN(net3721)
);

AOI21_X2 c3513(
.A(net1782),
.B1(net3712),
.B2(net11251),
.ZN(net3722)
);

INV_X1 c3514(
.A(net10484),
.ZN(net3723)
);

XOR2_X1 c3515(
.A(net2805),
.B(net2765),
.Z(net3724)
);

INV_X2 c3516(
.A(net10423),
.ZN(net3725)
);

NOR2_X1 c3517(
.A1(net2709),
.A2(net3708),
.ZN(net3726)
);

OR2_X2 c3518(
.A1(net3706),
.A2(net839),
.ZN(net3727)
);

NOR2_X4 c3519(
.A1(net1686),
.A2(net3725),
.ZN(net3728)
);

NOR2_X2 c3520(
.A1(net3712),
.A2(net3725),
.ZN(net3729)
);

XOR2_X2 c3521(
.A(net3720),
.B(net1791),
.Z(net3730)
);

INV_X8 c3522(
.A(net3722),
.ZN(net3731)
);

XNOR2_X1 c3523(
.A(net3731),
.B(net3723),
.ZN(net3732)
);

OR2_X4 c3524(
.A1(net3565),
.A2(net3704),
.ZN(net3733)
);

OR2_X1 c3525(
.A1(net2684),
.A2(net3731),
.ZN(net3734)
);

AOI21_X1 c3526(
.A(net1776),
.B1(net2768),
.B2(net11268),
.ZN(net3735)
);

XNOR2_X2 c3527(
.A(net2765),
.B(net2716),
.ZN(net3736)
);

AND2_X4 c3528(
.A1(net2747),
.A2(net3727),
.ZN(net3737)
);

AOI21_X4 c3529(
.A(net3732),
.B1(net3721),
.B2(net3718),
.ZN(net3738)
);

INV_X16 c3530(
.A(net11052),
.ZN(net3739)
);

AND2_X1 c3531(
.A1(net3696),
.A2(net2716),
.ZN(net3740)
);

AND3_X1 c3532(
.A1(net2733),
.A2(net3732),
.A3(net3708),
.ZN(net3741)
);

NAND2_X1 c3533(
.A1(net3738),
.A2(net3697),
.ZN(net3742)
);

NAND2_X2 c3534(
.A1(net3725),
.A2(net11524),
.ZN(net3743)
);

NAND2_X4 c3535(
.A1(net835),
.A2(net2799),
.ZN(net3744)
);

AND2_X2 c3536(
.A1(net3730),
.A2(net3615),
.ZN(net3745)
);

INV_X32 c3537(
.A(net11350),
.ZN(net3746)
);

XOR2_X1 c3538(
.A(net3705),
.B(net3732),
.Z(net3747)
);

INV_X4 c3539(
.A(net10451),
.ZN(net3748)
);

DFFS_X2 c3540(
.D(net3709),
.SN(net3732),
.CK(clk),
.Q(net3750),
.QN(net3749)
);

NOR2_X1 c3541(
.A1(net3744),
.A2(net2461),
.ZN(net3751)
);

OR2_X2 c3542(
.A1(net3716),
.A2(net3727),
.ZN(net3752)
);

NOR2_X4 c3543(
.A1(net3726),
.A2(net1675),
.ZN(net3753)
);

NAND3_X1 c3544(
.A1(net3734),
.A2(net3735),
.A3(net2605),
.ZN(net3754)
);

OAI222_X1 c3545(
.A1(net3743),
.A2(net3734),
.B1(net694),
.B2(net2709),
.C1(net3733),
.C2(net3723),
.ZN(net3755)
);

NOR2_X2 c3546(
.A1(net3753),
.A2(net3751),
.ZN(net3756)
);

DFFR_X1 c3547(
.D(net3719),
.RN(net2605),
.CK(clk),
.Q(net3758),
.QN(net3757)
);

XOR2_X2 c3548(
.A(net3713),
.B(net3712),
.Z(net3759)
);

NOR3_X4 c3549(
.A1(net3748),
.A2(net3757),
.A3(net3735),
.ZN(net3760)
);

XNOR2_X1 c3550(
.A(net3756),
.B(net2461),
.ZN(net3761)
);

OAI222_X4 c3551(
.A1(net3717),
.A2(net3756),
.B1(net3732),
.B2(net3742),
.C1(net3749),
.C2(net11525),
.ZN(net3762)
);

OR2_X4 c3552(
.A1(net3733),
.A2(net3717),
.ZN(net3763)
);

NOR3_X2 c3553(
.A1(net746),
.A2(net2535),
.A3(net3745),
.ZN(net3764)
);

INV_X1 c3554(
.A(net3708),
.ZN(net3765)
);

OAI221_X4 c3555(
.A(net2720),
.B1(net3759),
.B2(net3738),
.C1(net3723),
.C2(net1743),
.ZN(net3766)
);

DFFRS_X2 c3556(
.D(net3763),
.RN(net3709),
.SN(net3496),
.CK(clk),
.Q(net3768),
.QN(net3767)
);

OR2_X1 c3557(
.A1(net3629),
.A2(net3725),
.ZN(net3769)
);

AND3_X4 c3558(
.A1(net3758),
.A2(net3722),
.A3(net10854),
.ZN(net3770)
);

OAI211_X1 c3559(
.A(net3761),
.B(net3733),
.C1(net3724),
.C2(net3767),
.ZN(net3771)
);

OAI221_X2 c3560(
.A(net2771),
.B1(net3749),
.B2(net2754),
.C1(net3723),
.C2(net11356),
.ZN(net3772)
);

NAND3_X2 c3561(
.A1(net3769),
.A2(net1732),
.A3(net2716),
.ZN(net3773)
);

INV_X2 c3562(
.A(net10338),
.ZN(net3774)
);

AOI221_X4 c3563(
.A(net3700),
.B1(net3731),
.B2(net3774),
.C1(net3723),
.C2(net1686),
.ZN(net3775)
);

OR3_X1 c3564(
.A1(net1643),
.A2(net3768),
.A3(net1806),
.ZN(net3776)
);

MUX2_X1 c3565(
.A(net3772),
.B(net3774),
.S(net11339),
.Z(net3777)
);

SDFFR_X1 c3566(
.D(net3735),
.RN(net2508),
.SE(net2724),
.SI(net3714),
.CK(clk),
.Q(net3779),
.QN(net3778)
);

NOR4_X4 c3567(
.A1(net3777),
.A2(net3778),
.A3(net3704),
.A4(net11339),
.ZN(net3780)
);

AOI221_X2 c3568(
.A(net3724),
.B1(net3779),
.B2(net2799),
.C1(net3774),
.C2(net11118),
.ZN(net3781)
);

NOR4_X2 c3569(
.A1(net3542),
.A2(net1892),
.A3(net3666),
.A4(net1857),
.ZN(net3782)
);

XNOR2_X2 c3570(
.A(net907),
.B(net3669),
.ZN(net3783)
);

AND2_X4 c3571(
.A1(net1893),
.A2(net774),
.ZN(net3784)
);

AND2_X1 c3572(
.A1(net1874),
.A2(net2891),
.ZN(net3785)
);

NAND2_X1 c3573(
.A1(net2853),
.A2(net2849),
.ZN(net3786)
);

INV_X8 c3574(
.A(net9658),
.ZN(net3787)
);

NAND2_X2 c3575(
.A1(net2891),
.A2(net1802),
.ZN(net3788)
);

INV_X16 c3576(
.A(net9804),
.ZN(net3789)
);

OAI21_X4 c3577(
.A(net877),
.B1(net2773),
.B2(net1870),
.ZN(net3790)
);

DFFR_X2 c3578(
.D(net2809),
.RN(net3704),
.CK(clk),
.Q(net3792),
.QN(net3791)
);

NAND2_X4 c3579(
.A1(net1824),
.A2(net2854),
.ZN(net3793)
);

AND2_X2 c3580(
.A1(net2811),
.A2(net3715),
.ZN(net3794)
);

XOR2_X1 c3581(
.A(net917),
.B(net11466),
.Z(net3795)
);

MUX2_X2 c3582(
.A(net3715),
.B(net3794),
.S(net3791),
.Z(net3796)
);

NOR2_X1 c3583(
.A1(net2807),
.A2(net11113),
.ZN(net3797)
);

OR2_X2 c3584(
.A1(net3797),
.A2(net3692),
.ZN(net3798)
);

NOR2_X4 c3585(
.A1(net2874),
.A2(net2753),
.ZN(net3799)
);

NOR2_X2 c3586(
.A1(net1828),
.A2(net1802),
.ZN(net3800)
);

SDFF_X1 c3587(
.D(net914),
.SE(net2749),
.SI(net2849),
.CK(clk),
.Q(net3802),
.QN(net3801)
);

XOR2_X2 c3588(
.A(net3784),
.B(net1870),
.Z(net3803)
);

NAND3_X4 c3589(
.A1(net2840),
.A2(net1802),
.A3(net2862),
.ZN(net3804)
);

XNOR2_X1 c3590(
.A(net1635),
.B(net10882),
.ZN(net3805)
);

INV_X32 c3591(
.A(net10298),
.ZN(net3806)
);

DFFS_X1 c3592(
.D(net2896),
.SN(net3798),
.CK(clk),
.Q(net3808),
.QN(net3807)
);

OR2_X4 c3593(
.A1(net2879),
.A2(net3698),
.ZN(net3809)
);

OR3_X4 c3594(
.A1(net3782),
.A2(net2860),
.A3(net1893),
.ZN(net3810)
);

OR2_X1 c3595(
.A1(net3699),
.A2(net2719),
.ZN(net3811)
);

XNOR2_X2 c3596(
.A(net1886),
.B(net3799),
.ZN(net3812)
);

AND2_X4 c3597(
.A1(net3787),
.A2(net10794),
.ZN(net3813)
);

AND2_X1 c3598(
.A1(net2836),
.A2(net1851),
.ZN(net3814)
);

AND3_X2 c3599(
.A1(net3812),
.A2(net3782),
.A3(net877),
.ZN(net3815)
);

NOR3_X1 c3600(
.A1(net3813),
.A2(net3812),
.A3(net2848),
.ZN(net3816)
);

NAND2_X1 c3601(
.A1(net2833),
.A2(net2862),
.ZN(net3817)
);

NAND2_X2 c3602(
.A1(net2781),
.A2(net1881),
.ZN(net3818)
);

OR3_X2 c3603(
.A1(net1858),
.A2(net2754),
.A3(net10674),
.ZN(net3819)
);

NAND2_X4 c3604(
.A1(net3616),
.A2(net2593),
.ZN(net3820)
);

INV_X4 c3605(
.A(net10375),
.ZN(net3821)
);

AND2_X2 c3606(
.A1(net2753),
.A2(net3788),
.ZN(net3822)
);

XOR2_X1 c3607(
.A(net2754),
.B(net879),
.Z(net3823)
);

SDFF_X2 c3608(
.D(net3815),
.SE(net3785),
.SI(net3542),
.CK(clk),
.Q(net3825),
.QN(net3824)
);

NOR2_X1 c3609(
.A1(net3787),
.A2(net3803),
.ZN(net3826)
);

OAI21_X2 c3610(
.A(net3806),
.B1(net3812),
.B2(net889),
.ZN(net3827)
);

DFFRS_X1 c3611(
.D(net3792),
.RN(net2809),
.SN(net2749),
.CK(clk),
.Q(net3829),
.QN(net3828)
);

OR2_X2 c3612(
.A1(net3811),
.A2(net11113),
.ZN(net3830)
);

OAI21_X1 c3613(
.A(net3695),
.B1(net3812),
.B2(net3820),
.ZN(net3831)
);

AOI21_X2 c3614(
.A(net3822),
.B1(net3824),
.B2(net2839),
.ZN(net3832)
);

NOR2_X4 c3615(
.A1(net2883),
.A2(net11466),
.ZN(net3833)
);

INV_X1 c3616(
.A(net10266),
.ZN(net3834)
);

NOR2_X2 c3617(
.A1(net3739),
.A2(net2860),
.ZN(net3835)
);

AOI21_X1 c3618(
.A(net2839),
.B1(net2819),
.B2(net3812),
.ZN(net3836)
);

AOI21_X4 c3619(
.A(net2833),
.B1(net3807),
.B2(net10904),
.ZN(net3837)
);

XOR2_X2 c3620(
.A(net1870),
.B(net2829),
.Z(net3838)
);

XNOR2_X1 c3621(
.A(net889),
.B(net3768),
.ZN(net3839)
);

OR2_X4 c3622(
.A1(net2820),
.A2(net3834),
.ZN(net3840)
);

OR2_X1 c3623(
.A1(net3805),
.A2(net3835),
.ZN(net3841)
);

AND3_X1 c3624(
.A1(net1865),
.A2(net3803),
.A3(net3801),
.ZN(net3842)
);

DFFS_X2 c3625(
.D(net3842),
.SN(net1851),
.CK(clk),
.Q(net3844),
.QN(net3843)
);

XNOR2_X2 c3626(
.A(net3704),
.B(net3834),
.ZN(net3845)
);

NAND3_X1 c3627(
.A1(net2749),
.A2(net3837),
.A3(net3834),
.ZN(net3846)
);

AND2_X4 c3628(
.A1(net1730),
.A2(net3845),
.ZN(net3847)
);

AND2_X1 c3629(
.A1(net1701),
.A2(net2853),
.ZN(net3848)
);

AOI211_X4 c3630(
.A(net3817),
.B(net3840),
.C1(net3829),
.C2(net3542),
.ZN(net3849)
);

DFFR_X1 c3631(
.D(net3831),
.RN(net3841),
.CK(clk),
.Q(net3851),
.QN(net3850)
);

NAND2_X1 c3632(
.A1(net774),
.A2(net2900),
.ZN(net3852)
);

OAI222_X2 c3633(
.A1(net1877),
.A2(net3852),
.B1(net3828),
.B2(net863),
.C1(net2848),
.C2(net2894),
.ZN(net3853)
);

SDFFR_X2 c3634(
.D(net3845),
.RN(net3835),
.SE(net3842),
.SI(net3704),
.CK(clk),
.Q(net3855),
.QN(net3854)
);

NOR4_X1 c3635(
.A1(net3827),
.A2(net3616),
.A3(net2719),
.A4(net3849),
.ZN(net3856)
);

SDFFS_X1 c3636(
.D(net3800),
.SE(net3854),
.SI(net3841),
.SN(net1824),
.CK(clk),
.Q(net3858),
.QN(net3857)
);

AOI211_X2 c3637(
.A(net2869),
.B(net3823),
.C1(net2844),
.C2(net1885),
.ZN(net3859)
);

NAND2_X2 c3638(
.A1(net3852),
.A2(net10950),
.ZN(net3860)
);

NOR3_X4 c3639(
.A1(net3795),
.A2(net3819),
.A3(net3835),
.ZN(net3861)
);

SDFFS_X2 c3640(
.D(net3845),
.SE(net3849),
.SI(net2849),
.SN(net10878),
.CK(clk),
.Q(net3863),
.QN(net3862)
);

INV_X2 c3641(
.A(net9657),
.ZN(net3864)
);

NOR3_X2 c3642(
.A1(net3783),
.A2(net2881),
.A3(net3811),
.ZN(net3865)
);

SDFFR_X1 c3643(
.D(net3847),
.RN(net3858),
.SE(net2861),
.SI(net3828),
.CK(clk),
.Q(net3867),
.QN(net3866)
);

AOI22_X1 c3644(
.A1(net2810),
.A2(net3838),
.B1(net3834),
.B2(net10877),
.ZN(net3868)
);

AND3_X4 c3645(
.A1(net3698),
.A2(net3848),
.A3(net3820),
.ZN(net3869)
);

SDFFR_X2 c3646(
.D(net3819),
.RN(net3839),
.SE(net3866),
.SI(net1870),
.CK(clk),
.Q(net3871),
.QN(net3870)
);

AND4_X4 c3647(
.A1(net3803),
.A2(net3863),
.A3(net3857),
.A4(net3670),
.ZN(net3872)
);

DFFRS_X2 c3648(
.D(net2857),
.RN(net3808),
.SN(net2873),
.CK(clk),
.Q(net3874),
.QN(net3873)
);

SDFF_X1 c3649(
.D(net3868),
.SE(net3872),
.SI(net3862),
.CK(clk),
.Q(net3876),
.QN(net3875)
);

NAND4_X1 c3650(
.A1(net3852),
.A2(net3867),
.A3(net3872),
.A4(net3834),
.ZN(net3877)
);

NAND3_X2 c3651(
.A1(net899),
.A2(net720),
.A3(net10995),
.ZN(net3878)
);

INV_X8 c3652(
.A(net9761),
.ZN(net3879)
);

INV_X16 c3653(
.A(net1000),
.ZN(net3880)
);

INV_X32 c3654(
.A(net9762),
.ZN(net3881)
);

INV_X4 c3655(
.A(net2906),
.ZN(net3882)
);

INV_X1 c3656(
.A(net1955),
.ZN(net3883)
);

DFFR_X2 c3657(
.D(net1011),
.RN(net2976),
.CK(clk),
.Q(net3885),
.QN(net3884)
);

NAND2_X4 c3658(
.A1(net3879),
.A2(net3880),
.ZN(net3886)
);

AND2_X2 c3659(
.A1(net1927),
.A2(net2926),
.ZN(net3887)
);

INV_X2 c3660(
.A(net2976),
.ZN(net3888)
);

INV_X8 c3661(
.A(net3882),
.ZN(net3889)
);

XOR2_X1 c3662(
.A(net3889),
.B(net1020),
.Z(net3890)
);

NOR2_X1 c3663(
.A1(net954),
.A2(net3889),
.ZN(net3891)
);

INV_X16 c3664(
.A(net2912),
.ZN(net3892)
);

OR2_X2 c3665(
.A1(net1986),
.A2(net2986),
.ZN(net3893)
);

INV_X32 c3666(
.A(net29),
.ZN(net3894)
);

INV_X4 c3667(
.A(net3879),
.ZN(net3895)
);

NOR2_X4 c3668(
.A1(net3886),
.A2(net3892),
.ZN(net3896)
);

INV_X1 c3669(
.A(net3894),
.ZN(net3897)
);

INV_X2 c3670(
.A(net3880),
.ZN(net3898)
);

NOR2_X2 c3671(
.A1(net2005),
.A2(net3886),
.ZN(net3899)
);

INV_X8 c3672(
.A(net9897),
.ZN(net3900)
);

INV_X16 c3673(
.A(net9898),
.ZN(net3901)
);

INV_X32 c3674(
.A(net991),
.ZN(net3902)
);

INV_X4 c3675(
.A(net3900),
.ZN(net3903)
);

XOR2_X2 c3676(
.A(net3898),
.B(net3892),
.Z(net3904)
);

DFFS_X1 c3677(
.D(net3896),
.SN(net3888),
.CK(clk),
.Q(net3906),
.QN(net3905)
);

XNOR2_X1 c3678(
.A(net3905),
.B(net2926),
.ZN(net3907)
);

INV_X1 c3679(
.A(net3895),
.ZN(net3908)
);

INV_X2 c3680(
.A(net1956),
.ZN(net3909)
);

DFFS_X2 c3681(
.D(net2990),
.SN(net3895),
.CK(clk),
.Q(net3911),
.QN(net3910)
);

OR2_X4 c3682(
.A1(net3907),
.A2(net1989),
.ZN(net3912)
);

INV_X8 c3683(
.A(net9930),
.ZN(net3913)
);

INV_X16 c3684(
.A(net2954),
.ZN(net3914)
);

DFFR_X1 c3685(
.D(net3913),
.RN(net3904),
.CK(clk),
.Q(net3916),
.QN(net3915)
);

INV_X32 c3686(
.A(net1987),
.ZN(net3917)
);

DFFR_X2 c3687(
.D(net2908),
.RN(net3899),
.CK(clk),
.Q(net3919),
.QN(net3918)
);

INV_X4 c3688(
.A(net9943),
.ZN(net3920)
);

INV_X1 c3689(
.A(net3908),
.ZN(net3921)
);

DFFS_X1 c3690(
.D(net3889),
.SN(net3896),
.CK(clk),
.Q(net3923),
.QN(net3922)
);

INV_X2 c3691(
.A(net3923),
.ZN(net3924)
);

INV_X8 c3692(
.A(net3919),
.ZN(net3925)
);

INV_X16 c3693(
.A(net3925),
.ZN(net3926)
);

OR2_X1 c3694(
.A1(net942),
.A2(net3894),
.ZN(net3927)
);

INV_X32 c3695(
.A(net9942),
.ZN(net3928)
);

INV_X4 c3696(
.A(net3901),
.ZN(net3929)
);

INV_X1 c3697(
.A(net3903),
.ZN(net3930)
);

INV_X2 c3698(
.A(net10643),
.ZN(net3931)
);

XNOR2_X2 c3699(
.A(net1980),
.B(net3909),
.ZN(net3932)
);

AND2_X4 c3700(
.A1(net3929),
.A2(net2912),
.ZN(net3933)
);

INV_X8 c3701(
.A(net3923),
.ZN(net3934)
);

OR3_X1 c3702(
.A1(net2926),
.A2(net3918),
.A3(net3902),
.ZN(net3935)
);

AND2_X1 c3703(
.A1(net3894),
.A2(net3914),
.ZN(net3936)
);

SDFF_X2 c3704(
.D(net2966),
.SE(net3932),
.SI(net3908),
.CK(clk),
.Q(net3938),
.QN(net3937)
);

INV_X16 c3705(
.A(net3931),
.ZN(net3939)
);

INV_X32 c3706(
.A(net3927),
.ZN(net3940)
);

INV_X4 c3707(
.A(net3890),
.ZN(net3941)
);

NAND2_X1 c3708(
.A1(net3930),
.A2(net3926),
.ZN(net3942)
);

INV_X1 c3709(
.A(net10644),
.ZN(net3943)
);

AOI222_X1 c3710(
.A1(net3926),
.A2(net3929),
.B1(net3907),
.B2(net3913),
.C1(net3902),
.C2(net2912),
.ZN(net3944)
);

NAND2_X2 c3711(
.A1(net3926),
.A2(net3908),
.ZN(net3945)
);

AOI222_X4 c3712(
.A1(net3892),
.A2(net3925),
.B1(net3884),
.B2(net2926),
.C1(net3904),
.C2(net3902),
.ZN(net3946)
);

INV_X2 c3713(
.A(net3924),
.ZN(net3947)
);

NAND2_X4 c3714(
.A1(net3939),
.A2(net3917),
.ZN(net3948)
);

INV_X8 c3715(
.A(net9984),
.ZN(net3949)
);

INV_X16 c3716(
.A(net3945),
.ZN(net3950)
);

MUX2_X1 c3717(
.A(net3949),
.B(net3914),
.S(net3920),
.Z(net3951)
);

AND2_X2 c3718(
.A1(net3943),
.A2(net3922),
.ZN(net3952)
);

INV_X32 c3719(
.A(net9929),
.ZN(net3953)
);

XOR2_X1 c3720(
.A(net3944),
.B(net2926),
.Z(net3954)
);

NOR2_X1 c3721(
.A1(net3883),
.A2(net3930),
.ZN(net3955)
);

OR2_X2 c3722(
.A1(net2983),
.A2(net3904),
.ZN(net3956)
);

OAI21_X4 c3723(
.A(net3932),
.B1(net2954),
.B2(net2965),
.ZN(net3957)
);

NOR2_X4 c3724(
.A1(net3935),
.A2(net3920),
.ZN(net3958)
);

DFFS_X2 c3725(
.D(net3927),
.SN(net3940),
.CK(clk),
.Q(net3960),
.QN(net3959)
);

INV_X4 c3726(
.A(net3941),
.ZN(net3961)
);

INV_X1 c3727(
.A(net3938),
.ZN(net3962)
);

NOR2_X2 c3728(
.A1(net3894),
.A2(net10880),
.ZN(net3963)
);

MUX2_X2 c3729(
.A(net3947),
.B(net3921),
.S(net2942),
.Z(net3964)
);

XOR2_X2 c3730(
.A(net3951),
.B(net3954),
.Z(net3965)
);

XNOR2_X1 c3731(
.A(net3953),
.B(net3961),
.ZN(net3966)
);

NAND3_X4 c3732(
.A1(net3966),
.A2(net3944),
.A3(net3937),
.ZN(net3967)
);

OR2_X4 c3733(
.A1(net3958),
.A2(net10879),
.ZN(net3968)
);

OR2_X1 c3734(
.A1(net3965),
.A2(net3955),
.ZN(net3969)
);

INV_X2 c3735(
.A(net3061),
.ZN(net3970)
);

XNOR2_X2 c3736(
.A(net3085),
.B(net3940),
.ZN(net3971)
);

INV_X8 c3737(
.A(net2067),
.ZN(net3972)
);

AND2_X4 c3738(
.A1(net3064),
.A2(net2067),
.ZN(net3973)
);

INV_X16 c3739(
.A(net3028),
.ZN(net3974)
);

INV_X32 c3740(
.A(net10301),
.ZN(net3975)
);

OR3_X4 c3741(
.A1(net3059),
.A2(net2964),
.A3(net3063),
.ZN(net3976)
);

AND2_X1 c3742(
.A1(net2052),
.A2(net942),
.ZN(net3977)
);

AND3_X2 c3743(
.A1(net3952),
.A2(net3064),
.A3(net2052),
.ZN(net3978)
);

INV_X4 c3744(
.A(net3963),
.ZN(net3979)
);

INV_X1 c3745(
.A(net9730),
.ZN(net3980)
);

DFFR_X1 c3746(
.D(net3917),
.RN(net1936),
.CK(clk),
.Q(net3982),
.QN(net3981)
);

DFFR_X2 c3747(
.D(net3978),
.RN(net3043),
.CK(clk),
.Q(net3984),
.QN(net3983)
);

NAND2_X1 c3748(
.A1(net3031),
.A2(net3917),
.ZN(net3985)
);

NAND2_X2 c3749(
.A1(net3979),
.A2(net2987),
.ZN(net3986)
);

NAND2_X4 c3750(
.A1(net3928),
.A2(net2980),
.ZN(net3987)
);

AND2_X2 c3751(
.A1(net3972),
.A2(net3028),
.ZN(net3988)
);

INV_X2 c3752(
.A(net11527),
.ZN(net3989)
);

INV_X8 c3753(
.A(net10668),
.ZN(net3990)
);

INV_X16 c3754(
.A(net1118),
.ZN(net3991)
);

NOR3_X1 c3755(
.A1(net1113),
.A2(net2098),
.A3(net3031),
.ZN(net3992)
);

INV_X32 c3756(
.A(net11056),
.ZN(net3993)
);

OR3_X2 c3757(
.A1(net3984),
.A2(net3970),
.A3(net3967),
.ZN(net3994)
);

OAI21_X2 c3758(
.A(net3043),
.B1(net3060),
.B2(net3987),
.ZN(net3995)
);

INV_X4 c3759(
.A(net3958),
.ZN(net3996)
);

XOR2_X1 c3760(
.A(net3970),
.B(net10715),
.Z(net3997)
);

INV_X1 c3761(
.A(net3010),
.ZN(net3998)
);

NOR2_X1 c3762(
.A1(net2076),
.A2(net3987),
.ZN(net3999)
);

INV_X2 c3763(
.A(net3060),
.ZN(net4000)
);

INV_X8 c3764(
.A(net3961),
.ZN(net4001)
);

OR2_X2 c3765(
.A1(net3881),
.A2(net3982),
.ZN(net4002)
);

INV_X16 c3766(
.A(net2013),
.ZN(net4003)
);

INV_X32 c3767(
.A(net3996),
.ZN(net4004)
);

NOR2_X4 c3768(
.A1(net3994),
.A2(net11019),
.ZN(net4005)
);

OAI21_X1 c3769(
.A(net3017),
.B1(net3988),
.B2(net3060),
.ZN(net4006)
);

NOR2_X2 c3770(
.A1(net3995),
.A2(net4005),
.ZN(net4007)
);

XOR2_X2 c3771(
.A(net3998),
.B(net3958),
.Z(net4008)
);

INV_X4 c3772(
.A(net3993),
.ZN(net4009)
);

XNOR2_X1 c3773(
.A(net3047),
.B(net3060),
.ZN(net4010)
);

OR2_X4 c3774(
.A1(net4005),
.A2(net4010),
.ZN(net4011)
);

INV_X1 c3775(
.A(net4002),
.ZN(net4012)
);

OR2_X1 c3776(
.A1(net4009),
.A2(net3884),
.ZN(net4013)
);

INV_X2 c3777(
.A(net11472),
.ZN(net4014)
);

OR4_X1 c3778(
.A1(net4010),
.A2(net3948),
.A3(net2962),
.A4(net3967),
.ZN(net4015)
);

XNOR2_X2 c3779(
.A(net1021),
.B(net3995),
.ZN(net4016)
);

AOI21_X2 c3780(
.A(net1936),
.B1(net3882),
.B2(net1944),
.ZN(net4017)
);

INV_X8 c3781(
.A(net4013),
.ZN(net4018)
);

INV_X16 c3782(
.A(net4008),
.ZN(net4019)
);

DFFS_X1 c3783(
.D(net3978),
.SN(net3010),
.CK(clk),
.Q(net4021),
.QN(net4020)
);

INV_X32 c3784(
.A(net9729),
.ZN(net4022)
);

AND2_X4 c3785(
.A1(net2980),
.A2(net10763),
.ZN(net4023)
);

AND2_X1 c3786(
.A1(net78),
.A2(net4015),
.ZN(net4024)
);

INV_X4 c3787(
.A(net10416),
.ZN(net4025)
);

INV_X1 c3788(
.A(net3980),
.ZN(net4026)
);

INV_X2 c3789(
.A(net4025),
.ZN(net4027)
);

NAND2_X1 c3790(
.A1(net4012),
.A2(net4005),
.ZN(net4028)
);

SDFFS_X1 c3791(
.D(net1927),
.SE(net4023),
.SI(net3028),
.SN(net3981),
.CK(clk),
.Q(net4030),
.QN(net4029)
);

NAND2_X2 c3792(
.A1(net4022),
.A2(net10667),
.ZN(net4031)
);

AOI21_X1 c3793(
.A(net3009),
.B1(net4029),
.B2(net3010),
.ZN(net4032)
);

NAND2_X4 c3794(
.A1(net2906),
.A2(net3902),
.ZN(net4033)
);

AOI21_X4 c3795(
.A(net4016),
.B1(net4026),
.B2(net11526),
.ZN(net4034)
);

SDFFS_X2 c3796(
.D(net4023),
.SE(net4025),
.SI(net4015),
.SN(net3904),
.CK(clk),
.Q(net4036),
.QN(net4035)
);

INV_X8 c3797(
.A(net10501),
.ZN(net4037)
);

AND2_X2 c3798(
.A1(net3970),
.A2(net4005),
.ZN(net4038)
);

AND3_X1 c3799(
.A1(net3990),
.A2(net4021),
.A3(net3988),
.ZN(net4039)
);

XOR2_X1 c3800(
.A(net3991),
.B(net4002),
.Z(net4040)
);

OAI33_X1 c3801(
.A1(net4027),
.A2(net4002),
.A3(net3992),
.B1(net4000),
.B2(net2077),
.B3(net3084),
.ZN(net4041)
);

INV_X16 c3802(
.A(net10299),
.ZN(net4042)
);

NAND3_X1 c3803(
.A1(net4000),
.A2(net3058),
.A3(net10764),
.ZN(net4043)
);

DFFS_X2 c3804(
.D(net4007),
.SN(net4013),
.CK(clk),
.Q(net4045),
.QN(net4044)
);

NOR2_X1 c3805(
.A1(net4031),
.A2(net3983),
.ZN(net4046)
);

OR2_X2 c3806(
.A1(net4042),
.A2(net4035),
.ZN(net4047)
);

NOR2_X4 c3807(
.A1(net3027),
.A2(net3061),
.ZN(net4048)
);

NOR2_X2 c3808(
.A1(net4034),
.A2(net3975),
.ZN(net4049)
);

INV_X32 c3809(
.A(net10826),
.ZN(net4050)
);

XOR2_X2 c3810(
.A(net1000),
.B(net4000),
.Z(net4051)
);

XNOR2_X1 c3811(
.A(net4051),
.B(net3980),
.ZN(net4052)
);

NOR3_X4 c3812(
.A1(net4047),
.A2(net4045),
.A3(net4015),
.ZN(net4053)
);

NOR3_X2 c3813(
.A1(net4032),
.A2(net3961),
.A3(net4049),
.ZN(net4054)
);

AND3_X4 c3814(
.A1(net4037),
.A2(net4049),
.A3(net4053),
.ZN(net4055)
);

NAND3_X2 c3815(
.A1(net3079),
.A2(net4053),
.A3(net10693),
.ZN(net4056)
);

OR2_X4 c3816(
.A1(net3997),
.A2(net11102),
.ZN(net4057)
);

OR3_X1 c3817(
.A1(net4044),
.A2(net4020),
.A3(net11102),
.ZN(net4058)
);

INV_X4 c3818(
.A(net9896),
.ZN(net4059)
);

OR2_X1 c3819(
.A1(net3137),
.A2(net2161),
.ZN(net4060)
);

XNOR2_X2 c3820(
.A(net3080),
.B(net3161),
.ZN(net4061)
);

AND2_X4 c3821(
.A1(net1173),
.A2(net2153),
.ZN(net4062)
);

AND2_X1 c3822(
.A1(net3119),
.A2(net4053),
.ZN(net4063)
);

NAND2_X1 c3823(
.A1(net3063),
.A2(net11238),
.ZN(net4064)
);

NAND2_X2 c3824(
.A1(net1174),
.A2(net3084),
.ZN(net4065)
);

NAND2_X4 c3825(
.A1(net3136),
.A2(net1141),
.ZN(net4066)
);

INV_X1 c3826(
.A(net3962),
.ZN(net4067)
);

AND2_X2 c3827(
.A1(net1192),
.A2(net4044),
.ZN(net4068)
);

INV_X2 c3828(
.A(net4053),
.ZN(net4069)
);

XOR2_X1 c3829(
.A(net1141),
.B(net4014),
.Z(net4070)
);

NOR2_X1 c3830(
.A1(net4070),
.A2(net3004),
.ZN(net4071)
);

OR2_X2 c3831(
.A1(net2088),
.A2(net2144),
.ZN(net4072)
);

INV_X8 c3832(
.A(net10610),
.ZN(net4073)
);

INV_X16 c3833(
.A(net9740),
.ZN(net4074)
);

INV_X32 c3834(
.A(net4072),
.ZN(net4075)
);

INV_X4 c3835(
.A(net10256),
.ZN(net4076)
);

NOR2_X4 c3836(
.A1(net4046),
.A2(net4049),
.ZN(net4077)
);

INV_X1 c3837(
.A(net11417),
.ZN(net4078)
);

NOR2_X2 c3838(
.A1(net4015),
.A2(net3004),
.ZN(net4079)
);

XOR2_X2 c3839(
.A(net4064),
.B(net3950),
.Z(net4080)
);

INV_X2 c3840(
.A(net11176),
.ZN(net4081)
);

INV_X8 c3841(
.A(net9740),
.ZN(net4082)
);

XNOR2_X1 c3842(
.A(net1922),
.B(net10714),
.ZN(net4083)
);

DFFR_X1 c3843(
.D(net4045),
.RN(net4049),
.CK(clk),
.Q(net4085),
.QN(net4084)
);

INV_X16 c3844(
.A(net9910),
.ZN(net4086)
);

OR2_X4 c3845(
.A1(net4083),
.A2(net11371),
.ZN(net4087)
);

OR2_X1 c3846(
.A1(net4081),
.A2(net3912),
.ZN(net4088)
);

INV_X32 c3847(
.A(net11107),
.ZN(net4089)
);

XNOR2_X2 c3848(
.A(net3093),
.B(net4085),
.ZN(net4090)
);

DFFR_X2 c3849(
.D(net4088),
.RN(net3165),
.CK(clk),
.Q(net4092),
.QN(net4091)
);

MUX2_X1 c3850(
.A(net3967),
.B(net3950),
.S(net3975),
.Z(net4093)
);

AND2_X4 c3851(
.A1(net4087),
.A2(net4075),
.ZN(net4094)
);

DFFRS_X1 c3852(
.D(net2077),
.RN(net3902),
.SN(net3084),
.CK(clk),
.Q(net4096),
.QN(net4095)
);

OAI21_X4 c3853(
.A(net4089),
.B1(net4093),
.B2(net4083),
.ZN(net4097)
);

INV_X4 c3854(
.A(net4060),
.ZN(net4098)
);

AND2_X1 c3855(
.A1(net4076),
.A2(net4079),
.ZN(net4099)
);

MUX2_X2 c3856(
.A(net4078),
.B(net4067),
.S(net3994),
.Z(net4100)
);

NAND2_X1 c3857(
.A1(net2122),
.A2(net4062),
.ZN(net4101)
);

NAND2_X2 c3858(
.A1(net4070),
.A2(net4095),
.ZN(net4102)
);

INV_X1 c3859(
.A(net4100),
.ZN(net4103)
);

NAND3_X4 c3860(
.A1(net4073),
.A2(net4080),
.A3(net4082),
.ZN(net4104)
);

OR3_X4 c3861(
.A1(net4074),
.A2(net4062),
.A3(net3989),
.ZN(net4105)
);

NAND2_X4 c3862(
.A1(net4022),
.A2(net4001),
.ZN(net4106)
);

INV_X2 c3863(
.A(net11106),
.ZN(net4107)
);

INV_X8 c3864(
.A(net4078),
.ZN(net4108)
);

INV_X16 c3865(
.A(net11084),
.ZN(net4109)
);

DFFS_X1 c3866(
.D(net4103),
.SN(net2987),
.CK(clk),
.Q(net4111),
.QN(net4110)
);

AND2_X2 c3867(
.A1(net4097),
.A2(net4073),
.ZN(net4112)
);

XOR2_X1 c3868(
.A(net4062),
.B(net4107),
.Z(net4113)
);

NOR2_X1 c3869(
.A1(net3989),
.A2(net11337),
.ZN(net4114)
);

INV_X32 c3870(
.A(net11130),
.ZN(net4115)
);

OR2_X2 c3871(
.A1(net4113),
.A2(net4089),
.ZN(net4116)
);

INV_X4 c3872(
.A(net11320),
.ZN(net4117)
);

INV_X1 c3873(
.A(net11338),
.ZN(net4118)
);

INV_X2 c3874(
.A(net11417),
.ZN(net4119)
);

AND3_X2 c3875(
.A1(net3950),
.A2(net4101),
.A3(net4119),
.ZN(net4120)
);

NOR2_X4 c3876(
.A1(net4106),
.A2(net3950),
.ZN(net4121)
);

NOR3_X1 c3877(
.A1(net4118),
.A2(net3120),
.A3(net4107),
.ZN(net4122)
);

NOR2_X2 c3878(
.A1(net4014),
.A2(net11176),
.ZN(net4123)
);

OR3_X2 c3879(
.A1(net2964),
.A2(net4024),
.A3(net4108),
.ZN(net4124)
);

AOI221_X1 c3880(
.A(net4057),
.B1(net4118),
.B2(net3977),
.C1(net4069),
.C2(net4084),
.ZN(net4125)
);

XOR2_X2 c3881(
.A(net4114),
.B(net3967),
.Z(net4126)
);

OAI21_X2 c3882(
.A(net4126),
.B1(net2144),
.B2(net3136),
.ZN(net4127)
);

OAI21_X1 c3883(
.A(net3122),
.B1(net4073),
.B2(net4108),
.ZN(net4128)
);

INV_X8 c3884(
.A(net10481),
.ZN(net4129)
);

XNOR2_X1 c3885(
.A(net4098),
.B(net4070),
.ZN(net4130)
);

AOI21_X2 c3886(
.A(net4129),
.B1(net4126),
.B2(net1193),
.ZN(net4131)
);

OR2_X4 c3887(
.A1(net4123),
.A2(net4095),
.ZN(net4132)
);

AOI21_X1 c3888(
.A(net4096),
.B1(net3063),
.B2(net4087),
.ZN(net4133)
);

AOI222_X2 c3889(
.A1(net4063),
.A2(net3108),
.B1(net4108),
.B2(net3156),
.C1(net3084),
.C2(net11422),
.ZN(net4134)
);

DFFRS_X2 c3890(
.D(net4036),
.RN(net3165),
.SN(net4109),
.CK(clk),
.Q(net4136),
.QN(net4135)
);

SDFF_X1 c3891(
.D(net4131),
.SE(net4074),
.SI(net4063),
.CK(clk),
.Q(net4138),
.QN(net4137)
);

INV_X16 c3892(
.A(net10387),
.ZN(net4139)
);

AOI21_X4 c3893(
.A(net4094),
.B1(net2964),
.B2(net4133),
.ZN(net4140)
);

OR2_X1 c3894(
.A1(net4139),
.A2(net11422),
.ZN(net4141)
);

OAI221_X1 c3895(
.A(net4109),
.B1(net4108),
.B2(net4088),
.C1(net4059),
.C2(net2153),
.ZN(net4142)
);

AND3_X1 c3896(
.A1(net3100),
.A2(net4141),
.A3(net11529),
.ZN(net4143)
);

OAI221_X4 c3897(
.A(net4093),
.B1(net4133),
.B2(net4141),
.C1(net4084),
.C2(net3981),
.ZN(net4144)
);

OAI22_X1 c3898(
.A1(net4104),
.A2(net4105),
.B1(net4015),
.B2(net11529),
.ZN(net4145)
);

XNOR2_X2 c3899(
.A(net4132),
.B(net11528),
.ZN(net4146)
);

NAND3_X1 c3900(
.A1(net4136),
.A2(net4146),
.A3(net10797),
.ZN(net4147)
);

AND2_X4 c3901(
.A1(net3154),
.A2(net4147),
.ZN(net4148)
);

AND2_X1 c3902(
.A1(net4121),
.A2(net4029),
.ZN(net4149)
);

INV_X32 c3903(
.A(net11093),
.ZN(net4150)
);

INV_X4 c3904(
.A(net10333),
.ZN(net4151)
);

NAND2_X1 c3905(
.A1(net2144),
.A2(net3258),
.ZN(net4152)
);

INV_X1 c3906(
.A(net4082),
.ZN(net4153)
);

NAND2_X2 c3907(
.A1(net86),
.A2(net2035),
.ZN(net4154)
);

NAND2_X4 c3908(
.A1(net1129),
.A2(net4110),
.ZN(net4155)
);

INV_X2 c3909(
.A(net11462),
.ZN(net4156)
);

AND2_X2 c3910(
.A1(net3163),
.A2(net3180),
.ZN(net4157)
);

XOR2_X1 c3911(
.A(net1951),
.B(net4030),
.Z(net4158)
);

NOR2_X1 c3912(
.A1(net2035),
.A2(net3243),
.ZN(net4159)
);

INV_X8 c3913(
.A(net4149),
.ZN(net4160)
);

INV_X16 c3914(
.A(net10443),
.ZN(net4161)
);

OR2_X2 c3915(
.A1(net3261),
.A2(net3149),
.ZN(net4162)
);

NOR2_X4 c3916(
.A1(net4066),
.A2(net3128),
.ZN(net4163)
);

INV_X32 c3917(
.A(net11276),
.ZN(net4164)
);

NOR2_X2 c3918(
.A1(net3191),
.A2(net3912),
.ZN(net4165)
);

XOR2_X2 c3919(
.A(net3084),
.B(net4079),
.Z(net4166)
);

XNOR2_X1 c3920(
.A(net2098),
.B(net4137),
.ZN(net4167)
);

NOR3_X4 c3921(
.A1(net3156),
.A2(net2098),
.A3(net3994),
.ZN(net4168)
);

NOR3_X2 c3922(
.A1(net4151),
.A2(net3915),
.A3(net2265),
.ZN(net4169)
);

OAI222_X1 c3923(
.A1(net3087),
.A2(net4159),
.B1(net1129),
.B2(net2098),
.C1(net4167),
.C2(net3235),
.ZN(net4170)
);

DFFS_X2 c3924(
.D(net3104),
.SN(net4160),
.CK(clk),
.Q(net4172),
.QN(net4171)
);

OR2_X4 c3925(
.A1(net4154),
.A2(net4164),
.ZN(net4173)
);

OR2_X1 c3926(
.A1(net3216),
.A2(net4167),
.ZN(net4174)
);

XNOR2_X2 c3927(
.A(net4059),
.B(net10686),
.ZN(net4175)
);

AND2_X4 c3928(
.A1(net4172),
.A2(net3915),
.ZN(net4176)
);

AND2_X1 c3929(
.A1(net4161),
.A2(net3993),
.ZN(net4177)
);

NAND2_X1 c3930(
.A1(net4177),
.A2(net11530),
.ZN(net4178)
);

AND3_X4 c3931(
.A1(net4172),
.A2(net3004),
.A3(net4167),
.ZN(net4179)
);

NAND2_X2 c3932(
.A1(net4162),
.A2(net4079),
.ZN(net4180)
);

NAND3_X2 c3933(
.A1(net4030),
.A2(net4178),
.A3(net11531),
.ZN(net4181)
);

OR3_X1 c3934(
.A1(net3167),
.A2(net2016),
.A3(net4181),
.ZN(net4182)
);

INV_X4 c3935(
.A(net11300),
.ZN(net4183)
);

INV_X1 c3936(
.A(net2231),
.ZN(net4184)
);

NAND2_X4 c3937(
.A1(net4148),
.A2(net3163),
.ZN(net4185)
);

AND2_X2 c3938(
.A1(net4176),
.A2(net4175),
.ZN(net4186)
);

XOR2_X1 c3939(
.A(net3054),
.B(net3063),
.Z(net4187)
);

MUX2_X1 c3940(
.A(net4102),
.B(net1220),
.S(net4107),
.Z(net4188)
);

INV_X2 c3941(
.A(net11472),
.ZN(net4189)
);

NOR2_X1 c3942(
.A1(net4184),
.A2(net1109),
.ZN(net4190)
);

OR2_X2 c3943(
.A1(net4165),
.A2(net11531),
.ZN(net4191)
);

INV_X8 c3944(
.A(net10445),
.ZN(net4192)
);

INV_X16 c3945(
.A(net11277),
.ZN(net4193)
);

NOR2_X4 c3946(
.A1(net4192),
.A2(net3207),
.ZN(net4194)
);

NOR2_X2 c3947(
.A1(net4193),
.A2(net4181),
.ZN(net4195)
);

XOR2_X2 c3948(
.A(net4164),
.B(net2198),
.Z(net4196)
);

XNOR2_X1 c3949(
.A(net4186),
.B(net4195),
.ZN(net4197)
);

OR2_X4 c3950(
.A1(net4195),
.A2(net4176),
.ZN(net4198)
);

INV_X32 c3951(
.A(net11182),
.ZN(net4199)
);

OR2_X1 c3952(
.A1(net3200),
.A2(net4183),
.ZN(net4200)
);

XNOR2_X2 c3953(
.A(net4115),
.B(net4052),
.ZN(net4201)
);

SDFF_X2 c3954(
.D(net4198),
.SE(net4167),
.SI(net3217),
.CK(clk),
.Q(net4203),
.QN(net4202)
);

AND2_X4 c3955(
.A1(net3180),
.A2(net4202),
.ZN(net4204)
);

AND2_X1 c3956(
.A1(net3253),
.A2(net11335),
.ZN(net4205)
);

NAND2_X1 c3957(
.A1(net4199),
.A2(net4082),
.ZN(net4206)
);

OAI21_X4 c3958(
.A(net4197),
.B1(net4196),
.B2(net4171),
.ZN(net4207)
);

INV_X4 c3959(
.A(net11056),
.ZN(net4208)
);

INV_X1 c3960(
.A(net11284),
.ZN(net4209)
);

NAND2_X2 c3961(
.A1(net4196),
.A2(net4079),
.ZN(net4210)
);

INV_X2 c3962(
.A(net11327),
.ZN(net4211)
);

NAND2_X4 c3963(
.A1(net4191),
.A2(net3969),
.ZN(net4212)
);

MUX2_X2 c3964(
.A(net4211),
.B(net4150),
.S(net2203),
.Z(net4213)
);

AND2_X2 c3965(
.A1(net3253),
.A2(net4193),
.ZN(net4214)
);

XOR2_X1 c3966(
.A(net3063),
.B(net4209),
.Z(net4215)
);

NAND3_X4 c3967(
.A1(net4204),
.A2(net4176),
.A3(net4214),
.ZN(net4216)
);

OR3_X4 c3968(
.A1(net4189),
.A2(net4198),
.A3(net4193),
.ZN(net4217)
);

NOR2_X1 c3969(
.A1(net4183),
.A2(net4206),
.ZN(net4218)
);

OR2_X2 c3970(
.A1(net4064),
.A2(net4197),
.ZN(net4219)
);

NOR2_X4 c3971(
.A1(net4085),
.A2(net10796),
.ZN(net4220)
);

INV_X8 c3972(
.A(net11301),
.ZN(net4221)
);

AND3_X2 c3973(
.A1(net4217),
.A2(net2153),
.A3(net4220),
.ZN(net4222)
);

NOR3_X1 c3974(
.A1(net4152),
.A2(net1269),
.A3(net4214),
.ZN(net4223)
);

OAI222_X4 c3975(
.A1(net4157),
.A2(net2261),
.B1(net4197),
.B2(net4159),
.C1(net4158),
.C2(net4167),
.ZN(net4224)
);

NOR2_X2 c3976(
.A1(net4185),
.A2(net4197),
.ZN(net4225)
);

OR3_X2 c3977(
.A1(net4222),
.A2(net4140),
.A3(net4210),
.ZN(net4226)
);

INV_X16 c3978(
.A(net11300),
.ZN(net4227)
);

OAI21_X2 c3979(
.A(net4184),
.B1(net4227),
.B2(net11191),
.ZN(net4228)
);

INV_X32 c3980(
.A(net10039),
.ZN(net4229)
);

OAI21_X1 c3981(
.A(net283),
.B1(net4217),
.B2(net4214),
.ZN(net4230)
);

INV_X4 c3982(
.A(net11462),
.ZN(net4231)
);

AOI21_X2 c3983(
.A(net4209),
.B1(net4221),
.B2(net10886),
.ZN(net4232)
);

XOR2_X2 c3984(
.A(net3207),
.B(net3994),
.Z(net4233)
);

INV_X1 c3985(
.A(net3349),
.ZN(net4234)
);

INV_X2 c3986(
.A(net11080),
.ZN(net4235)
);

OAI221_X2 c3987(
.A(net4203),
.B1(net4234),
.B2(net4110),
.C1(net4160),
.C2(net1217),
.ZN(net4236)
);

INV_X8 c3988(
.A(net10469),
.ZN(net4237)
);

XNOR2_X1 c3989(
.A(net2142),
.B(net4052),
.ZN(net4238)
);

AOI21_X1 c3990(
.A(net3330),
.B1(net3913),
.B2(net3328),
.ZN(net4239)
);

OR2_X4 c3991(
.A1(net4146),
.A2(net2277),
.ZN(net4240)
);

INV_X16 c3992(
.A(net10108),
.ZN(net4241)
);

OR2_X1 c3993(
.A1(net4218),
.A2(net3256),
.ZN(net4242)
);

INV_X32 c3994(
.A(net3333),
.ZN(net4243)
);

XNOR2_X2 c3995(
.A(net4138),
.B(net4235),
.ZN(net4244)
);

INV_X4 c3996(
.A(net4243),
.ZN(net4245)
);

AND2_X4 c3997(
.A1(net4233),
.A2(net4059),
.ZN(net4246)
);

AND2_X1 c3998(
.A1(net3291),
.A2(net1297),
.ZN(net4247)
);

AOI21_X4 c3999(
.A(net4238),
.B1(net3314),
.B2(net4233),
.ZN(net4248)
);

INV_X1 c4000(
.A(net3243),
.ZN(net4249)
);

INV_X2 c4001(
.A(net10694),
.ZN(net4250)
);

INV_X8 c4002(
.A(net11358),
.ZN(net4251)
);

INV_X16 c4003(
.A(net4175),
.ZN(net4252)
);

INV_X32 c4004(
.A(net2296),
.ZN(net4253)
);

NAND2_X1 c4005(
.A1(net1341),
.A2(net2317),
.ZN(net4254)
);

NAND2_X2 c4006(
.A1(net3994),
.A2(net4210),
.ZN(net4255)
);

INV_X4 c4007(
.A(net4080),
.ZN(net4256)
);

AND3_X1 c4008(
.A1(net4247),
.A2(net3349),
.A3(net10635),
.ZN(net4257)
);

NAND2_X4 c4009(
.A1(net3268),
.A2(net2153),
.ZN(net4258)
);

AND2_X2 c4010(
.A1(net4141),
.A2(net10952),
.ZN(net4259)
);

INV_X1 c4011(
.A(net3292),
.ZN(net4260)
);

INV_X2 c4012(
.A(net11358),
.ZN(net4261)
);

NAND3_X1 c4013(
.A1(net4052),
.A2(net3312),
.A3(net4254),
.ZN(net4262)
);

INV_X8 c4014(
.A(net10892),
.ZN(net4263)
);

XOR2_X1 c4015(
.A(net4260),
.B(net3330),
.Z(net4264)
);

NOR2_X1 c4016(
.A1(net4150),
.A2(net3326),
.ZN(net4265)
);

INV_X16 c4017(
.A(net11109),
.ZN(net4266)
);

NOR3_X4 c4018(
.A1(net4209),
.A2(net2277),
.A3(net11220),
.ZN(net4267)
);

INV_X32 c4019(
.A(net3312),
.ZN(net4268)
);

OR2_X2 c4020(
.A1(net4241),
.A2(net4254),
.ZN(net4269)
);

INV_X4 c4021(
.A(net4266),
.ZN(net4270)
);

NOR2_X4 c4022(
.A1(net3108),
.A2(net11191),
.ZN(net4271)
);

NOR3_X2 c4023(
.A1(net3328),
.A2(net4270),
.A3(net3264),
.ZN(net4272)
);

INV_X1 c4024(
.A(net10155),
.ZN(net4273)
);

NOR2_X2 c4025(
.A1(net4058),
.A2(net4260),
.ZN(net4274)
);

XOR2_X2 c4026(
.A(net4253),
.B(net4265),
.Z(net4275)
);

INV_X2 c4027(
.A(net4275),
.ZN(net4276)
);

INV_X8 c4028(
.A(net11338),
.ZN(net4277)
);

XNOR2_X1 c4029(
.A(net3309),
.B(net3305),
.ZN(net4278)
);

OR2_X4 c4030(
.A1(net4252),
.A2(net4235),
.ZN(net4279)
);

OR2_X1 c4031(
.A1(net4271),
.A2(net4274),
.ZN(net4280)
);

INV_X16 c4032(
.A(net10409),
.ZN(net4281)
);

XNOR2_X2 c4033(
.A(net4229),
.B(net4272),
.ZN(net4282)
);

AND2_X4 c4034(
.A1(net3912),
.A2(net4277),
.ZN(net4283)
);

DFFRS_X1 c4035(
.D(net4246),
.RN(net4158),
.SN(net4254),
.CK(clk),
.Q(net4285),
.QN(net4284)
);

AND2_X1 c4036(
.A1(net4231),
.A2(net4277),
.ZN(net4286)
);

AND3_X4 c4037(
.A1(net4141),
.A2(net4111),
.A3(net4253),
.ZN(net4287)
);

INV_X32 c4038(
.A(net10261),
.ZN(net4288)
);

NAND2_X1 c4039(
.A1(net4268),
.A2(net4156),
.ZN(net4289)
);

DFFRS_X2 c4040(
.D(net4284),
.RN(net4071),
.SN(net10687),
.CK(clk),
.Q(net4291),
.QN(net4290)
);

NAND3_X2 c4041(
.A1(net4247),
.A2(net2351),
.A3(net4284),
.ZN(net4292)
);

NAND2_X2 c4042(
.A1(net4278),
.A2(net4279),
.ZN(net4293)
);

NAND2_X4 c4043(
.A1(net4270),
.A2(net4282),
.ZN(net4294)
);

AND2_X2 c4044(
.A1(net4079),
.A2(net4272),
.ZN(net4295)
);

DFFR_X1 c4045(
.D(net4254),
.RN(net4295),
.CK(clk),
.Q(net4297),
.QN(net4296)
);

OR3_X1 c4046(
.A1(net4296),
.A2(net4260),
.A3(net11323),
.ZN(net4298)
);

INV_X4 c4047(
.A(net10107),
.ZN(net4299)
);

AND4_X2 c4048(
.A1(net4299),
.A2(net4293),
.A3(net4273),
.A4(net4277),
.ZN(net4300)
);

MUX2_X1 c4049(
.A(net4300),
.B(net4263),
.S(net4298),
.Z(net4301)
);

OAI21_X4 c4050(
.A(net4240),
.B1(net4296),
.B2(net11323),
.ZN(net4302)
);

XOR2_X1 c4051(
.A(net3243),
.B(net11220),
.Z(net4303)
);

NOR2_X1 c4052(
.A1(net3263),
.A2(net2296),
.ZN(net4304)
);

MUX2_X2 c4053(
.A(net4215),
.B(net4295),
.S(net4254),
.Z(net4305)
);

OR2_X2 c4054(
.A1(net3166),
.A2(net4263),
.ZN(net4306)
);

SDFF_X1 c4055(
.D(net4167),
.SE(net4306),
.SI(net4297),
.CK(clk),
.Q(net4308),
.QN(net4307)
);

NAND3_X4 c4056(
.A1(net3314),
.A2(net4298),
.A3(net4273),
.ZN(net4309)
);

OR3_X4 c4057(
.A1(net4294),
.A2(net4291),
.A3(net4273),
.ZN(net4310)
);

SDFFR_X1 c4058(
.D(net4297),
.RN(net4194),
.SE(net4168),
.SI(net10748),
.CK(clk),
.Q(net4312),
.QN(net4311)
);

AND3_X2 c4059(
.A1(net4310),
.A2(net4277),
.A3(net4303),
.ZN(net4313)
);

NOR3_X1 c4060(
.A1(net4288),
.A2(net3170),
.A3(net4311),
.ZN(net4314)
);

OR3_X2 c4061(
.A1(net4308),
.A2(net4313),
.A3(net4168),
.ZN(net4315)
);

OAI21_X2 c4062(
.A(net4289),
.B1(net4279),
.B2(net4313),
.ZN(net4316)
);

SDFF_X2 c4063(
.D(net4313),
.SE(net4309),
.SI(net4303),
.CK(clk),
.Q(net4318),
.QN(net4317)
);

OAI222_X2 c4064(
.A1(net4314),
.A2(net4168),
.B1(net4307),
.B2(net4306),
.C1(net4263),
.C2(net4245),
.ZN(net4319)
);

OAI21_X1 c4065(
.A(net4257),
.B1(net4290),
.B2(net10951),
.ZN(net4320)
);

DFFRS_X1 c4066(
.D(net4168),
.RN(net4270),
.SN(net11405),
.CK(clk),
.Q(net4322),
.QN(net4321)
);

AOI222_X1 c4067(
.A1(net4389),
.A2(net3356),
.B1(net3413),
.B2(net4407),
.C1(net3341),
.C2(net2280),
.ZN(net4323)
);

NOR2_X4 c4068(
.A1(net4387),
.A2(net4407),
.ZN(net4324)
);

NOR2_X2 c4069(
.A1(net4406),
.A2(net4405),
.ZN(net4325)
);

XOR2_X2 c4070(
.A(net4382),
.B(net4362),
.Z(net4326)
);

DFFRS_X2 c4071(
.D(net4377),
.RN(net3413),
.SN(net3408),
.CK(clk),
.Q(net4328),
.QN(net4327)
);

AND4_X1 c4072(
.A1(net2265),
.A2(net4405),
.A3(net4364),
.A4(net4158),
.ZN(net4329)
);

AOI21_X2 c4073(
.A(net4309),
.B1(net4326),
.B2(net4355),
.ZN(net4330)
);

XNOR2_X1 c4074(
.A(net4409),
.B(net4362),
.ZN(net4331)
);

OR2_X4 c4075(
.A1(net4402),
.A2(net4372),
.ZN(net4332)
);

OR2_X1 c4076(
.A1(net4326),
.A2(net3382),
.ZN(net4333)
);

AOI21_X1 c4077(
.A(net4411),
.B1(net4333),
.B2(net4332),
.ZN(net4334)
);

AOI21_X4 c4078(
.A(net4400),
.B1(net4286),
.B2(net11311),
.ZN(net4335)
);

XNOR2_X2 c4079(
.A(net4386),
.B(net4249),
.ZN(net4336)
);

AND2_X4 c4080(
.A1(net4359),
.A2(net4293),
.ZN(net4337)
);

AND2_X1 c4081(
.A1(net4329),
.A2(net4407),
.ZN(net4338)
);

NAND2_X1 c4082(
.A1(net4325),
.A2(net4402),
.ZN(net4339)
);

NAND2_X2 c4083(
.A1(net4372),
.A2(net4333),
.ZN(net4340)
);

INV_X1 c4084(
.A(net4356),
.ZN(net4341)
);

DFFR_X2 c4085(
.D(net4338),
.RN(net3397),
.CK(clk),
.Q(net4343),
.QN(net4342)
);

AND3_X1 c4086(
.A1(net3408),
.A2(net4329),
.A3(net4302),
.ZN(net4344)
);

NAND3_X1 c4087(
.A1(net4343),
.A2(net4356),
.A3(net4397),
.ZN(net4345)
);

NOR3_X4 c4088(
.A1(net4390),
.A2(net4379),
.A3(net4340),
.ZN(net4346)
);

INV_X2 c4089(
.A(net4370),
.ZN(net4347)
);

NAND2_X4 c4090(
.A1(net4335),
.A2(net3332),
.ZN(net4348)
);

AOI222_X4 c4091(
.A1(net4287),
.A2(net4327),
.B1(net3407),
.B2(net4298),
.C1(net4272),
.C2(net3425),
.ZN(net4349)
);

NOR3_X2 c4092(
.A1(net2383),
.A2(net4342),
.A3(net4348),
.ZN(net4350)
);

AND3_X4 c4093(
.A1(net4345),
.A2(net4371),
.A3(net11311),
.ZN(net4351)
);

NAND3_X2 c4094(
.A1(net4339),
.A2(net4345),
.A3(net4349),
.ZN(net4352)
);

OR3_X1 c4095(
.A1(net4339),
.A2(net4258),
.A3(net11290),
.ZN(net4353)
);

AND2_X2 c4096(
.A1(net4333),
.A2(net11290),
.ZN(net4354)
);

SDFF_X1 c4097(
.D(net4028),
.SE(net3424),
.SI(net10636),
.CK(clk),
.Q(net4356),
.QN(net4355)
);

XOR2_X1 c4098(
.A(net1922),
.B(net4298),
.Z(net4357)
);

NOR2_X1 c4099(
.A1(net4111),
.A2(net4272),
.ZN(net4358)
);

INV_X8 c4100(
.A(net4358),
.ZN(net4359)
);

INV_X16 c4101(
.A(net11016),
.ZN(net4360)
);

INV_X32 c4102(
.A(net2280),
.ZN(net4361)
);

INV_X4 c4103(
.A(net9722),
.ZN(net4362)
);

INV_X1 c4104(
.A(net9721),
.ZN(net4363)
);

INV_X2 c4105(
.A(net11410),
.ZN(net4364)
);

OR2_X2 c4106(
.A1(net3383),
.A2(net1254),
.ZN(net4365)
);

INV_X8 c4107(
.A(net3424),
.ZN(net4366)
);

INV_X16 c4108(
.A(net9842),
.ZN(net4367)
);

INV_X32 c4109(
.A(net11079),
.ZN(net4368)
);

NOR2_X4 c4110(
.A1(net4259),
.A2(net4272),
.ZN(net4369)
);

INV_X4 c4111(
.A(net4286),
.ZN(net4370)
);

NOR2_X2 c4112(
.A1(net3390),
.A2(net3406),
.ZN(net4371)
);

XOR2_X2 c4113(
.A(net4318),
.B(net1412),
.Z(net4372)
);

XNOR2_X1 c4114(
.A(net3433),
.B(net4360),
.ZN(net4373)
);

MUX2_X1 c4115(
.A(net3334),
.B(net4285),
.S(net3982),
.Z(net4374)
);

OR2_X4 c4116(
.A1(net4371),
.A2(net4317),
.ZN(net4375)
);

INV_X1 c4117(
.A(net3356),
.ZN(net4376)
);

OR2_X1 c4118(
.A1(net4281),
.A2(net4245),
.ZN(net4377)
);

INV_X2 c4119(
.A(net2382),
.ZN(net4378)
);

DFFS_X1 c4120(
.D(net4377),
.SN(net4301),
.CK(clk),
.Q(net4380),
.QN(net4379)
);

OAI21_X4 c4121(
.A(net369),
.B1(net4370),
.B2(net4085),
.ZN(net4381)
);

XNOR2_X2 c4122(
.A(net4380),
.B(net4158),
.ZN(net4382)
);

MUX2_X2 c4123(
.A(net4304),
.B(net4377),
.S(net3433),
.Z(net4383)
);

NAND3_X4 c4124(
.A1(net3332),
.A2(net4279),
.A3(net2382),
.ZN(net4384)
);

AND2_X4 c4125(
.A1(net4370),
.A2(net2382),
.ZN(net4385)
);

INV_X8 c4126(
.A(net10319),
.ZN(net4386)
);

AOI22_X4 c4127(
.A1(net4368),
.A2(net3433),
.B1(net4384),
.B2(net2328),
.ZN(net4387)
);

AND2_X1 c4128(
.A1(net4361),
.A2(net3334),
.ZN(net4388)
);

NAND2_X1 c4129(
.A1(net4387),
.A2(net2411),
.ZN(net4389)
);

NAND2_X2 c4130(
.A1(net4279),
.A2(net4318),
.ZN(net4390)
);

INV_X16 c4131(
.A(net4385),
.ZN(net4391)
);

INV_X32 c4132(
.A(net4362),
.ZN(net4392)
);

NAND2_X4 c4133(
.A1(net3982),
.A2(net3390),
.ZN(net4393)
);

AND2_X2 c4134(
.A1(net4285),
.A2(net4378),
.ZN(net4394)
);

XOR2_X1 c4135(
.A(net4385),
.B(net4376),
.Z(net4395)
);

INV_X4 c4136(
.A(net10440),
.ZN(net4396)
);

NOR2_X1 c4137(
.A1(net1466),
.A2(net4382),
.ZN(net4397)
);

INV_X1 c4138(
.A(net11285),
.ZN(net4398)
);

INV_X2 c4139(
.A(net11081),
.ZN(net4399)
);

SDFF_X2 c4140(
.D(net4357),
.SE(net3355),
.SI(net2328),
.CK(clk),
.Q(net4401),
.QN(net4400)
);

INV_X8 c4141(
.A(net3382),
.ZN(net4402)
);

INV_X16 c4142(
.A(net10028),
.ZN(net4403)
);

DFFRS_X1 c4143(
.D(net1434),
.RN(net4395),
.SN(net3371),
.CK(clk),
.Q(net4405),
.QN(net4404)
);

OR2_X2 c4144(
.A1(net4272),
.A2(net4369),
.ZN(net4406)
);

NOR2_X4 c4145(
.A1(net4395),
.A2(net10899),
.ZN(net4407)
);

NOR2_X2 c4146(
.A1(net3365),
.A2(net2328),
.ZN(net4408)
);

XOR2_X2 c4147(
.A(net4369),
.B(net3258),
.Z(net4409)
);

XNOR2_X1 c4148(
.A(net4398),
.B(net467),
.ZN(net4410)
);

INV_X32 c4149(
.A(net10358),
.ZN(net4411)
);

INV_X4 c4150(
.A(net10285),
.ZN(net4412)
);

OR3_X4 c4151(
.A1(net4092),
.A2(net3407),
.A3(net10806),
.ZN(net4413)
);

INV_X1 c4152(
.A(net11179),
.ZN(net4414)
);

OR2_X4 c4153(
.A1(net3511),
.A2(net3520),
.ZN(net4415)
);

OR2_X1 c4154(
.A1(net3455),
.A2(net4410),
.ZN(net4416)
);

INV_X2 c4155(
.A(net4303),
.ZN(net4417)
);

XNOR2_X2 c4156(
.A(net3499),
.B(net4395),
.ZN(net4418)
);

AND2_X4 c4157(
.A1(net4332),
.A2(net4316),
.ZN(net4419)
);

INV_X8 c4158(
.A(net4378),
.ZN(net4420)
);

AND2_X1 c4159(
.A1(net3414),
.A2(net4331),
.ZN(net4421)
);

INV_X16 c4160(
.A(net4298),
.ZN(net4422)
);

INV_X32 c4161(
.A(net4348),
.ZN(net4423)
);

AND3_X2 c4162(
.A1(net4414),
.A2(net3520),
.A3(net4392),
.ZN(net4424)
);

NAND2_X1 c4163(
.A1(net3521),
.A2(net3397),
.ZN(net4425)
);

INV_X4 c4164(
.A(net11221),
.ZN(net4426)
);

NOR3_X1 c4165(
.A1(net4425),
.A2(net4349),
.A3(net4303),
.ZN(net4427)
);

OR3_X2 c4166(
.A1(net3460),
.A2(net4391),
.A3(net1513),
.ZN(net4428)
);

NAND2_X2 c4167(
.A1(net3457),
.A2(net2526),
.ZN(net4429)
);

NAND2_X4 c4168(
.A1(net4424),
.A2(net4360),
.ZN(net4430)
);

AND2_X2 c4169(
.A1(net4419),
.A2(net2469),
.ZN(net4431)
);

XOR2_X1 c4170(
.A(net4391),
.B(net4425),
.Z(net4432)
);

INV_X1 c4171(
.A(net466),
.ZN(net4433)
);

INV_X2 c4172(
.A(net10341),
.ZN(net4434)
);

NOR2_X1 c4173(
.A1(net4331),
.A2(net4426),
.ZN(net4435)
);

OR2_X2 c4174(
.A1(net4395),
.A2(net4396),
.ZN(net4436)
);

INV_X8 c4175(
.A(net3454),
.ZN(net4437)
);

INV_X16 c4176(
.A(net4367),
.ZN(net4438)
);

INV_X32 c4177(
.A(net10334),
.ZN(net4439)
);

INV_X4 c4178(
.A(net4429),
.ZN(net4440)
);

INV_X1 c4179(
.A(net10017),
.ZN(net4441)
);

INV_X2 c4180(
.A(net4354),
.ZN(net4442)
);

NOR2_X4 c4181(
.A1(net4439),
.A2(net4245),
.ZN(net4443)
);

NOR2_X2 c4182(
.A1(net3407),
.A2(net4245),
.ZN(net4444)
);

XOR2_X2 c4183(
.A(net4436),
.B(net4442),
.Z(net4445)
);

INV_X8 c4184(
.A(net4433),
.ZN(net4446)
);

OAI21_X2 c4185(
.A(net2485),
.B1(net1530),
.B2(net4442),
.ZN(net4447)
);

XNOR2_X1 c4186(
.A(net4417),
.B(net4423),
.ZN(net4448)
);

DFFRS_X2 c4187(
.D(net3476),
.RN(net4425),
.SN(net372),
.CK(clk),
.Q(net4450),
.QN(net4449)
);

INV_X16 c4188(
.A(net4418),
.ZN(net4451)
);

OR2_X4 c4189(
.A1(net2542),
.A2(net3520),
.ZN(net4452)
);

OAI21_X1 c4190(
.A(net3410),
.B1(net4378),
.B2(net3448),
.ZN(net4453)
);

AOI21_X2 c4191(
.A(net4448),
.B1(net3477),
.B2(net3460),
.ZN(net4454)
);

SDFF_X1 c4192(
.D(net2371),
.SE(net4431),
.SI(net4416),
.CK(clk),
.Q(net4456),
.QN(net4455)
);

OR2_X1 c4193(
.A1(net4450),
.A2(net4332),
.ZN(net4457)
);

XNOR2_X2 c4194(
.A(net4453),
.B(net4451),
.ZN(net4458)
);

AND2_X4 c4195(
.A1(net4454),
.A2(net11457),
.ZN(net4459)
);

AOI21_X1 c4196(
.A(net4433),
.B1(net4454),
.B2(net10949),
.ZN(net4460)
);

INV_X32 c4197(
.A(net10433),
.ZN(net4461)
);

INV_X4 c4198(
.A(net9905),
.ZN(net4462)
);

INV_X1 c4199(
.A(net4454),
.ZN(net4463)
);

AOI21_X4 c4200(
.A(net4444),
.B1(net4434),
.B2(net4303),
.ZN(net4464)
);

AND2_X1 c4201(
.A1(net4456),
.A2(net4441),
.ZN(net4465)
);

NAND2_X1 c4202(
.A1(net3509),
.A2(net11467),
.ZN(net4466)
);

INV_X2 c4203(
.A(net10156),
.ZN(net4467)
);

AND3_X1 c4204(
.A1(net4440),
.A2(net4220),
.A3(net4302),
.ZN(net4468)
);

NAND3_X1 c4205(
.A1(net4466),
.A2(net4454),
.A3(net4449),
.ZN(net4469)
);

NAND2_X2 c4206(
.A1(net4467),
.A2(net4448),
.ZN(net4470)
);

NOR3_X4 c4207(
.A1(net4344),
.A2(net4412),
.A3(net3414),
.ZN(net4471)
);

NAND2_X4 c4208(
.A1(net4468),
.A2(net4426),
.ZN(net4472)
);

AND2_X2 c4209(
.A1(net4420),
.A2(net4454),
.ZN(net4473)
);

SDFF_X2 c4210(
.D(net3264),
.SE(net4467),
.SI(net2520),
.CK(clk),
.Q(net4475),
.QN(net4474)
);

XOR2_X1 c4211(
.A(net4443),
.B(net4455),
.Z(net4476)
);

NOR2_X1 c4212(
.A1(net4451),
.A2(net11278),
.ZN(net4477)
);

INV_X8 c4213(
.A(net11459),
.ZN(net4478)
);

INV_X16 c4214(
.A(net11179),
.ZN(net4479)
);

AOI221_X4 c4215(
.A(net1418),
.B1(net4456),
.B2(net4476),
.C1(net3264),
.C2(net2461),
.ZN(net4480)
);

DFFRS_X1 c4216(
.D(net4412),
.RN(net3341),
.SN(net2351),
.CK(clk),
.Q(net4482),
.QN(net4481)
);

OR2_X2 c4217(
.A1(net4461),
.A2(net4462),
.ZN(net4483)
);

NOR3_X2 c4218(
.A1(net4462),
.A2(net4448),
.A3(net4483),
.ZN(net4484)
);

AND3_X4 c4219(
.A1(net4422),
.A2(net4472),
.A3(net4470),
.ZN(net4485)
);

NOR2_X4 c4220(
.A1(net4421),
.A2(net4472),
.ZN(net4486)
);

NOR2_X2 c4221(
.A1(net4469),
.A2(net4486),
.ZN(net4487)
);

NAND3_X2 c4222(
.A1(net4478),
.A2(net4450),
.A3(net4452),
.ZN(net4488)
);

OR3_X1 c4223(
.A1(net3477),
.A2(net4467),
.A3(net4474),
.ZN(net4489)
);

XOR2_X2 c4224(
.A(net4484),
.B(net4489),
.Z(net4490)
);

MUX2_X1 c4225(
.A(net4441),
.B(net4490),
.S(net3264),
.Z(net4491)
);

OAI21_X4 c4226(
.A(net4473),
.B1(net4486),
.B2(net11352),
.ZN(net4492)
);

XNOR2_X1 c4227(
.A(net4490),
.B(net4473),
.ZN(net4493)
);

MUX2_X2 c4228(
.A(net4475),
.B(net4493),
.S(net4488),
.Z(net4494)
);

OR2_X4 c4229(
.A1(net4433),
.A2(net11476),
.ZN(net4495)
);

NAND3_X4 c4230(
.A1(net4494),
.A2(net4490),
.A3(net4483),
.ZN(net4496)
);

DFFRS_X2 c4231(
.D(net4306),
.RN(net4489),
.SN(net4491),
.CK(clk),
.Q(net4498),
.QN(net4497)
);

OR3_X4 c4232(
.A1(net4492),
.A2(net4498),
.A3(net4495),
.ZN(net4499)
);

AND3_X2 c4233(
.A1(net4491),
.A2(net4316),
.A3(net1513),
.ZN(net4500)
);

INV_X32 c4234(
.A(net4470),
.ZN(net4501)
);

NOR3_X1 c4235(
.A1(net4293),
.A2(net3548),
.A3(net3604),
.ZN(net4502)
);

INV_X4 c4236(
.A(net3591),
.ZN(net4503)
);

INV_X1 c4237(
.A(net3509),
.ZN(net4504)
);

OR2_X1 c4238(
.A1(net4457),
.A2(net11532),
.ZN(net4505)
);

XNOR2_X2 c4239(
.A(net4489),
.B(net4487),
.ZN(net4506)
);

AND2_X4 c4240(
.A1(net3547),
.A2(net11523),
.ZN(net4507)
);

OR3_X2 c4241(
.A1(net2551),
.A2(net4458),
.A3(net654),
.ZN(net4508)
);

AND2_X1 c4242(
.A1(net3601),
.A2(net4470),
.ZN(net4509)
);

INV_X2 c4243(
.A(net4509),
.ZN(net4510)
);

OAI21_X2 c4244(
.A(net654),
.B1(net3600),
.B2(net2630),
.ZN(net4511)
);

NAND2_X1 c4245(
.A1(net3458),
.A2(net3547),
.ZN(net4512)
);

INV_X8 c4246(
.A(net11446),
.ZN(net4513)
);

NAND2_X2 c4247(
.A1(net2377),
.A2(net4428),
.ZN(net4514)
);

AOI221_X2 c4248(
.A(net4459),
.B1(net3543),
.B2(net2629),
.C1(net3594),
.C2(net11533),
.ZN(net4515)
);

NAND2_X4 c4249(
.A1(net589),
.A2(net4384),
.ZN(net4516)
);

AND2_X2 c4250(
.A1(net2532),
.A2(net4491),
.ZN(net4517)
);

XOR2_X1 c4251(
.A(net4428),
.B(net3555),
.Z(net4518)
);

INV_X16 c4252(
.A(net3471),
.ZN(net4519)
);

NOR2_X1 c4253(
.A1(net3341),
.A2(net4428),
.ZN(net4520)
);

INV_X32 c4254(
.A(net3567),
.ZN(net4521)
);

OR2_X2 c4255(
.A1(net1513),
.A2(net11532),
.ZN(net4522)
);

SDFFRS_X2 c4256(
.D(net4503),
.RN(net4500),
.SE(net3509),
.SI(net3341),
.SN(net3594),
.CK(clk),
.Q(net4524),
.QN(net4523)
);

NOR2_X4 c4257(
.A1(net4513),
.A2(net3598),
.ZN(net4525)
);

NOR2_X2 c4258(
.A1(net2567),
.A2(net3594),
.ZN(net4526)
);

OAI22_X4 c4259(
.A1(net1646),
.A2(net3585),
.B1(net3393),
.B2(net2593),
.ZN(net4527)
);

INV_X4 c4260(
.A(net4507),
.ZN(net4528)
);

XOR2_X2 c4261(
.A(net4510),
.B(net4501),
.Z(net4529)
);

INV_X1 c4262(
.A(net10254),
.ZN(net4530)
);

INV_X2 c4263(
.A(net4486),
.ZN(net4531)
);

INV_X8 c4264(
.A(net4376),
.ZN(net4532)
);

XNOR2_X1 c4265(
.A(net4464),
.B(net4505),
.ZN(net4533)
);

OR2_X4 c4266(
.A1(net4516),
.A2(net4302),
.ZN(net4534)
);

INV_X16 c4267(
.A(net2535),
.ZN(net4535)
);

INV_X32 c4268(
.A(net10227),
.ZN(net4536)
);

OR2_X1 c4269(
.A1(net4536),
.A2(net11372),
.ZN(net4537)
);

XNOR2_X2 c4270(
.A(net4529),
.B(net3567),
.ZN(net4538)
);

INV_X4 c4271(
.A(net10361),
.ZN(net4539)
);

AND2_X4 c4272(
.A1(net4452),
.A2(net4483),
.ZN(net4540)
);

AND2_X1 c4273(
.A1(net4522),
.A2(net4540),
.ZN(net4541)
);

NAND2_X1 c4274(
.A1(net3543),
.A2(net4540),
.ZN(net4542)
);

NAND2_X2 c4275(
.A1(net3526),
.A2(net4529),
.ZN(net4543)
);

NAND2_X4 c4276(
.A1(net4535),
.A2(net4526),
.ZN(net4544)
);

AND2_X2 c4277(
.A1(net4501),
.A2(net344),
.ZN(net4545)
);

INV_X1 c4278(
.A(net4511),
.ZN(net4546)
);

INV_X2 c4279(
.A(net4536),
.ZN(net4547)
);

SDFFR_X2 c4280(
.D(net4538),
.RN(net285),
.SE(net4501),
.SI(net3594),
.CK(clk),
.Q(net4549),
.QN(net4548)
);

INV_X8 c4281(
.A(net4528),
.ZN(net4550)
);

INV_X16 c4282(
.A(net11419),
.ZN(net4551)
);

XOR2_X1 c4283(
.A(net4521),
.B(net11372),
.Z(net4552)
);

NOR2_X1 c4284(
.A1(net4552),
.A2(net2380),
.ZN(net4553)
);

INV_X32 c4285(
.A(net11115),
.ZN(net4554)
);

OAI21_X1 c4286(
.A(net4505),
.B1(net4465),
.B2(net4452),
.ZN(net4555)
);

INV_X4 c4287(
.A(net4532),
.ZN(net4556)
);

OR2_X2 c4288(
.A1(net1530),
.A2(net4529),
.ZN(net4557)
);

INV_X1 c4289(
.A(net4531),
.ZN(net4558)
);

INV_X2 c4290(
.A(net11296),
.ZN(net4559)
);

AOI22_X2 c4291(
.A1(net4497),
.A2(net4541),
.B1(net4557),
.B2(net11457),
.ZN(net4560)
);

INV_X8 c4292(
.A(net11233),
.ZN(net4561)
);

NOR2_X4 c4293(
.A1(net4559),
.A2(net4442),
.ZN(net4562)
);

NOR2_X2 c4294(
.A1(net4546),
.A2(net4158),
.ZN(net4563)
);

AOI221_X1 c4295(
.A(net4553),
.B1(net3341),
.B2(net4561),
.C1(net3586),
.C2(net3594),
.ZN(net4564)
);

XOR2_X2 c4296(
.A(net4505),
.B(net10676),
.Z(net4565)
);

NAND4_X4 c4297(
.A1(net4551),
.A2(net3591),
.A3(net4487),
.A4(net3451),
.ZN(net4566)
);

AOI21_X2 c4298(
.A(net4556),
.B1(net3602),
.B2(net3418),
.ZN(net4567)
);

INV_X16 c4299(
.A(net10253),
.ZN(net4568)
);

INV_X32 c4300(
.A(net10398),
.ZN(net4569)
);

INV_X4 c4301(
.A(net11446),
.ZN(net4570)
);

SDFFS_X1 c4302(
.D(net4508),
.SE(net4558),
.SI(net4561),
.SN(net4539),
.CK(clk),
.Q(net4572),
.QN(net4571)
);

XNOR2_X1 c4303(
.A(net4549),
.B(net10876),
.ZN(net4573)
);

INV_X1 c4304(
.A(net11420),
.ZN(net4574)
);

AOI21_X1 c4305(
.A(net4515),
.B1(net4574),
.B2(net3341),
.ZN(net4575)
);

OAI211_X2 c4306(
.A(net4575),
.B(net4524),
.C1(net4539),
.C2(net4526),
.ZN(net4576)
);

INV_X2 c4307(
.A(net10384),
.ZN(net4577)
);

AOI21_X4 c4308(
.A(net4577),
.B1(net4574),
.B2(net4549),
.ZN(net4578)
);

OR2_X4 c4309(
.A1(net4545),
.A2(net11345),
.ZN(net4579)
);

OAI221_X1 c4310(
.A(net4561),
.B1(net4565),
.B2(net4536),
.C1(net4265),
.C2(net4542),
.ZN(net4580)
);

OR2_X1 c4311(
.A1(net4574),
.A2(net11038),
.ZN(net4581)
);

INV_X8 c4312(
.A(net10195),
.ZN(net4582)
);

XNOR2_X2 c4313(
.A(net4579),
.B(net4581),
.ZN(net4583)
);

OR4_X2 c4314(
.A1(net4582),
.A2(net4581),
.A3(net4565),
.A4(net4541),
.ZN(net4584)
);

AND2_X4 c4315(
.A1(net4561),
.A2(net11394),
.ZN(net4585)
);

DFFS_X2 c4316(
.D(net1728),
.SN(net3691),
.CK(clk),
.Q(net4587),
.QN(net4586)
);

AND2_X1 c4317(
.A1(net4463),
.A2(net4526),
.ZN(net4588)
);

AND3_X1 c4318(
.A1(net3660),
.A2(net654),
.A3(net4526),
.ZN(net4589)
);

INV_X16 c4319(
.A(net3129),
.ZN(net4590)
);

INV_X32 c4320(
.A(net9723),
.ZN(net4591)
);

INV_X4 c4321(
.A(net11490),
.ZN(net4592)
);

INV_X1 c4322(
.A(net4568),
.ZN(net4593)
);

NAND3_X1 c4323(
.A1(net3681),
.A2(net4590),
.A3(net4520),
.ZN(net4594)
);

INV_X2 c4324(
.A(net4580),
.ZN(net4595)
);

INV_X8 c4325(
.A(net2681),
.ZN(net4596)
);

INV_X16 c4326(
.A(net11471),
.ZN(net4597)
);

INV_X32 c4327(
.A(net9859),
.ZN(net4598)
);

INV_X4 c4328(
.A(net3652),
.ZN(net4599)
);

NAND2_X1 c4329(
.A1(net4598),
.A2(net10614),
.ZN(net4600)
);

NAND2_X2 c4330(
.A1(net4587),
.A2(net4588),
.ZN(net4601)
);

INV_X1 c4331(
.A(net9859),
.ZN(net4602)
);

INV_X2 c4332(
.A(net11533),
.ZN(net4603)
);

INV_X8 c4333(
.A(net9857),
.ZN(net4604)
);

INV_X16 c4334(
.A(net4599),
.ZN(net4605)
);

INV_X32 c4335(
.A(net9858),
.ZN(net4606)
);

INV_X4 c4336(
.A(net3585),
.ZN(net4607)
);

INV_X1 c4337(
.A(net9848),
.ZN(net4608)
);

INV_X2 c4338(
.A(net11449),
.ZN(net4609)
);

INV_X8 c4339(
.A(net4596),
.ZN(net4610)
);

AOI211_X1 c4340(
.A(net3637),
.B(net4465),
.C1(net4522),
.C2(net4598),
.ZN(net4611)
);

NAND2_X4 c4341(
.A1(net1729),
.A2(net4568),
.ZN(net4612)
);

INV_X16 c4342(
.A(net4487),
.ZN(net4613)
);

INV_X32 c4343(
.A(net2661),
.ZN(net4614)
);

INV_X4 c4344(
.A(net4498),
.ZN(net4615)
);

AND2_X2 c4345(
.A1(net3662),
.A2(net3635),
.ZN(net4616)
);

INV_X1 c4346(
.A(net9806),
.ZN(net4617)
);

XOR2_X1 c4347(
.A(net4598),
.B(net10779),
.Z(net4618)
);

INV_X2 c4348(
.A(net4316),
.ZN(net4619)
);

NOR3_X4 c4349(
.A1(net4600),
.A2(net4539),
.A3(net4522),
.ZN(net4620)
);

NOR3_X2 c4350(
.A1(net696),
.A2(net4608),
.A3(net4500),
.ZN(net4621)
);

AND3_X4 c4351(
.A1(net4609),
.A2(net3635),
.A3(net4619),
.ZN(net4622)
);

INV_X8 c4352(
.A(net9806),
.ZN(net4623)
);

NOR2_X1 c4353(
.A1(net4526),
.A2(net4590),
.ZN(net4624)
);

INV_X16 c4354(
.A(net3640),
.ZN(net4625)
);

INV_X32 c4355(
.A(net10446),
.ZN(net4626)
);

INV_X4 c4356(
.A(net9976),
.ZN(net4627)
);

INV_X1 c4357(
.A(net11360),
.ZN(net4628)
);

OR2_X2 c4358(
.A1(net2700),
.A2(net4620),
.ZN(net4629)
);

NOR2_X4 c4359(
.A1(net4522),
.A2(net4438),
.ZN(net4630)
);

INV_X2 c4360(
.A(net4570),
.ZN(net4631)
);

NOR2_X2 c4361(
.A1(net2380),
.A2(net10971),
.ZN(net4632)
);

XOR2_X2 c4362(
.A(net727),
.B(net2669),
.Z(net4633)
);

XNOR2_X1 c4363(
.A(net4324),
.B(net4633),
.ZN(net4634)
);

INV_X8 c4364(
.A(net4632),
.ZN(net4635)
);

OR2_X4 c4365(
.A1(net4593),
.A2(net4602),
.ZN(net4636)
);

INV_X16 c4366(
.A(net11031),
.ZN(net4637)
);

INV_X32 c4367(
.A(net10009),
.ZN(net4638)
);

INV_X4 c4368(
.A(net10948),
.ZN(net4639)
);

INV_X1 c4369(
.A(net10900),
.ZN(net4640)
);

INV_X2 c4370(
.A(net4634),
.ZN(net4641)
);

INV_X8 c4371(
.A(net4619),
.ZN(net4642)
);

INV_X16 c4372(
.A(net4302),
.ZN(net4643)
);

OR2_X1 c4373(
.A1(net4625),
.A2(net4599),
.ZN(net4644)
);

XNOR2_X2 c4374(
.A(net3555),
.B(net3662),
.ZN(net4645)
);

INV_X32 c4375(
.A(net9723),
.ZN(net4646)
);

INV_X4 c4376(
.A(net4631),
.ZN(net4647)
);

OAI221_X4 c4377(
.A(net4639),
.B1(net2719),
.B2(net4637),
.C1(net4588),
.C2(net4495),
.ZN(net4648)
);

AND2_X4 c4378(
.A1(net4606),
.A2(net3692),
.ZN(net4649)
);

NAND3_X2 c4379(
.A1(net4607),
.A2(net4638),
.A3(net2594),
.ZN(net4650)
);

AND2_X1 c4380(
.A1(net4618),
.A2(net4488),
.ZN(net4651)
);

INV_X1 c4381(
.A(net4645),
.ZN(net4652)
);

OAI33_X1 c4382(
.A1(net4651),
.A2(net4334),
.A3(net4620),
.B1(net4526),
.B2(net3691),
.B3(net4592),
.ZN(net4653)
);

OR3_X1 c4383(
.A1(net4624),
.A2(net4649),
.A3(net4640),
.ZN(net4654)
);

MUX2_X1 c4384(
.A(net4617),
.B(net4639),
.S(net10793),
.Z(net4655)
);

INV_X2 c4385(
.A(net11189),
.ZN(net4656)
);

INV_X8 c4386(
.A(net11411),
.ZN(net4657)
);

NAND2_X1 c4387(
.A1(net4617),
.A2(net4643),
.ZN(net4658)
);

INV_X16 c4388(
.A(net11490),
.ZN(net4659)
);

NAND2_X2 c4389(
.A1(net4647),
.A2(net4658),
.ZN(net4660)
);

NAND2_X4 c4390(
.A1(net4602),
.A2(net4643),
.ZN(net4661)
);

OAI21_X4 c4391(
.A(net4644),
.B1(net4586),
.B2(net11452),
.ZN(net4662)
);

AND2_X2 c4392(
.A1(net4630),
.A2(net11232),
.ZN(net4663)
);

MUX2_X2 c4393(
.A(net1309),
.B(net4625),
.S(net11232),
.Z(net4664)
);

OAI221_X2 c4394(
.A(net4605),
.B1(net4316),
.B2(net4568),
.C1(net4608),
.C2(net3615),
.ZN(net4665)
);

AOI221_X4 c4395(
.A(net2669),
.B1(net4641),
.B2(net4664),
.C1(net4526),
.C2(net11485),
.ZN(net4666)
);

NAND4_X2 c4396(
.A1(net4656),
.A2(net4660),
.A3(net4598),
.A4(net4664),
.ZN(net4667)
);

NAND3_X4 c4397(
.A1(net4640),
.A2(net4651),
.A3(net4664),
.ZN(net4668)
);

AOI222_X2 c4398(
.A1(net4657),
.A2(net4656),
.B1(net4665),
.B2(net4614),
.C1(net4620),
.C2(net4664),
.ZN(net4669)
);

OR3_X4 c4399(
.A1(net3746),
.A2(net4542),
.A3(net3767),
.ZN(net4670)
);

XOR2_X1 c4400(
.A(net4572),
.B(net4334),
.Z(net4671)
);

SDFF_X1 c4401(
.D(net2606),
.SE(net2806),
.SI(net11030),
.CK(clk),
.Q(net4673),
.QN(net4672)
);

INV_X32 c4402(
.A(net4430),
.ZN(net4674)
);

NOR2_X1 c4403(
.A1(net2763),
.A2(net2670),
.ZN(out1)
);

OR2_X2 c4404(
.A1(net2670),
.A2(net1636),
.ZN(net4675)
);

INV_X4 c4405(
.A(net11456),
.ZN(net4676)
);

NOR2_X4 c4406(
.A1(net4675),
.A2(net10592),
.ZN(net4677)
);

NOR2_X2 c4407(
.A1(net4590),
.A2(net4643),
.ZN(net4678)
);

XOR2_X2 c4408(
.A(net4671),
.B(net3626),
.Z(net4679)
);

INV_X1 c4409(
.A(net10118),
.ZN(net4680)
);

INV_X2 c4410(
.A(net1816),
.ZN(net4681)
);

DFFR_X1 c4411(
.D(net3635),
.RN(net3767),
.CK(clk),
.Q(net4683),
.QN(net4682)
);

XNOR2_X1 c4412(
.A(net4635),
.B(net1743),
.ZN(net4684)
);

INV_X8 c4413(
.A(net11379),
.ZN(net4685)
);

OR2_X4 c4414(
.A1(net4650),
.A2(net4542),
.ZN(net4686)
);

OR2_X1 c4415(
.A1(net4685),
.A2(net4680),
.ZN(net4687)
);

XNOR2_X2 c4416(
.A(net3619),
.B(net4665),
.ZN(net4688)
);

AND2_X4 c4417(
.A1(net2806),
.A2(net3541),
.ZN(net4689)
);

AND2_X1 c4418(
.A1(net701),
.A2(net1743),
.ZN(net4690)
);

AND3_X2 c4419(
.A1(net3728),
.A2(net4668),
.A3(net701),
.ZN(net4691)
);

INV_X16 c4420(
.A(net11364),
.ZN(net4692)
);

NAND2_X1 c4421(
.A1(net4585),
.A2(net701),
.ZN(net4693)
);

NOR3_X1 c4422(
.A1(net4686),
.A2(net1636),
.A3(net4321),
.ZN(net4694)
);

NAND2_X2 c4423(
.A1(net3752),
.A2(net826),
.ZN(net4695)
);

NAND2_X4 c4424(
.A1(net4643),
.A2(net4689),
.ZN(net4696)
);

OR3_X2 c4425(
.A1(net694),
.A2(net4675),
.A3(net4681),
.ZN(net4697)
);

INV_X32 c4426(
.A(net9880),
.ZN(net4698)
);

OAI21_X2 c4427(
.A(net4384),
.B1(net1816),
.B2(net4614),
.ZN(net4699)
);

INV_X4 c4428(
.A(net1687),
.ZN(net4700)
);

AND2_X2 c4429(
.A1(net2557),
.A2(net4590),
.ZN(net4701)
);

SDFF_X2 c4430(
.D(net3780),
.SE(net785),
.SI(net1562),
.CK(clk),
.Q(net4703),
.QN(net4702)
);

XOR2_X1 c4431(
.A(net826),
.B(net4693),
.Z(net4704)
);

NOR2_X1 c4432(
.A1(net3544),
.A2(net4700),
.ZN(net4705)
);

OR4_X4 c4433(
.A1(net3737),
.A2(net2719),
.A3(net4672),
.A4(net4571),
.ZN(net4706)
);

OR2_X2 c4434(
.A1(net4689),
.A2(net4697),
.ZN(net4707)
);

NOR2_X4 c4435(
.A1(net810),
.A2(net2799),
.ZN(net4708)
);

NOR2_X2 c4436(
.A1(net2461),
.A2(net4680),
.ZN(net4709)
);

INV_X1 c4437(
.A(net10114),
.ZN(net4710)
);

XOR2_X2 c4438(
.A(net4690),
.B(net3765),
.Z(net4711)
);

INV_X2 c4439(
.A(net11317),
.ZN(net4712)
);

XNOR2_X1 c4440(
.A(net4681),
.B(net3723),
.ZN(net4713)
);

DFFRS_X1 c4441(
.D(net3773),
.RN(net4674),
.SN(net3742),
.CK(clk),
.Q(net4715),
.QN(net4714)
);

OAI22_X2 c4442(
.A1(net4692),
.A2(net2771),
.B1(net4674),
.B2(net4704),
.ZN(net4716)
);

OR2_X4 c4443(
.A1(net1791),
.A2(net4438),
.ZN(net4717)
);

OR2_X1 c4444(
.A1(net4670),
.A2(net4673),
.ZN(net4718)
);

XNOR2_X2 c4445(
.A(net3541),
.B(net4713),
.ZN(net4719)
);

AND2_X4 c4446(
.A1(net4684),
.A2(net10528),
.ZN(net4720)
);

OAI21_X1 c4447(
.A(net2508),
.B1(net2670),
.B2(net4715),
.ZN(net4721)
);

AND2_X1 c4448(
.A1(net4698),
.A2(net4719),
.ZN(net4722)
);

NAND2_X1 c4449(
.A1(net4698),
.A2(net11485),
.ZN(net4723)
);

AOI21_X2 c4450(
.A(net4718),
.B1(net4711),
.B2(net4658),
.ZN(net4724)
);

NAND2_X2 c4451(
.A1(net4694),
.A2(net4717),
.ZN(net4725)
);

AOI21_X1 c4452(
.A(net4722),
.B1(net4723),
.B2(net4680),
.ZN(net4726)
);

INV_X8 c4453(
.A(net9920),
.ZN(net4727)
);

DFFRS_X2 c4454(
.D(net4550),
.RN(net4726),
.SN(net3775),
.CK(clk),
.Q(net4729),
.QN(net4728)
);

AOI21_X4 c4455(
.A(net4677),
.B1(net4728),
.B2(net4681),
.ZN(net4730)
);

NAND2_X4 c4456(
.A1(net2739),
.A2(net4728),
.ZN(net4731)
);

AND3_X1 c4457(
.A1(net4706),
.A2(net4650),
.A3(net4715),
.ZN(net4732)
);

SDFF_X1 c4458(
.D(net4588),
.SE(net4723),
.SI(net4683),
.CK(clk),
.Q(net4734),
.QN(net4733)
);

NAND3_X1 c4459(
.A1(net4701),
.A2(net4680),
.A3(net4717),
.ZN(net4735)
);

AND2_X2 c4460(
.A1(net4705),
.A2(net4735),
.ZN(net4736)
);

NOR3_X4 c4461(
.A1(net2704),
.A2(net4731),
.A3(net4670),
.ZN(net4737)
);

SDFF_X2 c4462(
.D(net4726),
.SE(net1802),
.SI(net4734),
.CK(clk),
.Q(net4739),
.QN(net4738)
);

XOR2_X1 c4463(
.A(net4696),
.B(net4733),
.Z(net4740)
);

DFFRS_X1 c4464(
.D(net4711),
.RN(net4737),
.SN(net4740),
.CK(clk),
.Q(net4742),
.QN(net4741)
);

AOI221_X2 c4465(
.A(net4695),
.B1(net4673),
.B2(net4741),
.C1(net3615),
.C2(net4684),
.ZN(net4743)
);

NOR3_X2 c4466(
.A1(net4709),
.A2(net4737),
.A3(net4741),
.ZN(net4744)
);

AND3_X4 c4467(
.A1(net4721),
.A2(net2735),
.A3(net1743),
.ZN(net4745)
);

NAND3_X2 c4468(
.A1(net4708),
.A2(net4738),
.A3(net4732),
.ZN(net4746)
);

OR3_X1 c4469(
.A1(net4734),
.A2(net4739),
.A3(net4743),
.ZN(net4747)
);

NOR2_X1 c4470(
.A1(net4743),
.A2(net4710),
.ZN(net4748)
);

MUX2_X1 c4471(
.A(net4748),
.B(net4747),
.S(net3728),
.Z(net4749)
);

INV_X16 c4472(
.A(net11456),
.ZN(net4750)
);

OAI21_X4 c4473(
.A(net2771),
.B1(net4678),
.B2(net4723),
.ZN(net4751)
);

MUX2_X2 c4474(
.A(net4746),
.B(net4684),
.S(net4698),
.Z(net4752)
);

OR2_X2 c4475(
.A1(net4750),
.A2(net4703),
.ZN(net4753)
);

NOR2_X4 c4476(
.A1(net4438),
.A2(net4727),
.ZN(net4754)
);

NAND3_X4 c4477(
.A1(net3745),
.A2(net4740),
.A3(net4719),
.ZN(net4755)
);

SDFFS_X2 c4478(
.D(net4649),
.SE(net4738),
.SI(net4755),
.SN(net10983),
.CK(clk),
.Q(net4757),
.QN(net4756)
);

OR3_X4 c4479(
.A1(net4730),
.A2(net4757),
.A3(net10901),
.ZN(net4758)
);

OAI211_X4 c4480(
.A(net4754),
.B(net4758),
.C1(net4755),
.C2(net4665),
.ZN(net4759)
);

OAI211_X1 c4481(
.A(net4752),
.B(net4743),
.C1(net4755),
.C2(net11037),
.ZN(net4760)
);

NOR2_X2 c4482(
.A1(net3670),
.A2(net2822),
.ZN(net4761)
);

XOR2_X2 c4483(
.A(net3666),
.B(net819),
.Z(net4762)
);

XNOR2_X1 c4484(
.A(net3697),
.B(net3855),
.ZN(net4763)
);

OR2_X4 c4485(
.A1(net720),
.A2(net1840),
.ZN(net4764)
);

AND3_X2 c4486(
.A1(net4628),
.A2(net863),
.A3(net4756),
.ZN(net4765)
);

OR2_X1 c4487(
.A1(net2719),
.A2(net3849),
.ZN(net4766)
);

NOR3_X1 c4488(
.A1(net3809),
.A2(net3849),
.A3(net4732),
.ZN(net4767)
);

XNOR2_X2 c4489(
.A(net4716),
.B(net2892),
.ZN(net4768)
);

OR3_X2 c4490(
.A1(net3825),
.A2(net3809),
.A3(net4592),
.ZN(net4769)
);

DFFRS_X2 c4491(
.D(net2829),
.RN(net3856),
.SN(net3751),
.CK(clk),
.Q(net4771),
.QN(net4770)
);

OAI21_X2 c4492(
.A(net3856),
.B1(net4757),
.B2(net2849),
.ZN(net4772)
);

INV_X32 c4493(
.A(net9711),
.ZN(net4773)
);

OAI21_X1 c4494(
.A(net3671),
.B1(net2881),
.B2(net3697),
.ZN(net4774)
);

AND2_X4 c4495(
.A1(net863),
.A2(net3781),
.ZN(net4775)
);

AND2_X1 c4496(
.A1(net2855),
.A2(net2880),
.ZN(net4776)
);

NAND2_X1 c4497(
.A1(net3799),
.A2(net2855),
.ZN(net4777)
);

AOI21_X2 c4498(
.A(net4525),
.B1(net3826),
.B2(net10778),
.ZN(net4778)
);

AOI21_X1 c4499(
.A(net3858),
.B1(net3840),
.B2(net879),
.ZN(net4779)
);

AOI21_X4 c4500(
.A(net3727),
.B1(net4775),
.B2(net4716),
.ZN(net4780)
);

NAND2_X2 c4501(
.A1(net4707),
.A2(net3820),
.ZN(net4781)
);

NAND2_X4 c4502(
.A1(net4592),
.A2(net11070),
.ZN(net4782)
);

INV_X4 c4503(
.A(net10429),
.ZN(net4783)
);

AND3_X1 c4504(
.A1(net3802),
.A2(net3727),
.A3(net3846),
.ZN(net4784)
);

NAND3_X1 c4505(
.A1(net2817),
.A2(net3874),
.A3(net3789),
.ZN(net4785)
);

DFFR_X2 c4506(
.D(net4666),
.RN(net3751),
.CK(clk),
.Q(net4787),
.QN(net4786)
);

NOR3_X4 c4507(
.A1(net2880),
.A2(out1),
.A3(net4392),
.ZN(net4788)
);

NOR4_X4 c4508(
.A1(net4773),
.A2(net1802),
.A3(net785),
.A4(net3862),
.ZN(net4789)
);

NOR3_X2 c4509(
.A1(net785),
.A2(net4770),
.A3(net3789),
.ZN(net4790)
);

SDFF_X1 c4510(
.D(net3794),
.SE(net3793),
.SI(net4592),
.CK(clk),
.Q(net4792),
.QN(net4791)
);

AND3_X4 c4511(
.A1(net3851),
.A2(net3870),
.A3(net3834),
.ZN(net4793)
);

AND2_X2 c4512(
.A1(net917),
.A2(net3844),
.ZN(net4794)
);

SDFF_X2 c4513(
.D(net2877),
.SE(net4763),
.SI(net2892),
.CK(clk),
.Q(net4796),
.QN(net4795)
);

NAND3_X2 c4514(
.A1(net3781),
.A2(net4775),
.A3(net785),
.ZN(net4797)
);

NOR4_X2 c4515(
.A1(net4732),
.A2(net4777),
.A3(net3878),
.A4(net4795),
.ZN(net4798)
);

OR3_X1 c4516(
.A1(net3860),
.A2(net2848),
.A3(net3697),
.ZN(net4799)
);

XOR2_X1 c4517(
.A(net3768),
.B(net4796),
.Z(net4800)
);

NOR2_X1 c4518(
.A1(net4785),
.A2(net4762),
.ZN(net4801)
);

OR2_X2 c4519(
.A1(net4790),
.A2(net10846),
.ZN(net4802)
);

SDFFR_X1 c4520(
.D(net4761),
.RN(net1911),
.SE(net4716),
.SI(net2894),
.CK(clk),
.Q(net4804),
.QN(net4803)
);

MUX2_X1 c4521(
.A(net1860),
.B(net4802),
.S(net3850),
.Z(net4805)
);

AOI221_X1 c4522(
.A(net3760),
.B1(net4732),
.B2(net4775),
.C1(net4803),
.C2(net2751),
.ZN(net4806)
);

OAI21_X4 c4523(
.A(net2887),
.B1(net2725),
.B2(net4790),
.ZN(net4807)
);

MUX2_X2 c4524(
.A(net3669),
.B(net2751),
.S(net10596),
.Z(net4808)
);

NAND3_X4 c4525(
.A1(net3834),
.A2(net3860),
.A3(net2854),
.ZN(net4809)
);

OR3_X4 c4526(
.A1(net4790),
.A2(net4805),
.A3(net3837),
.ZN(net4810)
);

DFFRS_X1 c4527(
.D(net3864),
.RN(net4525),
.SN(net879),
.CK(clk),
.Q(net4812),
.QN(net4811)
);

NOR2_X4 c4528(
.A1(net3840),
.A2(net4796),
.ZN(net4813)
);

INV_X1 c4529(
.A(net9710),
.ZN(net4814)
);

AND3_X2 c4530(
.A1(net4767),
.A2(net3811),
.A3(net4539),
.ZN(net4815)
);

OAI222_X1 c4531(
.A1(net3793),
.A2(net3814),
.B1(net4795),
.B2(net3834),
.C1(net3794),
.C2(net3849),
.ZN(net4816)
);

NOR2_X2 c4532(
.A1(net4787),
.A2(net1911),
.ZN(net4817)
);

XOR2_X2 c4533(
.A(net1851),
.B(net2777),
.Z(net4818)
);

XNOR2_X1 c4534(
.A(net10739),
.B(net11535),
.ZN(net4819)
);

OR2_X4 c4535(
.A1(net4092),
.A2(net4813),
.ZN(net4820)
);

DFFRS_X2 c4536(
.D(net3665),
.RN(net4793),
.SN(net2831),
.CK(clk),
.Q(net4822),
.QN(net4821)
);

OR2_X1 c4537(
.A1(net3669),
.A2(net4822),
.ZN(net4823)
);

NOR3_X1 c4538(
.A1(net3718),
.A2(net3871),
.A3(net720),
.ZN(net4824)
);

OR3_X2 c4539(
.A1(net3826),
.A2(net4769),
.A3(net4819),
.ZN(net4825)
);

OAI21_X2 c4540(
.A(net3788),
.B1(net4819),
.B2(net4781),
.ZN(net4826)
);

OAI21_X1 c4541(
.A(net4794),
.B1(net4771),
.B2(net11534),
.ZN(net4827)
);

AOI21_X2 c4542(
.A(net3863),
.B1(net4796),
.B2(net4804),
.ZN(net4828)
);

OAI222_X4 c4543(
.A1(net2831),
.A2(net4704),
.B1(net4818),
.B2(net4803),
.C1(net2829),
.C2(net4819),
.ZN(net4829)
);

SDFF_X1 c4544(
.D(net4813),
.SE(net2894),
.SI(net4795),
.CK(clk),
.Q(net4831),
.QN(net4830)
);

AOI21_X1 c4545(
.A(net4782),
.B1(net4824),
.B2(net4786),
.ZN(net4832)
);

AOI21_X4 c4546(
.A(net4790),
.B1(net11023),
.B2(net11535),
.ZN(net4833)
);

AND3_X1 c4547(
.A1(net3821),
.A2(net4783),
.A3(net819),
.ZN(net4834)
);

NAND3_X1 c4548(
.A1(net4820),
.A2(net4834),
.A3(net11536),
.ZN(net4835)
);

NOR3_X4 c4549(
.A1(net3418),
.A2(net4771),
.A3(net840),
.ZN(net4836)
);

NOR3_X2 c4550(
.A1(net4765),
.A2(net4831),
.A3(net11024),
.ZN(net4837)
);

AND3_X4 c4551(
.A1(net4768),
.A2(net4797),
.A3(net4821),
.ZN(net4838)
);

SDFF_X2 c4552(
.D(net3830),
.SE(net3794),
.SI(net3864),
.CK(clk),
.Q(net4840),
.QN(net4839)
);

DFFRS_X1 c4553(
.D(net1868),
.RN(net4822),
.SN(net4819),
.CK(clk),
.Q(net4842),
.QN(net4841)
);

DFFRS_X2 c4554(
.D(net4828),
.RN(net4837),
.SN(net10595),
.CK(clk),
.Q(net4844),
.QN(net4843)
);

SDFF_X1 c4555(
.D(net2881),
.SE(net2894),
.SI(net3878),
.CK(clk),
.Q(net4846),
.QN(net4845)
);

NAND3_X2 c4556(
.A1(net4775),
.A2(net4814),
.A3(net4811),
.ZN(net4847)
);

OR3_X1 c4557(
.A1(net4807),
.A2(net10707),
.A3(net11071),
.ZN(net4848)
);

OAI222_X2 c4558(
.A1(net1903),
.A2(net4842),
.B1(net4818),
.B2(net4819),
.C1(net3849),
.C2(net3818),
.ZN(net4849)
);

MUX2_X1 c4559(
.A(net819),
.B(net4813),
.S(net4845),
.Z(net4850)
);

SDFF_X2 c4560(
.D(net4806),
.SE(net4848),
.SI(net4821),
.CK(clk),
.Q(net4852),
.QN(net4851)
);

OAI21_X4 c4561(
.A(net4852),
.B1(net4835),
.B2(net4846),
.ZN(net4853)
);

MUX2_X2 c4562(
.A(net4789),
.B(net4841),
.S(net10935),
.Z(net4854)
);

NAND3_X4 c4563(
.A1(net4854),
.A2(net4851),
.A3(net3810),
.ZN(net4855)
);

OR3_X4 c4564(
.A1(net3751),
.A2(net4853),
.A3(net10811),
.ZN(net4856)
);

INV_X2 c4565(
.A(net3885),
.ZN(net4857)
);

INV_X8 c4566(
.A(net3960),
.ZN(net4858)
);

INV_X16 c4567(
.A(net3914),
.ZN(net4859)
);

INV_X32 c4568(
.A(net3906),
.ZN(net4860)
);

XNOR2_X2 c4569(
.A(net1988),
.B(net3964),
.ZN(net4861)
);

INV_X4 c4570(
.A(net3903),
.ZN(net4862)
);

INV_X1 c4571(
.A(net1016),
.ZN(net4863)
);

INV_X2 c4572(
.A(net1990),
.ZN(net4864)
);

AND2_X4 c4573(
.A1(net1915),
.A2(in24),
.ZN(net4865)
);

INV_X8 c4574(
.A(net1021),
.ZN(net4866)
);

INV_X16 c4575(
.A(net3924),
.ZN(net4867)
);

INV_X32 c4576(
.A(net3964),
.ZN(net4868)
);

INV_X4 c4577(
.A(net3954),
.ZN(net4869)
);

INV_X1 c4578(
.A(net1932),
.ZN(net4870)
);

INV_X2 c4579(
.A(in7),
.ZN(net4871)
);

INV_X8 c4580(
.A(net3902),
.ZN(net4872)
);

INV_X16 c4581(
.A(net4865),
.ZN(net4873)
);

INV_X32 c4582(
.A(net3934),
.ZN(net4874)
);

AND2_X1 c4583(
.A1(net3911),
.A2(net3954),
.ZN(net4875)
);

INV_X4 c4584(
.A(net3942),
.ZN(net4876)
);

INV_X1 c4585(
.A(net1961),
.ZN(net4877)
);

INV_X2 c4586(
.A(net2963),
.ZN(net4878)
);

INV_X8 c4587(
.A(net3911),
.ZN(net4879)
);

NAND2_X1 c4588(
.A1(net4867),
.A2(net4879),
.ZN(net4880)
);

INV_X16 c4589(
.A(net2942),
.ZN(net4881)
);

INV_X32 c4590(
.A(net4875),
.ZN(net4882)
);

INV_X4 c4591(
.A(net4873),
.ZN(net4883)
);

NAND2_X2 c4592(
.A1(in24),
.A2(net3910),
.ZN(net4884)
);

INV_X1 c4593(
.A(net4858),
.ZN(net4885)
);

NAND2_X4 c4594(
.A1(net4859),
.A2(net4883),
.ZN(net4886)
);

INV_X2 c4595(
.A(net3914),
.ZN(net4887)
);

AND2_X2 c4596(
.A1(net4880),
.A2(net2924),
.ZN(net4888)
);

INV_X8 c4597(
.A(net4885),
.ZN(net4889)
);

XOR2_X1 c4598(
.A(net4882),
.B(net3969),
.Z(net4890)
);

NOR2_X1 c4599(
.A1(net4876),
.A2(net4881),
.ZN(net4891)
);

AND3_X2 c4600(
.A1(net4883),
.A2(net4884),
.A3(net4881),
.ZN(net4892)
);

INV_X16 c4601(
.A(net9648),
.ZN(net4893)
);

INV_X32 c4602(
.A(net3920),
.ZN(net4894)
);

OR2_X2 c4603(
.A1(net4874),
.A2(net4886),
.ZN(net4895)
);

NOR2_X4 c4604(
.A1(net4881),
.A2(net4868),
.ZN(net4896)
);

INV_X4 c4605(
.A(net4884),
.ZN(net4897)
);

NOR3_X1 c4606(
.A1(net4870),
.A2(net4873),
.A3(net4892),
.ZN(net4898)
);

NOR2_X2 c4607(
.A1(net2942),
.A2(net4896),
.ZN(net4899)
);

OR3_X2 c4608(
.A1(net4887),
.A2(net3933),
.A3(net4864),
.ZN(net4900)
);

OAI21_X2 c4609(
.A(net4876),
.B1(net4879),
.B2(net4887),
.ZN(net4901)
);

XOR2_X2 c4610(
.A(net4892),
.B(net4865),
.Z(net4902)
);

INV_X1 c4611(
.A(net2980),
.ZN(net4903)
);

DFFS_X1 c4612(
.D(net4890),
.SN(net4900),
.CK(clk),
.Q(net4905),
.QN(net4904)
);

INV_X2 c4613(
.A(net4889),
.ZN(net4906)
);

XNOR2_X1 c4614(
.A(net4895),
.B(net4889),
.ZN(net4907)
);

OR2_X4 c4615(
.A1(net4885),
.A2(net4886),
.ZN(net4908)
);

OR2_X1 c4616(
.A1(net4900),
.A2(net4859),
.ZN(net4909)
);

XNOR2_X2 c4617(
.A(net4906),
.B(net4894),
.ZN(net4910)
);

INV_X8 c4618(
.A(net9649),
.ZN(net4911)
);

AND2_X4 c4619(
.A1(net4858),
.A2(net3964),
.ZN(net4912)
);

AND2_X1 c4620(
.A1(net4912),
.A2(net4897),
.ZN(net4913)
);

NAND2_X1 c4621(
.A1(net4860),
.A2(net3959),
.ZN(net4914)
);

NAND2_X2 c4622(
.A1(net4901),
.A2(net3960),
.ZN(net4915)
);

NAND2_X4 c4623(
.A1(net4892),
.A2(net4915),
.ZN(net4916)
);

AND2_X2 c4624(
.A1(net3933),
.A2(net4916),
.ZN(net4917)
);

XOR2_X1 c4625(
.A(net4875),
.B(net4878),
.Z(net4918)
);

OAI21_X1 c4626(
.A(net4897),
.B1(net4861),
.B2(net4876),
.ZN(net4919)
);

AOI21_X2 c4627(
.A(net4911),
.B1(net3942),
.B2(net4919),
.ZN(net4920)
);

NOR2_X1 c4628(
.A1(net4917),
.A2(net4918),
.ZN(net4921)
);

OR2_X2 c4629(
.A1(net3888),
.A2(net4887),
.ZN(net4922)
);

NOR2_X4 c4630(
.A1(net4914),
.A2(net4915),
.ZN(net4923)
);

AOI21_X1 c4631(
.A(net4867),
.B1(net4909),
.B2(net10665),
.ZN(net4924)
);

DFFS_X2 c4632(
.D(net3934),
.SN(net4922),
.CK(clk),
.Q(net4926),
.QN(net4925)
);

AOI222_X1 c4633(
.A1(net4912),
.A2(net4879),
.B1(net4917),
.B2(net4925),
.C1(net4902),
.C2(net3904),
.ZN(net4927)
);

SDFFR_X2 c4634(
.D(net4857),
.RN(net4893),
.SE(net4922),
.SI(net3955),
.CK(clk),
.Q(net4929),
.QN(net4928)
);

AOI21_X4 c4635(
.A(net4926),
.B1(net4899),
.B2(net4881),
.ZN(net4930)
);

AND3_X1 c4636(
.A1(net4915),
.A2(net4924),
.A3(net4891),
.ZN(net4931)
);

NOR2_X2 c4637(
.A1(net4893),
.A2(net4923),
.ZN(net4932)
);

XOR2_X2 c4638(
.A(net4925),
.B(net10664),
.Z(net4933)
);

AOI211_X4 c4639(
.A(net4868),
.B(net4906),
.C1(net4876),
.C2(net3902),
.ZN(net4934)
);

XNOR2_X1 c4640(
.A(net4934),
.B(net3909),
.ZN(net4935)
);

SDFFS_X1 c4641(
.D(net4922),
.SE(net4932),
.SI(net4895),
.SN(net4935),
.CK(clk),
.Q(net4937),
.QN(net4936)
);

AOI222_X4 c4642(
.A1(net4931),
.A2(net4916),
.B1(net4936),
.B2(net4874),
.C1(net4909),
.C2(net3904),
.ZN(net4938)
);

OR2_X4 c4643(
.A1(net4919),
.A2(net4915),
.ZN(net4939)
);

OR2_X1 c4644(
.A1(net4924),
.A2(net4923),
.ZN(net4940)
);

DFFRS_X1 c4645(
.D(net4934),
.RN(net4940),
.SN(net11539),
.CK(clk),
.Q(net4942),
.QN(net4941)
);

DFFRS_X2 c4646(
.D(net4940),
.RN(net4928),
.SN(net11538),
.CK(clk),
.Q(net4944),
.QN(net4943)
);

SDFFRS_X1 c4647(
.D(net4939),
.RN(net4907),
.SE(net4940),
.SI(net4935),
.SN(net4866),
.CK(clk),
.Q(net4946),
.QN(net4945)
);

XNOR2_X2 c4648(
.A(net3987),
.B(net3003),
.ZN(net4947)
);

NAND3_X1 c4649(
.A1(net4019),
.A2(net4898),
.A3(net4886),
.ZN(net4948)
);

INV_X16 c4650(
.A(net4023),
.ZN(net4949)
);

NOR3_X4 c4651(
.A1(net2058),
.A2(net2924),
.A3(net3987),
.ZN(net4950)
);

INV_X32 c4652(
.A(net4886),
.ZN(net4951)
);

AND2_X4 c4653(
.A1(net3973),
.A2(net3975),
.ZN(net4952)
);

INV_X4 c4654(
.A(net4000),
.ZN(net4953)
);

INV_X1 c4655(
.A(net2096),
.ZN(net4954)
);

INV_X2 c4656(
.A(net10468),
.ZN(net4955)
);

INV_X8 c4657(
.A(net4954),
.ZN(net4956)
);

INV_X16 c4658(
.A(net4951),
.ZN(net4957)
);

INV_X32 c4659(
.A(net9778),
.ZN(net4958)
);

AND2_X1 c4660(
.A1(net4880),
.A2(net3909),
.ZN(net4959)
);

INV_X4 c4661(
.A(net3882),
.ZN(net4960)
);

NAND2_X1 c4662(
.A1(net3048),
.A2(net4898),
.ZN(net4961)
);

INV_X1 c4663(
.A(net9815),
.ZN(net4962)
);

INV_X2 c4664(
.A(net4003),
.ZN(net4963)
);

INV_X8 c4665(
.A(net4955),
.ZN(net4964)
);

NAND2_X2 c4666(
.A1(net3003),
.A2(net3079),
.ZN(net4965)
);

INV_X16 c4667(
.A(net4956),
.ZN(net4966)
);

DFFR_X1 c4668(
.D(net4890),
.RN(net4891),
.CK(clk),
.Q(net4968),
.QN(net4967)
);

INV_X32 c4669(
.A(net11020),
.ZN(net4969)
);

SDFF_X1 c4670(
.D(net4950),
.SE(net4966),
.SI(net4963),
.CK(clk),
.Q(net4971),
.QN(net4970)
);

INV_X4 c4671(
.A(net4021),
.ZN(net4972)
);

INV_X1 c4672(
.A(net4933),
.ZN(net4973)
);

INV_X2 c4673(
.A(net4959),
.ZN(net4974)
);

NAND2_X4 c4674(
.A1(net4899),
.A2(net4916),
.ZN(net4975)
);

SDFF_X2 c4675(
.D(net4916),
.SE(net2081),
.SI(net4948),
.CK(clk),
.Q(net4977),
.QN(net4976)
);

INV_X8 c4676(
.A(net2980),
.ZN(net4978)
);

AND2_X2 c4677(
.A1(net4972),
.A2(net4969),
.ZN(net4979)
);

XOR2_X1 c4678(
.A(net4944),
.B(net4916),
.Z(net4980)
);

INV_X16 c4679(
.A(net4960),
.ZN(net4981)
);

NOR2_X1 c4680(
.A1(net2924),
.A2(net3948),
.ZN(net4982)
);

INV_X32 c4681(
.A(net1932),
.ZN(net4983)
);

OR2_X2 c4682(
.A1(net4942),
.A2(net3993),
.ZN(net4984)
);

NOR2_X4 c4683(
.A1(net4971),
.A2(net4968),
.ZN(net4985)
);

NOR2_X2 c4684(
.A1(net4985),
.A2(net2096),
.ZN(net4986)
);

INV_X4 c4685(
.A(net4926),
.ZN(net4987)
);

INV_X1 c4686(
.A(net4981),
.ZN(net4988)
);

INV_X2 c4687(
.A(net4979),
.ZN(net4989)
);

INV_X8 c4688(
.A(net2066),
.ZN(net4990)
);

XOR2_X2 c4689(
.A(net4964),
.B(net4986),
.Z(net4991)
);

DFFR_X2 c4690(
.D(net4961),
.RN(net4984),
.CK(clk),
.Q(net4993),
.QN(net4992)
);

XNOR2_X1 c4691(
.A(net4991),
.B(net4866),
.ZN(net4994)
);

OR2_X4 c4692(
.A1(net4947),
.A2(net4994),
.ZN(net4995)
);

INV_X16 c4693(
.A(net10264),
.ZN(net4996)
);

INV_X32 c4694(
.A(net4879),
.ZN(net4997)
);

NOR3_X2 c4695(
.A1(net4986),
.A2(net4963),
.A3(net4970),
.ZN(net4998)
);

DFFRS_X1 c4696(
.D(net4989),
.RN(net3038),
.SN(net4974),
.CK(clk),
.Q(net5000),
.QN(net4999)
);

AND3_X4 c4697(
.A1(net3079),
.A2(net4923),
.A3(net4984),
.ZN(net5001)
);

INV_X4 c4698(
.A(net9778),
.ZN(net5002)
);

OR2_X1 c4699(
.A1(net4881),
.A2(net10903),
.ZN(net5003)
);

DFFS_X1 c4700(
.D(net4990),
.SN(net4943),
.CK(clk),
.Q(net5005),
.QN(net5004)
);

INV_X1 c4701(
.A(net10593),
.ZN(net5006)
);

XNOR2_X2 c4702(
.A(net4948),
.B(net4866),
.ZN(net5007)
);

INV_X2 c4703(
.A(net10240),
.ZN(net5008)
);

INV_X8 c4704(
.A(net4998),
.ZN(net5009)
);

AND2_X4 c4705(
.A1(net4994),
.A2(net4995),
.ZN(net5010)
);

NAND3_X2 c4706(
.A1(net5008),
.A2(net4959),
.A3(net4990),
.ZN(net5011)
);

AND2_X1 c4707(
.A1(net4987),
.A2(net3948),
.ZN(net5012)
);

NAND2_X1 c4708(
.A1(net4971),
.A2(net10798),
.ZN(net5013)
);

INV_X16 c4709(
.A(net4978),
.ZN(net5014)
);

INV_X32 c4710(
.A(net5014),
.ZN(net5015)
);

NAND2_X2 c4711(
.A1(net4866),
.A2(net5003),
.ZN(net5016)
);

OR3_X1 c4712(
.A1(net5013),
.A2(net5005),
.A3(net4969),
.ZN(net5017)
);

INV_X4 c4713(
.A(net10055),
.ZN(net5018)
);

NAND2_X4 c4714(
.A1(net4983),
.A2(net4973),
.ZN(net5019)
);

AND2_X2 c4715(
.A1(net5016),
.A2(net4994),
.ZN(net5020)
);

INV_X1 c4716(
.A(net11020),
.ZN(net5021)
);

XOR2_X1 c4717(
.A(net5003),
.B(net4897),
.Z(net5022)
);

MUX2_X1 c4718(
.A(net5018),
.B(net4001),
.S(net11103),
.Z(net5023)
);

NOR2_X1 c4719(
.A1(net5022),
.A2(net5015),
.ZN(net5024)
);

OR2_X2 c4720(
.A1(net5015),
.A2(net5000),
.ZN(net5025)
);

NOR2_X4 c4721(
.A1(net5019),
.A2(net4972),
.ZN(net5026)
);

NOR2_X2 c4722(
.A1(net4966),
.A2(net4024),
.ZN(net5027)
);

OAI21_X4 c4723(
.A(net3885),
.B1(net4994),
.B2(net5018),
.ZN(net5028)
);

OAI33_X1 c4724(
.A1(net4985),
.A2(net5028),
.A3(net4954),
.B1(net4999),
.B2(net3038),
.B3(net4994),
.ZN(net5029)
);

XOR2_X2 c4725(
.A(net5026),
.B(net5015),
.Z(net5030)
);

DFFRS_X2 c4726(
.D(net5020),
.RN(net5013),
.SN(net3902),
.CK(clk),
.Q(net5032),
.QN(net5031)
);

XNOR2_X1 c4727(
.A(net5030),
.B(net5004),
.ZN(net5033)
);

MUX2_X2 c4728(
.A(net5027),
.B(net4941),
.S(net11019),
.Z(net5034)
);

AOI222_X2 c4729(
.A1(net5027),
.A2(net5033),
.B1(net4999),
.B2(net3981),
.C1(net4964),
.C2(net10594),
.ZN(net5035)
);

SDFF_X1 c4730(
.D(net4891),
.SE(net5033),
.SI(net5030),
.CK(clk),
.Q(net5037),
.QN(net5036)
);

OR2_X4 c4731(
.A1(net3156),
.A2(net1951),
.ZN(net5038)
);

OR2_X1 c4732(
.A1(net2130),
.A2(net4996),
.ZN(net5039)
);

XNOR2_X2 c4733(
.A(net4143),
.B(net5039),
.ZN(net5040)
);

AND2_X4 c4734(
.A1(net3909),
.A2(net11504),
.ZN(net5041)
);

AND2_X1 c4735(
.A1(net4952),
.A2(net4014),
.ZN(net5042)
);

INV_X2 c4736(
.A(net2061),
.ZN(net5043)
);

INV_X8 c4737(
.A(net2928),
.ZN(net5044)
);

INV_X16 c4738(
.A(net4864),
.ZN(net5045)
);

INV_X32 c4739(
.A(net4033),
.ZN(net5046)
);

INV_X4 c4740(
.A(net10480),
.ZN(net5047)
);

INV_X1 c4741(
.A(net3100),
.ZN(net5048)
);

NAND2_X1 c4742(
.A1(net5041),
.A2(net4963),
.ZN(net5049)
);

INV_X2 c4743(
.A(net5039),
.ZN(net5050)
);

NAND2_X2 c4744(
.A1(net5045),
.A2(net4976),
.ZN(net5051)
);

NAND2_X4 c4745(
.A1(net4001),
.A2(net11371),
.ZN(net5052)
);

AND2_X2 c4746(
.A1(net5043),
.A2(net2130),
.ZN(net5053)
);

INV_X8 c4747(
.A(net10002),
.ZN(net5054)
);

INV_X16 c4748(
.A(net4117),
.ZN(net5055)
);

INV_X32 c4749(
.A(net5051),
.ZN(net5056)
);

INV_X4 c4750(
.A(net10830),
.ZN(net5057)
);

XOR2_X1 c4751(
.A(net2161),
.B(net4067),
.Z(net5058)
);

INV_X1 c4752(
.A(net3987),
.ZN(net5059)
);

INV_X2 c4753(
.A(net5058),
.ZN(net5060)
);

NAND3_X4 c4754(
.A1(net4861),
.A2(net5059),
.A3(net4024),
.ZN(net5061)
);

NOR2_X1 c4755(
.A1(net5049),
.A2(net5059),
.ZN(net5062)
);

INV_X8 c4756(
.A(net9769),
.ZN(net5063)
);

INV_X16 c4757(
.A(net5040),
.ZN(net5064)
);

INV_X32 c4758(
.A(net11079),
.ZN(net5065)
);

INV_X4 c4759(
.A(net5060),
.ZN(net5066)
);

OR2_X2 c4760(
.A1(net4086),
.A2(net5059),
.ZN(net5067)
);

INV_X1 c4761(
.A(net5040),
.ZN(net5068)
);

NOR2_X4 c4762(
.A1(net4898),
.A2(net5066),
.ZN(net5069)
);

INV_X2 c4763(
.A(net2963),
.ZN(net5070)
);

INV_X8 c4764(
.A(net9769),
.ZN(net5071)
);

INV_X16 c4765(
.A(net10141),
.ZN(net5072)
);

OR3_X4 c4766(
.A1(net5050),
.A2(net5009),
.A3(net5070),
.ZN(net5073)
);

INV_X32 c4767(
.A(net5070),
.ZN(net5074)
);

NOR2_X2 c4768(
.A1(net5074),
.A2(net5066),
.ZN(net5075)
);

AND3_X2 c4769(
.A1(net5059),
.A2(net5058),
.A3(net4902),
.ZN(net5076)
);

SDFF_X2 c4770(
.D(net4001),
.SE(net5061),
.SI(net4119),
.CK(clk),
.Q(net5078),
.QN(net5077)
);

XOR2_X2 c4771(
.A(net4127),
.B(net11177),
.Z(net5079)
);

OAI221_X1 c4772(
.A(net4977),
.B1(net5058),
.B2(net3969),
.C1(net5033),
.C2(net5060),
.ZN(net5080)
);

XNOR2_X1 c4773(
.A(net5072),
.B(net4970),
.ZN(net5081)
);

OR2_X4 c4774(
.A1(net5063),
.A2(net5036),
.ZN(net5082)
);

INV_X4 c4775(
.A(net10472),
.ZN(net5083)
);

OR2_X1 c4776(
.A1(net5067),
.A2(net5070),
.ZN(net5084)
);

NOR3_X1 c4777(
.A1(net4933),
.A2(net4107),
.A3(net5057),
.ZN(net5085)
);

INV_X1 c4778(
.A(net4144),
.ZN(net5086)
);

XNOR2_X2 c4779(
.A(net5068),
.B(net5060),
.ZN(net5087)
);

OR3_X2 c4780(
.A1(net5075),
.A2(net4122),
.A3(net4959),
.ZN(net5088)
);

AND2_X4 c4781(
.A1(net4119),
.A2(net4973),
.ZN(net5089)
);

AND2_X1 c4782(
.A1(net5065),
.A2(net4122),
.ZN(net5090)
);

INV_X2 c4783(
.A(net9875),
.ZN(net5091)
);

DFFRS_X1 c4784(
.D(net5075),
.RN(net3120),
.SN(net10559),
.CK(clk),
.Q(net5093),
.QN(net5092)
);

INV_X8 c4785(
.A(net5090),
.ZN(net5094)
);

INV_X16 c4786(
.A(net5084),
.ZN(net5095)
);

OAI221_X4 c4787(
.A(net5095),
.B1(net5060),
.B2(net5075),
.C1(net5070),
.C2(net4140),
.ZN(net5096)
);

INV_X32 c4788(
.A(net9874),
.ZN(net5097)
);

OAI21_X2 c4789(
.A(net5085),
.B1(net4952),
.B2(net5077),
.ZN(net5098)
);

OAI221_X2 c4790(
.A(net5060),
.B1(net3165),
.B2(net5053),
.C1(net3100),
.C2(net5057),
.ZN(net5099)
);

INV_X4 c4791(
.A(net3120),
.ZN(net5100)
);

DFFRS_X2 c4792(
.D(net4958),
.RN(net5092),
.SN(net5094),
.CK(clk),
.Q(net5102),
.QN(net5101)
);

INV_X1 c4793(
.A(net5054),
.ZN(net5103)
);

INV_X2 c4794(
.A(net5097),
.ZN(net5104)
);

INV_X8 c4795(
.A(net5043),
.ZN(net5105)
);

INV_X16 c4796(
.A(net10091),
.ZN(net5106)
);

INV_X32 c4797(
.A(net5106),
.ZN(net5107)
);

OAI21_X1 c4798(
.A(net3975),
.B1(net5040),
.B2(net5081),
.ZN(net5108)
);

NAND2_X1 c4799(
.A1(net5104),
.A2(net5057),
.ZN(net5109)
);

INV_X4 c4800(
.A(net9815),
.ZN(net5110)
);

INV_X1 c4801(
.A(net11223),
.ZN(net5111)
);

SDFF_X1 c4802(
.D(net5109),
.SE(net5094),
.SI(net5110),
.CK(clk),
.Q(net5113),
.QN(net5112)
);

NAND2_X2 c4803(
.A1(net5105),
.A2(net5110),
.ZN(net5114)
);

NAND2_X4 c4804(
.A1(net5108),
.A2(net5052),
.ZN(net5115)
);

AOI21_X2 c4805(
.A(net5046),
.B1(net4124),
.B2(net5107),
.ZN(net5116)
);

INV_X2 c4806(
.A(net10463),
.ZN(net5117)
);

AOI21_X1 c4807(
.A(net5055),
.B1(net5104),
.B2(net10860),
.ZN(net5118)
);

AOI21_X4 c4808(
.A(net5118),
.B1(net5070),
.B2(net4864),
.ZN(net5119)
);

AND2_X2 c4809(
.A1(net4144),
.A2(net11171),
.ZN(net5120)
);

INV_X8 c4810(
.A(net10001),
.ZN(net5121)
);

AND3_X1 c4811(
.A1(net4861),
.A2(net5120),
.A3(net10969),
.ZN(net5122)
);

INV_X16 c4812(
.A(net11222),
.ZN(net5123)
);

NAND3_X1 c4813(
.A1(net5123),
.A2(net5093),
.A3(net5109),
.ZN(net5124)
);

INV_X32 c4814(
.A(net11301),
.ZN(net5125)
);

XOR2_X1 c4815(
.A(net4193),
.B(net5083),
.Z(net5126)
);

NOR2_X1 c4816(
.A1(net4096),
.A2(net3201),
.ZN(net5127)
);

INV_X4 c4817(
.A(net4107),
.ZN(net5128)
);

OR2_X2 c4818(
.A1(net5005),
.A2(net1288),
.ZN(net5129)
);

NOR2_X4 c4819(
.A1(net5063),
.A2(net5125),
.ZN(net5130)
);

NOR2_X2 c4820(
.A1(net4208),
.A2(net4158),
.ZN(net5131)
);

XOR2_X2 c4821(
.A(net3993),
.B(net3149),
.Z(net5132)
);

INV_X1 c4822(
.A(net4191),
.ZN(net5133)
);

XNOR2_X1 c4823(
.A(net4959),
.B(net5000),
.ZN(net5134)
);

SDFF_X2 c4824(
.D(net5038),
.SE(net3259),
.SI(net3182),
.CK(clk),
.Q(net5136),
.QN(net5135)
);

INV_X2 c4825(
.A(net4122),
.ZN(net5137)
);

INV_X8 c4826(
.A(net11182),
.ZN(net5138)
);

OR2_X4 c4827(
.A1(net5133),
.A2(net11183),
.ZN(net5139)
);

OR2_X1 c4828(
.A1(net4061),
.A2(net4982),
.ZN(net5140)
);

INV_X16 c4829(
.A(net4118),
.ZN(net5141)
);

XNOR2_X2 c4830(
.A(net4147),
.B(net3913),
.ZN(net5142)
);

AND2_X4 c4831(
.A1(net5133),
.A2(net3148),
.ZN(net5143)
);

AND2_X1 c4832(
.A1(net3128),
.A2(net5006),
.ZN(net5144)
);

INV_X32 c4833(
.A(net4971),
.ZN(net5145)
);

NAND2_X1 c4834(
.A1(net258),
.A2(net5091),
.ZN(net5146)
);

NAND2_X2 c4835(
.A1(net4200),
.A2(net3108),
.ZN(net5147)
);

NAND2_X4 c4836(
.A1(net5125),
.A2(net5004),
.ZN(net5148)
);

AND2_X2 c4837(
.A1(net5147),
.A2(net5066),
.ZN(net5149)
);

XOR2_X1 c4838(
.A(net5091),
.B(net3004),
.Z(net5150)
);

NOR3_X4 c4839(
.A1(net5132),
.A2(net4140),
.A3(net5144),
.ZN(net5151)
);

INV_X4 c4840(
.A(net5111),
.ZN(net5152)
);

NOR2_X1 c4841(
.A1(net5148),
.A2(net5144),
.ZN(net5153)
);

OR2_X2 c4842(
.A1(net5134),
.A2(net3982),
.ZN(net5154)
);

NOR2_X4 c4843(
.A1(net5153),
.A2(net4091),
.ZN(net5155)
);

NOR2_X2 c4844(
.A1(net3148),
.A2(net3993),
.ZN(net5156)
);

XOR2_X2 c4845(
.A(net3969),
.B(net5053),
.Z(net5157)
);

XNOR2_X1 c4846(
.A(net5149),
.B(net2142),
.ZN(net5158)
);

NOR3_X2 c4847(
.A1(net5127),
.A2(net4194),
.A3(net5144),
.ZN(net5159)
);

INV_X1 c4848(
.A(net10487),
.ZN(net5160)
);

AND3_X4 c4849(
.A1(net3259),
.A2(net5149),
.A3(net3248),
.ZN(net5161)
);

NAND3_X2 c4850(
.A1(net5078),
.A2(net4213),
.A3(net5144),
.ZN(net5162)
);

OR2_X4 c4851(
.A1(net5138),
.A2(net5110),
.ZN(net5163)
);

OR3_X1 c4852(
.A1(net5150),
.A2(net4896),
.A3(net5126),
.ZN(net5164)
);

INV_X2 c4853(
.A(net11276),
.ZN(net5165)
);

OR2_X1 c4854(
.A1(net5127),
.A2(net11217),
.ZN(net5166)
);

INV_X8 c4855(
.A(net11192),
.ZN(net5167)
);

MUX2_X1 c4856(
.A(net5163),
.B(net5160),
.S(net4169),
.Z(net5168)
);

OAI21_X4 c4857(
.A(net4221),
.B1(net5164),
.B2(net5063),
.ZN(net5169)
);

XNOR2_X2 c4858(
.A(net4213),
.B(net5143),
.ZN(net5170)
);

AND2_X4 c4859(
.A1(net5160),
.A2(net11101),
.ZN(net5171)
);

AND2_X1 c4860(
.A1(net5170),
.A2(net5156),
.ZN(net5172)
);

NAND2_X1 c4861(
.A1(net4111),
.A2(net5107),
.ZN(net5173)
);

NAND2_X2 c4862(
.A1(net3916),
.A2(net5163),
.ZN(net5174)
);

NAND2_X4 c4863(
.A1(net5091),
.A2(net11505),
.ZN(net5175)
);

INV_X16 c4864(
.A(net11314),
.ZN(net5176)
);

INV_X32 c4865(
.A(net9764),
.ZN(net5177)
);

MUX2_X2 c4866(
.A(net5129),
.B(net5166),
.S(net5162),
.Z(net5178)
);

SDFFRS_X2 c4867(
.D(net5157),
.RN(net5078),
.SE(net4207),
.SI(net5144),
.SN(net5126),
.CK(clk),
.Q(net5180),
.QN(net5179)
);

INV_X4 c4868(
.A(net9980),
.ZN(net5181)
);

AND2_X2 c4869(
.A1(net4076),
.A2(net2153),
.ZN(net5182)
);

NAND3_X4 c4870(
.A1(net5176),
.A2(net5164),
.A3(net5111),
.ZN(net5183)
);

XOR2_X1 c4871(
.A(net5032),
.B(net5175),
.Z(net5184)
);

NOR2_X1 c4872(
.A1(net5145),
.A2(net5134),
.ZN(net5185)
);

OR2_X2 c4873(
.A1(net5006),
.A2(net5125),
.ZN(net5186)
);

NOR4_X1 c4874(
.A1(net5142),
.A2(net5175),
.A3(net5173),
.A4(net5174),
.ZN(net5187)
);

NOR2_X4 c4875(
.A1(net5163),
.A2(net5165),
.ZN(net5188)
);

OR3_X4 c4876(
.A1(net5186),
.A2(net5162),
.A3(net4208),
.ZN(net5189)
);

INV_X1 c4877(
.A(net10465),
.ZN(net5190)
);

NOR2_X2 c4878(
.A1(net5171),
.A2(net5143),
.ZN(net5191)
);

XOR2_X2 c4879(
.A(net5094),
.B(net5156),
.Z(net5192)
);

XNOR2_X1 c4880(
.A(net5134),
.B(net11239),
.ZN(net5193)
);

INV_X2 c4881(
.A(net10038),
.ZN(net5194)
);

AND3_X2 c4882(
.A1(net5165),
.A2(net5031),
.A3(net5193),
.ZN(net5195)
);

NOR3_X1 c4883(
.A1(net5152),
.A2(net5156),
.A3(net5185),
.ZN(net5196)
);

AOI211_X2 c4884(
.A(net5191),
.B(net3251),
.C1(net4155),
.C2(net5144),
.ZN(net5197)
);

OR2_X4 c4885(
.A1(net5173),
.A2(net5184),
.ZN(net5198)
);

OR3_X2 c4886(
.A1(net5140),
.A2(net5170),
.A3(net5137),
.ZN(net5199)
);

OR2_X1 c4887(
.A1(net5193),
.A2(net10911),
.ZN(net5200)
);

XNOR2_X2 c4888(
.A(net5055),
.B(net5163),
.ZN(net5201)
);

INV_X8 c4889(
.A(net9763),
.ZN(net5202)
);

OAI21_X2 c4890(
.A(net5167),
.B1(net5202),
.B2(net5195),
.ZN(net5203)
);

AOI22_X1 c4891(
.A1(net4187),
.A2(net5202),
.B1(net4194),
.B2(net11326),
.ZN(net5204)
);

AND4_X4 c4892(
.A1(net5201),
.A2(net5156),
.A3(net5133),
.A4(net5053),
.ZN(net5205)
);

NAND4_X1 c4893(
.A1(net5183),
.A2(net5137),
.A3(net4219),
.A4(net5091),
.ZN(net5206)
);

OAI21_X1 c4894(
.A(net5185),
.B1(net5190),
.B2(net11313),
.ZN(net5207)
);

AOI21_X2 c4895(
.A(net5053),
.B1(net4862),
.B2(net5195),
.ZN(net5208)
);

AOI21_X1 c4896(
.A(net5198),
.B1(net5201),
.B2(net5193),
.ZN(net5209)
);

INV_X16 c4897(
.A(net10749),
.ZN(net5210)
);

AND2_X4 c4898(
.A1(net5066),
.A2(net3327),
.ZN(net5211)
);

INV_X32 c4899(
.A(net9843),
.ZN(net5212)
);

INV_X4 c4900(
.A(net11541),
.ZN(net5213)
);

INV_X1 c4901(
.A(net9672),
.ZN(net5214)
);

AND2_X1 c4902(
.A1(net3348),
.A2(net5049),
.ZN(net5215)
);

INV_X2 c4903(
.A(net4232),
.ZN(net5216)
);

DFFS_X2 c4904(
.D(net4280),
.SN(net5160),
.CK(clk),
.Q(net5218),
.QN(net5217)
);

DFFR_X1 c4905(
.D(net5196),
.RN(net4084),
.CK(clk),
.Q(net5220),
.QN(net5219)
);

INV_X8 c4906(
.A(net9916),
.ZN(net5221)
);

NAND2_X1 c4907(
.A1(net3913),
.A2(net11540),
.ZN(net5222)
);

INV_X16 c4908(
.A(net11183),
.ZN(net5223)
);

INV_X32 c4909(
.A(net5025),
.ZN(net5224)
);

NAND2_X2 c4910(
.A1(net3252),
.A2(net5182),
.ZN(net5225)
);

NAND2_X4 c4911(
.A1(net1316),
.A2(net5025),
.ZN(net5226)
);

INV_X4 c4912(
.A(net5049),
.ZN(net5227)
);

AND2_X2 c4913(
.A1(net5169),
.A2(net5164),
.ZN(net5228)
);

XOR2_X1 c4914(
.A(net5227),
.B(net2928),
.Z(net5229)
);

NOR2_X1 c4915(
.A1(net5188),
.A2(net4251),
.ZN(net5230)
);

DFFRS_X1 c4916(
.D(net5223),
.RN(net4280),
.SN(net4277),
.CK(clk),
.Q(net5232),
.QN(net5231)
);

OR2_X2 c4917(
.A1(net4155),
.A2(net5213),
.ZN(net5233)
);

NOR2_X4 c4918(
.A1(net4963),
.A2(net3276),
.ZN(net5234)
);

NOR2_X2 c4919(
.A1(net3276),
.A2(net5234),
.ZN(net5235)
);

XOR2_X2 c4920(
.A(net4251),
.B(net5223),
.Z(net5236)
);

XNOR2_X1 c4921(
.A(net3327),
.B(net258),
.ZN(net5237)
);

INV_X1 c4922(
.A(net10389),
.ZN(net5238)
);

OR2_X4 c4923(
.A1(net4277),
.A2(net5228),
.ZN(net5239)
);

OR2_X1 c4924(
.A1(net5154),
.A2(net5235),
.ZN(net5240)
);

XNOR2_X2 c4925(
.A(net5220),
.B(net5217),
.ZN(net5241)
);

INV_X2 c4926(
.A(net5241),
.ZN(net5242)
);

AND2_X4 c4927(
.A1(net5185),
.A2(net5223),
.ZN(net5243)
);

AND2_X1 c4928(
.A1(net3317),
.A2(net1951),
.ZN(net5244)
);

INV_X8 c4929(
.A(net3235),
.ZN(net5245)
);

NAND2_X1 c4930(
.A1(net4896),
.A2(net5131),
.ZN(net5246)
);

AOI21_X4 c4931(
.A(net5044),
.B1(net5221),
.B2(net5218),
.ZN(net5247)
);

INV_X16 c4932(
.A(net3108),
.ZN(net5248)
);

INV_X32 c4933(
.A(net10497),
.ZN(net5249)
);

INV_X4 c4934(
.A(net10062),
.ZN(net5250)
);

AND3_X1 c4935(
.A1(net5182),
.A2(net2294),
.A3(net5196),
.ZN(net5251)
);

NAND2_X2 c4936(
.A1(net2277),
.A2(net5219),
.ZN(net5252)
);

NAND2_X4 c4937(
.A1(net5218),
.A2(net5225),
.ZN(net5253)
);

INV_X1 c4938(
.A(net9672),
.ZN(net5254)
);

INV_X2 c4939(
.A(net10365),
.ZN(net5255)
);

DFFRS_X2 c4940(
.D(net5233),
.RN(net5254),
.SN(net5205),
.CK(clk),
.Q(net5257),
.QN(net5256)
);

NAND3_X1 c4941(
.A1(net5143),
.A2(net5236),
.A3(net5221),
.ZN(net5258)
);

INV_X8 c4942(
.A(net4235),
.ZN(net5259)
);

AND2_X2 c4943(
.A1(net5164),
.A2(net5242),
.ZN(net5260)
);

XOR2_X1 c4944(
.A(net5214),
.B(net5243),
.Z(net5261)
);

NOR2_X1 c4945(
.A1(net5254),
.A2(net5213),
.ZN(net5262)
);

OR2_X2 c4946(
.A1(net4269),
.A2(net5230),
.ZN(net5263)
);

INV_X16 c4947(
.A(net11278),
.ZN(net5264)
);

NOR2_X4 c4948(
.A1(net5261),
.A2(net1247),
.ZN(net5265)
);

NOR2_X2 c4949(
.A1(net5257),
.A2(net5235),
.ZN(net5266)
);

INV_X32 c4950(
.A(net10246),
.ZN(net5267)
);

AOI221_X4 c4951(
.A(net5248),
.B1(net5267),
.B2(net5255),
.C1(net5233),
.C2(net3257),
.ZN(net5268)
);

NOR3_X4 c4952(
.A1(net5238),
.A2(net5166),
.A3(net5250),
.ZN(net5269)
);

OAI222_X1 c4953(
.A1(net4256),
.A2(net3317),
.B1(net4194),
.B2(net4245),
.C1(net5228),
.C2(net5234),
.ZN(net5270)
);

NOR3_X2 c4954(
.A1(net5229),
.A2(net5236),
.A3(net2294),
.ZN(net5271)
);

XOR2_X2 c4955(
.A(net1247),
.B(net5266),
.Z(net5272)
);

XNOR2_X1 c4956(
.A(net5263),
.B(net5254),
.ZN(net5273)
);

OR2_X4 c4957(
.A1(net5266),
.A2(net11040),
.ZN(net5274)
);

OR2_X1 c4958(
.A1(net5252),
.A2(net5230),
.ZN(net5275)
);

AND3_X4 c4959(
.A1(net5255),
.A2(net4267),
.A3(net5267),
.ZN(net5276)
);

NAND3_X2 c4960(
.A1(net5260),
.A2(net3235),
.A3(net11542),
.ZN(net5277)
);

INV_X4 c4961(
.A(net10392),
.ZN(net5278)
);

XNOR2_X2 c4962(
.A(net5233),
.B(net10569),
.ZN(net5279)
);

OR4_X1 c4963(
.A1(net5268),
.A2(net3317),
.A3(net5278),
.A4(net4245),
.ZN(net5280)
);

OR3_X1 c4964(
.A1(net5272),
.A2(net5233),
.A3(net11483),
.ZN(net5281)
);

MUX2_X1 c4965(
.A(net5128),
.B(net5256),
.S(net11543),
.Z(net5282)
);

OAI21_X4 c4966(
.A(net5282),
.B1(net2294),
.B2(net10768),
.ZN(net5283)
);

AND2_X4 c4967(
.A1(net5264),
.A2(net5278),
.ZN(net5284)
);

MUX2_X2 c4968(
.A(net5259),
.B(net5257),
.S(net5233),
.Z(net5285)
);

AND2_X1 c4969(
.A1(net5221),
.A2(net11386),
.ZN(net5286)
);

INV_X1 c4970(
.A(net10419),
.ZN(net5287)
);

NAND2_X1 c4971(
.A1(net5266),
.A2(net5287),
.ZN(net5288)
);

SDFF_X1 c4972(
.D(net5205),
.SE(net5268),
.SI(net3296),
.CK(clk),
.Q(net5290),
.QN(net5289)
);

NAND3_X4 c4973(
.A1(net4265),
.A2(net5290),
.A3(net10570),
.ZN(net5291)
);

OAI222_X4 c4974(
.A1(net5267),
.A2(net2277),
.B1(net5289),
.B2(net5234),
.C1(net3981),
.C2(net11386),
.ZN(net5292)
);

OR3_X4 c4975(
.A1(net5290),
.A2(net5292),
.A3(net5288),
.ZN(net5293)
);

NAND2_X2 c4976(
.A1(net5237),
.A2(net3306),
.ZN(net5294)
);

AND3_X2 c4977(
.A1(net5286),
.A2(net5290),
.A3(net11483),
.ZN(net5295)
);

OAI222_X2 c4978(
.A1(net3306),
.A2(net5284),
.B1(net5289),
.B2(net5092),
.C1(net4277),
.C2(net11542),
.ZN(net5296)
);

NOR3_X1 c4979(
.A1(net5292),
.A2(net5291),
.A3(net4090),
.ZN(net5297)
);

INV_X2 c4980(
.A(net5294),
.ZN(net5298)
);

NAND2_X4 c4981(
.A1(net5262),
.A2(net5265),
.ZN(net5299)
);

INV_X8 c4982(
.A(net2328),
.ZN(net5300)
);

AND2_X2 c4983(
.A1(net5249),
.A2(net3425),
.ZN(net5301)
);

XOR2_X1 c4984(
.A(net4263),
.B(net4392),
.Z(net5302)
);

SDFF_X2 c4985(
.D(net4363),
.SE(net5301),
.SI(net5275),
.CK(clk),
.Q(net5304),
.QN(net5303)
);

NOR2_X1 c4986(
.A1(net5291),
.A2(net4340),
.ZN(net5305)
);

INV_X16 c4987(
.A(net5265),
.ZN(net5306)
);

INV_X32 c4988(
.A(net9742),
.ZN(net5307)
);

OR2_X2 c4989(
.A1(net4258),
.A2(net4333),
.ZN(net5308)
);

INV_X4 c4990(
.A(net9742),
.ZN(net5309)
);

OR3_X2 c4991(
.A1(net5300),
.A2(net4267),
.A3(net4245),
.ZN(net5310)
);

OAI21_X2 c4992(
.A(net5305),
.B1(net5284),
.B2(net4374),
.ZN(net5311)
);

INV_X1 c4993(
.A(net11365),
.ZN(net5312)
);

INV_X2 c4994(
.A(net9826),
.ZN(net5313)
);

NOR2_X4 c4995(
.A1(net5311),
.A2(net5195),
.ZN(net5314)
);

INV_X8 c4996(
.A(net1297),
.ZN(net5315)
);

OAI21_X1 c4997(
.A(net3425),
.B1(net5298),
.B2(net5296),
.ZN(net5316)
);

NOR2_X2 c4998(
.A1(net4274),
.A2(net1412),
.ZN(net5317)
);

XOR2_X2 c4999(
.A(net5302),
.B(net4399),
.Z(net5318)
);

XNOR2_X1 c5000(
.A(net5212),
.B(net5307),
.ZN(net5319)
);

INV_X16 c5001(
.A(net5315),
.ZN(net5320)
);

OR2_X4 c5002(
.A1(net4380),
.A2(net4340),
.ZN(net5321)
);

INV_X32 c5003(
.A(net9843),
.ZN(net5322)
);

INV_X4 c5004(
.A(net5320),
.ZN(net5323)
);

OR2_X1 c5005(
.A1(net4301),
.A2(net5288),
.ZN(net5324)
);

INV_X1 c5006(
.A(net10281),
.ZN(net5325)
);

INV_X2 c5007(
.A(net5322),
.ZN(net5326)
);

AOI21_X2 c5008(
.A(net4353),
.B1(net5320),
.B2(net11421),
.ZN(net5327)
);

XNOR2_X2 c5009(
.A(net5265),
.B(net11421),
.ZN(net5328)
);

AOI21_X1 c5010(
.A(net5298),
.B1(net5309),
.B2(net3425),
.ZN(net5329)
);

AOI21_X4 c5011(
.A(net5314),
.B1(net5313),
.B2(net4374),
.ZN(net5330)
);

AND2_X4 c5012(
.A1(net5083),
.A2(net4237),
.ZN(net5331)
);

DFFRS_X1 c5013(
.D(net4237),
.RN(net5291),
.SN(net5330),
.CK(clk),
.Q(net5333),
.QN(net5332)
);

INV_X8 c5014(
.A(net5160),
.ZN(net5334)
);

INV_X16 c5015(
.A(net4381),
.ZN(net5335)
);

AND2_X1 c5016(
.A1(net5159),
.A2(net5331),
.ZN(net5336)
);

NAND2_X1 c5017(
.A1(net3411),
.A2(net5250),
.ZN(net5337)
);

INV_X32 c5018(
.A(net9853),
.ZN(net5338)
);

NAND2_X2 c5019(
.A1(net5326),
.A2(net4263),
.ZN(net5339)
);

NAND2_X4 c5020(
.A1(net5323),
.A2(net5334),
.ZN(net5340)
);

INV_X4 c5021(
.A(net10359),
.ZN(net5341)
);

AND2_X2 c5022(
.A1(net5328),
.A2(net11394),
.ZN(net5342)
);

INV_X1 c5023(
.A(net10421),
.ZN(net5343)
);

AND3_X1 c5024(
.A1(net5335),
.A2(net5331),
.A3(net5340),
.ZN(net5344)
);

NAND3_X1 c5025(
.A1(net5325),
.A2(net4340),
.A3(net4265),
.ZN(net5345)
);

INV_X2 c5026(
.A(net10208),
.ZN(net5346)
);

INV_X8 c5027(
.A(net10386),
.ZN(net5347)
);

NOR3_X4 c5028(
.A1(net5340),
.A2(net5328),
.A3(net5291),
.ZN(net5348)
);

AOI221_X2 c5029(
.A(net5330),
.B1(net4346),
.B2(net5274),
.C1(net5309),
.C2(net5307),
.ZN(net5349)
);

NOR3_X2 c5030(
.A1(net5327),
.A2(net5331),
.A3(net4346),
.ZN(net5350)
);

XOR2_X1 c5031(
.A(net3406),
.B(net4374),
.Z(net5351)
);

DFFR_X2 c5032(
.D(net2411),
.RN(net3217),
.CK(clk),
.Q(net5353),
.QN(net5352)
);

INV_X16 c5033(
.A(net11365),
.ZN(net5354)
);

NOR2_X1 c5034(
.A1(net5354),
.A2(net5200),
.ZN(net5355)
);

AND3_X4 c5035(
.A1(net4341),
.A2(net5355),
.A3(net5160),
.ZN(net5356)
);

OR2_X2 c5036(
.A1(net5338),
.A2(net3406),
.ZN(net5357)
);

NOR2_X4 c5037(
.A1(net4403),
.A2(net5340),
.ZN(net5358)
);

NOR2_X2 c5038(
.A1(net5316),
.A2(net5253),
.ZN(net5359)
);

DFFS_X1 c5039(
.D(net5301),
.SN(net5311),
.CK(clk),
.Q(net5361),
.QN(net5360)
);

NAND3_X2 c5040(
.A1(net4265),
.A2(net4399),
.A3(net11312),
.ZN(net5362)
);

XOR2_X2 c5041(
.A(net4373),
.B(net5287),
.Z(net5363)
);

OR3_X1 c5042(
.A1(net5361),
.A2(net5310),
.A3(net10970),
.ZN(net5364)
);

XNOR2_X1 c5043(
.A(net5361),
.B(net5012),
.ZN(net5365)
);

OR2_X4 c5044(
.A1(net5355),
.A2(net472),
.ZN(net5366)
);

MUX2_X1 c5045(
.A(net5363),
.B(net5362),
.S(net5083),
.Z(net5367)
);

OR2_X1 c5046(
.A1(net5365),
.A2(net5353),
.ZN(net5368)
);

XNOR2_X2 c5047(
.A(net4408),
.B(net5353),
.ZN(net5369)
);

AND2_X4 c5048(
.A1(net5319),
.A2(net5365),
.ZN(net5370)
);

INV_X32 c5049(
.A(net10280),
.ZN(net5371)
);

INV_X4 c5050(
.A(net11479),
.ZN(net5372)
);

DFFRS_X2 c5051(
.D(net5366),
.RN(net5365),
.SN(net5337),
.CK(clk),
.Q(net5374),
.QN(net5373)
);

AOI221_X1 c5052(
.A(net5203),
.B1(net5373),
.B2(net2411),
.C1(net5347),
.C2(net5321),
.ZN(net5375)
);

OAI221_X1 c5053(
.A(net4244),
.B1(net5166),
.B2(net4365),
.C1(net5347),
.C2(net3257),
.ZN(net5376)
);

OAI21_X4 c5054(
.A(net5308),
.B1(net5340),
.B2(net5365),
.ZN(net5377)
);

AND2_X1 c5055(
.A1(net5343),
.A2(net5370),
.ZN(net5378)
);

OAI221_X4 c5056(
.A(net5367),
.B1(net5378),
.B2(net5375),
.C1(net5334),
.C2(net5347),
.ZN(net5379)
);

NAND2_X1 c5057(
.A1(net5312),
.A2(net10745),
.ZN(net5380)
);

MUX2_X2 c5058(
.A(net5380),
.B(net5378),
.S(net5347),
.Z(net5381)
);

NAND3_X4 c5059(
.A1(net5341),
.A2(net5381),
.A3(net5354),
.ZN(net5382)
);

AOI222_X1 c5060(
.A1(net5346),
.A2(net5382),
.B1(net5339),
.B2(net5360),
.C1(net5332),
.C2(net5352),
.ZN(net5383)
);

NAND2_X2 c5061(
.A1(net5381),
.A2(net5382),
.ZN(net5384)
);

AOI222_X4 c5062(
.A1(net5384),
.A2(net5381),
.B1(net5382),
.B2(net4334),
.C1(net5352),
.C2(net10884),
.ZN(net5385)
);

NAND2_X4 c5063(
.A1(net4333),
.A2(net4426),
.ZN(net5386)
);

AND2_X2 c5064(
.A1(net5333),
.A2(net11348),
.ZN(net5387)
);

INV_X1 c5065(
.A(net949),
.ZN(net5388)
);

INV_X2 c5066(
.A(net4905),
.ZN(net5389)
);

INV_X8 c5067(
.A(net2490),
.ZN(net5390)
);

XOR2_X1 c5068(
.A(net4482),
.B(net5368),
.Z(net5391)
);

INV_X16 c5069(
.A(net5130),
.ZN(net5392)
);

NOR2_X1 c5070(
.A1(net4245),
.A2(net4477),
.ZN(net5393)
);

INV_X32 c5071(
.A(net4267),
.ZN(net5394)
);

INV_X4 c5072(
.A(net4982),
.ZN(net5395)
);

INV_X1 c5073(
.A(net9800),
.ZN(net5396)
);

OR2_X2 c5074(
.A1(net5331),
.A2(net4477),
.ZN(net5397)
);

NOR2_X4 c5075(
.A1(net4445),
.A2(net4267),
.ZN(net5398)
);

INV_X2 c5076(
.A(net9800),
.ZN(net5399)
);

INV_X8 c5077(
.A(net4477),
.ZN(net5400)
);

INV_X16 c5078(
.A(net5213),
.ZN(net5401)
);

INV_X32 c5079(
.A(net11460),
.ZN(net5402)
);

INV_X4 c5080(
.A(net4410),
.ZN(net5403)
);

INV_X1 c5081(
.A(net5339),
.ZN(net5404)
);

INV_X2 c5082(
.A(net5374),
.ZN(net5405)
);

INV_X8 c5083(
.A(net3436),
.ZN(net5406)
);

OR3_X4 c5084(
.A1(net5400),
.A2(net556),
.A3(net5406),
.ZN(net5407)
);

INV_X16 c5085(
.A(net5386),
.ZN(net5408)
);

NOR2_X2 c5086(
.A1(net5368),
.A2(net4472),
.ZN(net5409)
);

INV_X32 c5087(
.A(net9819),
.ZN(net5410)
);

INV_X4 c5088(
.A(net4426),
.ZN(net5411)
);

INV_X1 c5089(
.A(net5246),
.ZN(net5412)
);

SDFF_X1 c5090(
.D(net5395),
.SE(net5345),
.SI(net5275),
.CK(clk),
.Q(net5414),
.QN(net5413)
);

INV_X2 c5091(
.A(net11058),
.ZN(net5415)
);

INV_X8 c5092(
.A(net5397),
.ZN(net5416)
);

INV_X16 c5093(
.A(net10184),
.ZN(net5417)
);

OAI221_X2 c5094(
.A(net5195),
.B1(net3446),
.B2(net5414),
.C1(net5166),
.C2(net5389),
.ZN(net5418)
);

INV_X32 c5095(
.A(net4447),
.ZN(net5419)
);

XOR2_X2 c5096(
.A(net4407),
.B(net5417),
.Z(net5420)
);

OAI22_X1 c5097(
.A1(net5416),
.A2(net5406),
.B1(net5331),
.B2(net2527),
.ZN(net5421)
);

XNOR2_X1 c5098(
.A(net4337),
.B(net4445),
.ZN(net5422)
);

SDFFS_X2 c5099(
.D(net3478),
.SE(net5374),
.SI(net4476),
.SN(net5389),
.CK(clk),
.Q(net5424),
.QN(net5423)
);

OR2_X4 c5100(
.A1(net5415),
.A2(net4447),
.ZN(net5425)
);

OR2_X1 c5101(
.A1(net5345),
.A2(net4423),
.ZN(net5426)
);

INV_X4 c5102(
.A(net9856),
.ZN(net5427)
);

AND3_X2 c5103(
.A1(net5410),
.A2(net4337),
.A3(net4267),
.ZN(net5428)
);

XNOR2_X2 c5104(
.A(net1491),
.B(net5402),
.ZN(net5429)
);

INV_X1 c5105(
.A(net5372),
.ZN(net5430)
);

DFFS_X2 c5106(
.D(net5430),
.SN(net2509),
.CK(clk),
.Q(net5432),
.QN(net5431)
);

AND2_X4 c5107(
.A1(net5409),
.A2(net5428),
.ZN(net5433)
);

AND2_X1 c5108(
.A1(net5398),
.A2(net4495),
.ZN(net5434)
);

NAND2_X1 c5109(
.A1(net4446),
.A2(net5434),
.ZN(net5435)
);

INV_X2 c5110(
.A(net10269),
.ZN(net5436)
);

NAND2_X2 c5111(
.A1(net5387),
.A2(net5347),
.ZN(net5437)
);

NOR3_X1 c5112(
.A1(net5418),
.A2(net5436),
.A3(net5332),
.ZN(net5438)
);

NAND2_X4 c5113(
.A1(net5369),
.A2(net4447),
.ZN(net5439)
);

INV_X8 c5114(
.A(net10431),
.ZN(net5440)
);

SDFFR_X1 c5115(
.D(net5428),
.RN(net5333),
.SE(net5434),
.SI(net5389),
.CK(clk),
.Q(net5442),
.QN(net5441)
);

AND2_X2 c5116(
.A1(net5438),
.A2(net5304),
.ZN(net5443)
);

XOR2_X1 c5117(
.A(net5411),
.B(net5422),
.Z(net5444)
);

NOR2_X1 c5118(
.A1(net5404),
.A2(net4360),
.ZN(net5445)
);

INV_X16 c5119(
.A(net10157),
.ZN(net5446)
);

OR2_X2 c5120(
.A1(net5440),
.A2(net5445),
.ZN(net5447)
);

INV_X32 c5121(
.A(net10574),
.ZN(net5448)
);

OR3_X2 c5122(
.A1(net3397),
.A2(net5436),
.A3(net5441),
.ZN(net5449)
);

DFFR_X1 c5123(
.D(net5447),
.RN(net5434),
.CK(clk),
.Q(net5451),
.QN(net5450)
);

INV_X4 c5124(
.A(net5451),
.ZN(net5452)
);

INV_X1 c5125(
.A(net5442),
.ZN(net5453)
);

NOR2_X4 c5126(
.A1(net5436),
.A2(net4245),
.ZN(net5454)
);

NOR2_X2 c5127(
.A1(net5392),
.A2(net5303),
.ZN(net5455)
);

AND4_X2 c5128(
.A1(net5288),
.A2(net4337),
.A3(net5436),
.A4(net5373),
.ZN(net5456)
);

OAI21_X2 c5129(
.A(net5426),
.B1(net4263),
.B2(net5451),
.ZN(net5457)
);

XOR2_X2 c5130(
.A(net5457),
.B(net5448),
.Z(net5458)
);

AND4_X1 c5131(
.A1(net5175),
.A2(net2517),
.A3(net5446),
.A4(net5234),
.ZN(net5459)
);

XNOR2_X1 c5132(
.A(net5394),
.B(net5454),
.ZN(net5460)
);

INV_X2 c5133(
.A(net10401),
.ZN(net5461)
);

OAI21_X1 c5134(
.A(net4360),
.B1(net5457),
.B2(net5454),
.ZN(net5462)
);

OR2_X4 c5135(
.A1(net5461),
.A2(net5452),
.ZN(net5463)
);

SDFF_X2 c5136(
.D(net5460),
.SE(net5309),
.SI(net10573),
.CK(clk),
.Q(net5465),
.QN(net5464)
);

OR2_X1 c5137(
.A1(net5450),
.A2(net10985),
.ZN(net5466)
);

DFFR_X2 c5138(
.D(net5462),
.RN(net5424),
.CK(clk),
.Q(net5468),
.QN(net5467)
);

DFFS_X1 c5139(
.D(net5421),
.SN(net4493),
.CK(clk),
.Q(net5470),
.QN(net5469)
);

AOI21_X2 c5140(
.A(net5459),
.B1(net5468),
.B2(net4481),
.ZN(net5471)
);

INV_X8 c5141(
.A(net10428),
.ZN(net5472)
);

AOI21_X1 c5142(
.A(net5471),
.B1(net5465),
.B2(net4407),
.ZN(net5473)
);

XNOR2_X2 c5143(
.A(net5466),
.B(net5465),
.ZN(net5474)
);

INV_X16 c5144(
.A(net11228),
.ZN(net5475)
);

AND2_X4 c5145(
.A1(net5474),
.A2(net5475),
.ZN(net5476)
);

INV_X32 c5146(
.A(net5452),
.ZN(net5477)
);

INV_X4 c5147(
.A(net9734),
.ZN(net5478)
);

INV_X1 c5148(
.A(net5439),
.ZN(net5479)
);

INV_X2 c5149(
.A(net5406),
.ZN(net5480)
);

INV_X8 c5150(
.A(net10355),
.ZN(net5481)
);

AND2_X1 c5151(
.A1(net5437),
.A2(net5449),
.ZN(net5482)
);

NAND2_X1 c5152(
.A1(net4578),
.A2(net5407),
.ZN(net5483)
);

AOI21_X4 c5153(
.A(net2630),
.B1(net4483),
.B2(net4524),
.ZN(net5484)
);

INV_X16 c5154(
.A(net9734),
.ZN(net5485)
);

INV_X32 c5155(
.A(net4519),
.ZN(net5486)
);

NAND2_X2 c5156(
.A1(net4396),
.A2(net5401),
.ZN(net5487)
);

AND3_X1 c5157(
.A1(net5481),
.A2(net5309),
.A3(net5472),
.ZN(net5488)
);

INV_X4 c5158(
.A(net11266),
.ZN(net5489)
);

NAND2_X4 c5159(
.A1(net5486),
.A2(net5347),
.ZN(net5490)
);

INV_X1 c5160(
.A(net5275),
.ZN(net5491)
);

INV_X2 c5161(
.A(net9856),
.ZN(net5492)
);

AND2_X2 c5162(
.A1(net4581),
.A2(net5353),
.ZN(net5493)
);

INV_X8 c5163(
.A(net5487),
.ZN(net5494)
);

XOR2_X1 c5164(
.A(net5429),
.B(net4540),
.Z(net5495)
);

INV_X16 c5165(
.A(net10314),
.ZN(net5496)
);

INV_X32 c5166(
.A(net4472),
.ZN(net5497)
);

INV_X4 c5167(
.A(net5493),
.ZN(net5498)
);

INV_X1 c5168(
.A(net5489),
.ZN(net5499)
);

INV_X2 c5169(
.A(net3588),
.ZN(net5500)
);

INV_X8 c5170(
.A(net11312),
.ZN(net5501)
);

NOR2_X1 c5171(
.A1(net5480),
.A2(net4434),
.ZN(net5502)
);

OR2_X2 c5172(
.A1(net5501),
.A2(net10677),
.ZN(net5503)
);

INV_X16 c5173(
.A(net10153),
.ZN(net5504)
);

NAND3_X1 c5174(
.A1(net5420),
.A2(net5321),
.A3(net5502),
.ZN(net5505)
);

NOR2_X4 c5175(
.A1(net5497),
.A2(net3594),
.ZN(net5506)
);

NOR2_X2 c5176(
.A1(net5501),
.A2(net5309),
.ZN(net5507)
);

INV_X32 c5177(
.A(net3571),
.ZN(net5508)
);

XOR2_X2 c5178(
.A(net5492),
.B(net4458),
.Z(net5509)
);

DFFRS_X1 c5179(
.D(net5479),
.RN(net4534),
.SN(net5485),
.CK(clk),
.Q(net5511),
.QN(net5510)
);

XNOR2_X1 c5180(
.A(net5494),
.B(net5509),
.ZN(net5512)
);

OR2_X4 c5181(
.A1(net5495),
.A2(net5321),
.ZN(net5513)
);

OR2_X1 c5182(
.A1(net5512),
.A2(net5493),
.ZN(net5514)
);

XNOR2_X2 c5183(
.A(net4434),
.B(net5493),
.ZN(net5515)
);

AND2_X4 c5184(
.A1(net2628),
.A2(net5502),
.ZN(net5516)
);

AND2_X1 c5185(
.A1(net4220),
.A2(net5495),
.ZN(net5517)
);

NAND2_X1 c5186(
.A1(net5499),
.A2(net2582),
.ZN(net5518)
);

NAND2_X2 c5187(
.A1(net5488),
.A2(net5448),
.ZN(net5519)
);

NAND2_X4 c5188(
.A1(net5517),
.A2(net5510),
.ZN(net5520)
);

AND2_X2 c5189(
.A1(net5490),
.A2(net4504),
.ZN(net5521)
);

XOR2_X1 c5190(
.A(net5484),
.B(net5347),
.Z(net5522)
);

INV_X4 c5191(
.A(net9904),
.ZN(net5523)
);

INV_X1 c5192(
.A(net5347),
.ZN(net5524)
);

NOR2_X1 c5193(
.A1(net5475),
.A2(net5509),
.ZN(net5525)
);

NOR3_X4 c5194(
.A1(net5500),
.A2(net3598),
.A3(net3594),
.ZN(net5526)
);

INV_X2 c5195(
.A(net10406),
.ZN(net5527)
);

INV_X8 c5196(
.A(net11419),
.ZN(net5528)
);

INV_X16 c5197(
.A(net11442),
.ZN(net5529)
);

OR2_X2 c5198(
.A1(net5407),
.A2(net5515),
.ZN(net5530)
);

INV_X32 c5199(
.A(net4504),
.ZN(net5531)
);

NOR2_X4 c5200(
.A1(net5521),
.A2(net10544),
.ZN(net5532)
);

NOR2_X2 c5201(
.A1(net5529),
.A2(net5477),
.ZN(net5533)
);

XOR2_X2 c5202(
.A(net5533),
.B(net2629),
.Z(net5534)
);

NOR3_X2 c5203(
.A1(net5519),
.A2(net5449),
.A3(net5427),
.ZN(net5535)
);

XNOR2_X1 c5204(
.A(net1412),
.B(net5529),
.ZN(net5536)
);

INV_X4 c5205(
.A(net5309),
.ZN(net5537)
);

OR2_X4 c5206(
.A1(net4554),
.A2(net1562),
.ZN(net5538)
);

OR2_X1 c5207(
.A1(net5491),
.A2(net5501),
.ZN(net5539)
);

AOI22_X4 c5208(
.A1(net5267),
.A2(net5523),
.B1(net5179),
.B2(net5352),
.ZN(net5540)
);

XNOR2_X2 c5209(
.A(net5521),
.B(net5539),
.ZN(net5541)
);

INV_X1 c5210(
.A(net11416),
.ZN(net5542)
);

AND3_X4 c5211(
.A1(net5539),
.A2(net4488),
.A3(net4458),
.ZN(net5543)
);

NAND3_X2 c5212(
.A1(net5541),
.A2(net5527),
.A3(net5542),
.ZN(net5544)
);

AND2_X4 c5213(
.A1(net5543),
.A2(net5531),
.ZN(net5545)
);

AND2_X1 c5214(
.A1(net5528),
.A2(net5545),
.ZN(net5546)
);

NAND2_X1 c5215(
.A1(net5401),
.A2(net5539),
.ZN(net5547)
);

OR3_X1 c5216(
.A1(net4537),
.A2(net5508),
.A3(net3588),
.ZN(net5548)
);

NAND2_X2 c5217(
.A1(net5509),
.A2(net5486),
.ZN(net5549)
);

MUX2_X1 c5218(
.A(net5503),
.B(net5495),
.S(net10844),
.Z(net5550)
);

DFFRS_X2 c5219(
.D(net5550),
.RN(net5548),
.SN(net5547),
.CK(clk),
.Q(net5552),
.QN(net5551)
);

NAND2_X4 c5220(
.A1(net4158),
.A2(net5517),
.ZN(net5553)
);

OAI33_X1 c5221(
.A1(net5549),
.A2(net5527),
.A3(net5540),
.B1(net5509),
.B2(net4523),
.B3(net5542),
.ZN(net5554)
);

AND2_X2 c5222(
.A1(net5504),
.A2(net5542),
.ZN(net5555)
);

SDFFRS_X1 c5223(
.D(net5485),
.RN(net5506),
.SE(net5548),
.SI(net5545),
.SN(net5488),
.CK(clk),
.Q(net5557),
.QN(net5556)
);

XOR2_X1 c5224(
.A(net4483),
.B(net5550),
.Z(net5558)
);

SDFFRS_X2 c5225(
.D(net5523),
.RN(net5448),
.SE(net5550),
.SI(net5510),
.SN(net5545),
.CK(clk),
.Q(net5560),
.QN(net5559)
);

AOI221_X4 c5226(
.A(net5544),
.B1(net4504),
.B2(net5511),
.C1(net5542),
.C2(net5352),
.ZN(net5561)
);

SDFF_X1 c5227(
.D(net5558),
.SE(net5547),
.SI(net5557),
.CK(clk),
.Q(net5563),
.QN(net5562)
);

SDFF_X2 c5228(
.D(net5561),
.SE(net5525),
.SI(net5232),
.CK(clk),
.Q(net5565),
.QN(net5564)
);

NOR2_X1 c5229(
.A1(net4660),
.A2(net5506),
.ZN(net5566)
);

OR2_X2 c5230(
.A1(net4633),
.A2(net1130),
.ZN(net5567)
);

INV_X2 c5231(
.A(net10232),
.ZN(out25)
);

NOR2_X4 c5232(
.A1(net5505),
.A2(net2526),
.ZN(net5568)
);

INV_X8 c5233(
.A(net11403),
.ZN(net5569)
);

OAI21_X4 c5234(
.A(net3607),
.B1(net5513),
.B2(net5566),
.ZN(net5570)
);

INV_X16 c5235(
.A(net11175),
.ZN(net5571)
);

NOR2_X2 c5236(
.A1(net5555),
.A2(net5547),
.ZN(net5572)
);

XOR2_X2 c5237(
.A(net5569),
.B(net4608),
.Z(net5573)
);

XNOR2_X1 c5238(
.A(net3645),
.B(net11440),
.ZN(net5574)
);

OR2_X4 c5239(
.A1(net2528),
.A2(net5564),
.ZN(net5575)
);

OR2_X1 c5240(
.A1(net5571),
.A2(net5353),
.ZN(net5576)
);

XNOR2_X2 c5241(
.A(net4662),
.B(net5574),
.ZN(net5577)
);

INV_X32 c5242(
.A(net5516),
.ZN(net5578)
);

AND2_X4 c5243(
.A1(net4659),
.A2(net4633),
.ZN(net5579)
);

AND2_X1 c5244(
.A1(net4591),
.A2(net4615),
.ZN(net5580)
);

NAND2_X1 c5245(
.A1(net4524),
.A2(net10638),
.ZN(net5581)
);

NAND2_X2 c5246(
.A1(net4465),
.A2(net2528),
.ZN(net5582)
);

INV_X4 c5247(
.A(net4637),
.ZN(net5583)
);

NAND2_X4 c5248(
.A1(net5472),
.A2(net5583),
.ZN(net5584)
);

AND2_X2 c5249(
.A1(net4597),
.A2(net4562),
.ZN(net5585)
);

XOR2_X1 c5250(
.A(net720),
.B(net10972),
.Z(net5586)
);

NOR2_X1 c5251(
.A1(net5568),
.A2(net5542),
.ZN(net5587)
);

INV_X1 c5252(
.A(net5577),
.ZN(net5588)
);

OR2_X2 c5253(
.A1(net5506),
.A2(net3676),
.ZN(net5589)
);

NOR2_X4 c5254(
.A1(net5588),
.A2(net4562),
.ZN(net5590)
);

NOR2_X2 c5255(
.A1(net4641),
.A2(net3622),
.ZN(net5591)
);

INV_X2 c5256(
.A(net4265),
.ZN(net5592)
);

XOR2_X2 c5257(
.A(net4615),
.B(net10613),
.Z(net5593)
);

XNOR2_X1 c5258(
.A(net5507),
.B(net3668),
.ZN(net5594)
);

INV_X8 c5259(
.A(net4530),
.ZN(net5595)
);

OR2_X4 c5260(
.A1(net4667),
.A2(net5228),
.ZN(net5596)
);

INV_X16 c5261(
.A(net9998),
.ZN(net5597)
);

INV_X32 c5262(
.A(net11390),
.ZN(net5598)
);

OR2_X1 c5263(
.A1(net5538),
.A2(net3627),
.ZN(net5599)
);

INV_X4 c5264(
.A(net11484),
.ZN(net5600)
);

XNOR2_X2 c5265(
.A(net5572),
.B(net4334),
.ZN(net5601)
);

AND2_X4 c5266(
.A1(net4603),
.A2(net10637),
.ZN(net5602)
);

AND2_X1 c5267(
.A1(net5524),
.A2(net4641),
.ZN(net5603)
);

NAND2_X1 c5268(
.A1(net5592),
.A2(net4392),
.ZN(net5604)
);

NAND2_X2 c5269(
.A1(net5585),
.A2(net5602),
.ZN(net5605)
);

INV_X1 c5270(
.A(net11411),
.ZN(net5606)
);

NAND2_X4 c5271(
.A1(net5573),
.A2(net5567),
.ZN(net5607)
);

INV_X2 c5272(
.A(net10233),
.ZN(net5608)
);

INV_X8 c5273(
.A(net10394),
.ZN(net5609)
);

AND2_X2 c5274(
.A1(net4623),
.A2(net4542),
.ZN(net5610)
);

XOR2_X1 c5275(
.A(net5594),
.B(net5583),
.Z(net5611)
);

INV_X16 c5276(
.A(net10094),
.ZN(net5612)
);

MUX2_X2 c5277(
.A(net4569),
.B(net711),
.S(net4658),
.Z(net5613)
);

NOR2_X1 c5278(
.A1(net5611),
.A2(net5093),
.ZN(net5614)
);

DFFS_X2 c5279(
.D(net4661),
.SN(net5596),
.CK(clk),
.Q(net5616),
.QN(net5615)
);

INV_X32 c5280(
.A(net5600),
.ZN(net5617)
);

INV_X4 c5281(
.A(net5607),
.ZN(net5618)
);

OR2_X2 c5282(
.A1(net5613),
.A2(net5616),
.ZN(net5619)
);

NOR2_X4 c5283(
.A1(net5593),
.A2(net4615),
.ZN(net5620)
);

NOR2_X2 c5284(
.A1(net5620),
.A2(net5563),
.ZN(net5621)
);

XOR2_X2 c5285(
.A(net5582),
.B(net5619),
.Z(net5622)
);

XNOR2_X1 c5286(
.A(net4603),
.B(net5609),
.ZN(net5623)
);

OR2_X4 c5287(
.A1(net2526),
.A2(net5419),
.ZN(net5624)
);

OR2_X1 c5288(
.A1(net4646),
.A2(net5616),
.ZN(net5625)
);

XNOR2_X2 c5289(
.A(net5618),
.B(net5563),
.ZN(net5626)
);

NAND3_X4 c5290(
.A1(net5603),
.A2(net5621),
.A3(net5616),
.ZN(net5627)
);

AND2_X4 c5291(
.A1(net5619),
.A2(net5627),
.ZN(net5628)
);

AND2_X1 c5292(
.A1(net4495),
.A2(net5506),
.ZN(net5629)
);

INV_X1 c5293(
.A(net11382),
.ZN(net5630)
);

NAND2_X1 c5294(
.A1(net5617),
.A2(net5455),
.ZN(net5631)
);

AOI222_X2 c5295(
.A1(net5567),
.A2(net5631),
.B1(net4614),
.B2(net5580),
.C1(net5559),
.C2(net11231),
.ZN(net5632)
);

NAND2_X2 c5296(
.A1(net5624),
.A2(net5623),
.ZN(net5633)
);

INV_X2 c5297(
.A(net10171),
.ZN(net5634)
);

OR3_X4 c5298(
.A1(net5632),
.A2(net5595),
.A3(net4091),
.ZN(net5635)
);

OAI222_X1 c5299(
.A1(net3611),
.A2(net5631),
.B1(net5632),
.B2(out25),
.C1(net5615),
.C2(net4608),
.ZN(net5636)
);

AND3_X2 c5300(
.A1(net5630),
.A2(net5240),
.A3(net5625),
.ZN(net5637)
);

INV_X8 c5301(
.A(net11403),
.ZN(net5638)
);

NOR3_X1 c5302(
.A1(net5579),
.A2(net5635),
.A3(net5638),
.ZN(net5639)
);

DFFRS_X1 c5303(
.D(net5622),
.RN(net5619),
.SN(net5638),
.CK(clk),
.Q(net5641),
.QN(net5640)
);

AOI221_X2 c5304(
.A(net5093),
.B1(net5631),
.B2(net5634),
.C1(net5615),
.C2(out25),
.ZN(net5642)
);

OAI222_X4 c5305(
.A1(net5597),
.A2(net5637),
.B1(net5638),
.B2(net4495),
.C1(net5413),
.C2(net11231),
.ZN(net5643)
);

NAND2_X4 c5306(
.A1(net5598),
.A2(net5638),
.ZN(net5644)
);

OAI222_X2 c5307(
.A1(net5644),
.A2(net4534),
.B1(net5580),
.B2(net4523),
.C1(net5615),
.C2(net10771),
.ZN(net5645)
);

OR3_X2 c5308(
.A1(net5427),
.A2(net5639),
.A3(net11345),
.ZN(net5646)
);

AOI221_X1 c5309(
.A(net5642),
.B1(net5632),
.B2(net4633),
.C1(net5638),
.C2(net4592),
.ZN(net5647)
);

OAI21_X2 c5310(
.A(net5645),
.B1(net5646),
.B2(net5612),
.ZN(net5648)
);

DFFRS_X2 c5311(
.D(net5648),
.RN(net5638),
.SN(net5516),
.CK(clk),
.Q(net5650),
.QN(net5649)
);

AND2_X2 c5312(
.A1(net4614),
.A2(net3723),
.ZN(net5651)
);

OAI221_X1 c5313(
.A(net4679),
.B1(net4614),
.B2(net4680),
.C1(net5464),
.C2(net3742),
.ZN(net5652)
);

INV_X16 c5314(
.A(net10491),
.ZN(net5653)
);

XOR2_X1 c5315(
.A(net4739),
.B(net3741),
.Z(net5654)
);

INV_X32 c5316(
.A(net11363),
.ZN(net5655)
);

OAI21_X1 c5317(
.A(net5655),
.B1(net4664),
.B2(net5333),
.ZN(net5656)
);

NOR2_X1 c5318(
.A1(net5575),
.A2(net3749),
.ZN(net5657)
);

OR2_X2 c5319(
.A1(net4562),
.A2(net5654),
.ZN(net5658)
);

INV_X4 c5320(
.A(net10047),
.ZN(net5659)
);

INV_X1 c5321(
.A(net11228),
.ZN(net5660)
);

NOR2_X4 c5322(
.A1(net3779),
.A2(net3765),
.ZN(net5661)
);

NOR2_X2 c5323(
.A1(net4699),
.A2(net5583),
.ZN(net5662)
);

INV_X2 c5324(
.A(net11298),
.ZN(net5663)
);

XOR2_X2 c5325(
.A(net5433),
.B(net5654),
.Z(net5664)
);

XNOR2_X1 c5326(
.A(net3765),
.B(net5604),
.ZN(net5665)
);

OR2_X4 c5327(
.A1(net5606),
.A2(net5625),
.ZN(net5666)
);

OR2_X1 c5328(
.A1(net3496),
.A2(net5639),
.ZN(net5667)
);

XNOR2_X2 c5329(
.A(net3729),
.B(net840),
.ZN(net5668)
);

AND2_X4 c5330(
.A1(net5513),
.A2(net5666),
.ZN(net5669)
);

AND2_X1 c5331(
.A1(net5542),
.A2(net5660),
.ZN(net5670)
);

NAND2_X1 c5332(
.A1(net5639),
.A2(net4664),
.ZN(net5671)
);

NAND2_X2 c5333(
.A1(net5670),
.A2(net5655),
.ZN(net5672)
);

NAND2_X4 c5334(
.A1(net5567),
.A2(net5639),
.ZN(net5673)
);

INV_X8 c5335(
.A(net11252),
.ZN(net5674)
);

INV_X16 c5336(
.A(net9834),
.ZN(net5675)
);

AOI21_X2 c5337(
.A(net5419),
.B1(net2517),
.B2(net5560),
.ZN(net5676)
);

AND2_X2 c5338(
.A1(net472),
.A2(net5667),
.ZN(net5677)
);

AOI21_X1 c5339(
.A(net3741),
.B1(net5650),
.B2(net4714),
.ZN(net5678)
);

XOR2_X1 c5340(
.A(net3747),
.B(net3155),
.Z(net5679)
);

NOR2_X1 c5341(
.A1(net4676),
.A2(net5608),
.ZN(net5680)
);

INV_X32 c5342(
.A(net11464),
.ZN(net5681)
);

OR2_X2 c5343(
.A1(net3758),
.A2(net4334),
.ZN(net5682)
);

NOR2_X4 c5344(
.A1(net5626),
.A2(net4740),
.ZN(net5683)
);

AOI21_X4 c5345(
.A(net3770),
.B1(net3496),
.B2(net10520),
.ZN(net5684)
);

NOR2_X2 c5346(
.A1(net4745),
.A2(net4715),
.ZN(net5685)
);

XOR2_X2 c5347(
.A(net5667),
.B(net5685),
.Z(net5686)
);

AND3_X1 c5348(
.A1(net4615),
.A2(net5580),
.A3(net5604),
.ZN(net5687)
);

XNOR2_X1 c5349(
.A(net4658),
.B(net5662),
.ZN(net5688)
);

OR2_X4 c5350(
.A1(net5680),
.A2(net4676),
.ZN(net5689)
);

NAND3_X1 c5351(
.A1(net5654),
.A2(net5681),
.A3(net5240),
.ZN(net5690)
);

SDFF_X1 c5352(
.D(net1743),
.SE(net5669),
.SI(net3692),
.CK(clk),
.Q(net5692),
.QN(net5691)
);

OR2_X1 c5353(
.A1(net4687),
.A2(net5590),
.ZN(net5693)
);

XNOR2_X2 c5354(
.A(net5653),
.B(net5667),
.ZN(net5694)
);

AND2_X4 c5355(
.A1(net5675),
.A2(net5692),
.ZN(net5695)
);

INV_X4 c5356(
.A(net9805),
.ZN(net5696)
);

AND2_X1 c5357(
.A1(net5673),
.A2(net5681),
.ZN(net5697)
);

NAND2_X1 c5358(
.A1(net5689),
.A2(net10615),
.ZN(net5698)
);

NAND2_X2 c5359(
.A1(net5659),
.A2(net10708),
.ZN(net5699)
);

NAND2_X4 c5360(
.A1(net5682),
.A2(net5668),
.ZN(net5700)
);

SDFF_X2 c5361(
.D(net5414),
.SE(net5691),
.SI(net3747),
.CK(clk),
.Q(net5702),
.QN(net5701)
);

AND2_X2 c5362(
.A1(net5672),
.A2(net5700),
.ZN(net5703)
);

NOR3_X4 c5363(
.A1(net783),
.A2(net5668),
.A3(net5542),
.ZN(net5704)
);

XOR2_X1 c5364(
.A(net4334),
.B(net5701),
.Z(net5705)
);

DFFR_X1 c5365(
.D(net5566),
.RN(net5698),
.CK(clk),
.Q(net5707),
.QN(net5706)
);

INV_X1 c5366(
.A(net10183),
.ZN(net5708)
);

NOR2_X1 c5367(
.A1(net5657),
.A2(net5655),
.ZN(net5709)
);

OR2_X2 c5368(
.A1(net5697),
.A2(net5709),
.ZN(net5710)
);

NOR2_X4 c5369(
.A1(net5560),
.A2(net5709),
.ZN(net5711)
);

NOR3_X2 c5370(
.A1(net4668),
.A2(net5709),
.A3(net5707),
.ZN(net5712)
);

NOR2_X2 c5371(
.A1(net3497),
.A2(net5655),
.ZN(net5713)
);

DFFR_X2 c5372(
.D(net2517),
.RN(net5683),
.CK(clk),
.Q(net5715),
.QN(net5714)
);

INV_X2 c5373(
.A(net10270),
.ZN(net5716)
);

AND3_X4 c5374(
.A1(net4649),
.A2(net5686),
.A3(net5654),
.ZN(net5717)
);

DFFRS_X1 c5375(
.D(net5674),
.RN(net5716),
.SN(net5710),
.CK(clk),
.Q(net5719),
.QN(net5718)
);

INV_X8 c5376(
.A(net10308),
.ZN(net5720)
);

XOR2_X2 c5377(
.A(net5651),
.B(net5661),
.Z(net5721)
);

XNOR2_X1 c5378(
.A(net5477),
.B(net5711),
.ZN(net5722)
);

OR2_X4 c5379(
.A1(net5711),
.A2(net5700),
.ZN(net5723)
);

NAND3_X2 c5380(
.A1(net5608),
.A2(net5696),
.A3(net5722),
.ZN(net5724)
);

OR2_X1 c5381(
.A1(net5724),
.A2(net5483),
.ZN(net5725)
);

XNOR2_X2 c5382(
.A(net5455),
.B(net5703),
.ZN(net5726)
);

AND2_X4 c5383(
.A1(net5718),
.A2(net10519),
.ZN(net5727)
);

OAI221_X4 c5384(
.A(net5686),
.B1(net5727),
.B2(net4679),
.C1(net5654),
.C2(net5712),
.ZN(net5728)
);

SDFFRS_X1 c5385(
.D(net5712),
.RN(net5663),
.SE(net5727),
.SI(net5711),
.SN(net5704),
.CK(clk),
.Q(net5730),
.QN(net5729)
);

AND2_X1 c5386(
.A1(net5665),
.A2(net5671),
.ZN(net5731)
);

NAND2_X1 c5387(
.A1(net5720),
.A2(net10752),
.ZN(net5732)
);

NAND2_X2 c5388(
.A1(net5713),
.A2(net5687),
.ZN(net5733)
);

NAND2_X4 c5389(
.A1(net2735),
.A2(net5722),
.ZN(net5734)
);

OR3_X1 c5390(
.A1(net5681),
.A2(net5710),
.A3(net5729),
.ZN(net5735)
);

MUX2_X1 c5391(
.A(net5731),
.B(net5667),
.S(net11045),
.Z(net5736)
);

OAI221_X2 c5392(
.A(net4751),
.B1(net5723),
.B2(net4704),
.C1(net5729),
.C2(net5706),
.ZN(net5737)
);

AND2_X2 c5393(
.A1(net5625),
.A2(net5732),
.ZN(net5738)
);

INV_X16 c5394(
.A(net11363),
.ZN(net5739)
);

OAI21_X4 c5395(
.A(net1881),
.B1(net3820),
.B2(net5714),
.ZN(net5740)
);

XOR2_X1 c5396(
.A(net3702),
.B(net5464),
.Z(net5741)
);

NOR2_X1 c5397(
.A1(net4539),
.A2(net11521),
.ZN(net5742)
);

OR2_X2 c5398(
.A1(net5737),
.A2(net3789),
.ZN(net5743)
);

NOR2_X4 c5399(
.A1(net5715),
.A2(net4665),
.ZN(net5744)
);

INV_X32 c5400(
.A(net9760),
.ZN(net5745)
);

OAI22_X4 c5401(
.A1(net4817),
.A2(net4779),
.B1(net2848),
.B2(net4764),
.ZN(net5746)
);

AOI222_X1 c5402(
.A1(net3818),
.A2(net4757),
.B1(net4747),
.B2(net5649),
.C1(net4819),
.C2(net11534),
.ZN(net5747)
);

DFFS_X1 c5403(
.D(net5578),
.SN(net4766),
.CK(clk),
.Q(net5749),
.QN(net5748)
);

MUX2_X2 c5404(
.A(net5465),
.B(net4850),
.S(net4837),
.Z(net5750)
);

NAND3_X4 c5405(
.A1(net1840),
.A2(net3873),
.A3(net3723),
.ZN(net5751)
);

OR3_X4 c5406(
.A1(net4788),
.A2(net4850),
.A3(net11536),
.ZN(net5752)
);

DFFRS_X2 c5407(
.D(net4833),
.RN(net4776),
.SN(net5734),
.CK(clk),
.Q(net5754),
.QN(net5753)
);

INV_X4 c5408(
.A(net10294),
.ZN(net5755)
);

NOR2_X2 c5409(
.A1(net4763),
.A2(net3875),
.ZN(net5756)
);

XOR2_X2 c5410(
.A(net4850),
.B(net4788),
.Z(net5757)
);

XNOR2_X1 c5411(
.A(net2725),
.B(net4592),
.ZN(net5758)
);

OR2_X4 c5412(
.A1(net4665),
.A2(net10738),
.ZN(net5759)
);

OR2_X1 c5413(
.A1(net5756),
.A2(net5578),
.ZN(out16)
);

AND3_X2 c5414(
.A1(net5734),
.A2(net3865),
.A3(net10881),
.ZN(net5760)
);

NOR3_X1 c5415(
.A1(net2822),
.A2(net5734),
.A3(net5754),
.ZN(net5761)
);

OR3_X2 c5416(
.A1(net4747),
.A2(net5752),
.A3(net2713),
.ZN(net5762)
);

XNOR2_X2 c5417(
.A(net5741),
.B(net2854),
.ZN(net5763)
);

AND2_X4 c5418(
.A1(net4840),
.A2(net5719),
.ZN(net5764)
);

AND2_X1 c5419(
.A1(net4800),
.A2(net4812),
.ZN(net5765)
);

NAND2_X1 c5420(
.A1(net3838),
.A2(net11537),
.ZN(net5766)
);

OAI21_X2 c5421(
.A(net3865),
.B1(net3818),
.B2(net4818),
.ZN(net5767)
);

SDFF_X1 c5422(
.D(net3844),
.SE(net5737),
.SI(net3878),
.CK(clk),
.Q(net5769),
.QN(net5768)
);

NAND2_X2 c5423(
.A1(net4680),
.A2(net711),
.ZN(net5770)
);

NAND2_X4 c5424(
.A1(net5757),
.A2(net5751),
.ZN(net5771)
);

AND2_X2 c5425(
.A1(net5752),
.A2(net5580),
.ZN(net5772)
);

OAI21_X1 c5426(
.A(net5668),
.B1(net4713),
.B2(net4756),
.ZN(net5773)
);

AOI21_X2 c5427(
.A(net3837),
.B1(net5753),
.B2(net10845),
.ZN(net5774)
);

AOI21_X1 c5428(
.A(net5695),
.B1(net2751),
.B2(net4321),
.ZN(net5775)
);

XOR2_X1 c5429(
.A(net5751),
.B(net11537),
.Z(net5776)
);

NOR2_X1 c5430(
.A1(net5773),
.A2(net3846),
.ZN(net5777)
);

AOI21_X4 c5431(
.A(net5765),
.B1(net2821),
.B2(net3833),
.ZN(net5778)
);

DFFS_X2 c5432(
.D(net3798),
.SN(net5668),
.CK(clk),
.Q(net5780),
.QN(net5779)
);

AND3_X1 c5433(
.A1(net4826),
.A2(net2849),
.A3(net3833),
.ZN(net5781)
);

INV_X1 c5434(
.A(net10115),
.ZN(net5782)
);

OR2_X2 c5435(
.A1(net3874),
.A2(net11509),
.ZN(net5783)
);

NAND3_X1 c5436(
.A1(net1802),
.A2(net5776),
.A3(net10632),
.ZN(net5784)
);

SDFF_X2 c5437(
.D(net4818),
.SE(net5773),
.SI(net3849),
.CK(clk),
.Q(net5786),
.QN(net5785)
);

NOR3_X4 c5438(
.A1(net4713),
.A2(net2713),
.A3(net4665),
.ZN(net5787)
);

NOR2_X4 c5439(
.A1(net2594),
.A2(net5784),
.ZN(net5788)
);

NOR3_X2 c5440(
.A1(net5755),
.A2(net4781),
.A3(net11535),
.ZN(net5789)
);

AND3_X4 c5441(
.A1(net4780),
.A2(net4818),
.A3(net4776),
.ZN(net5790)
);

DFFRS_X1 c5442(
.D(net5690),
.RN(net5780),
.SN(net5773),
.CK(clk),
.Q(net5792),
.QN(net5791)
);

NOR2_X2 c5443(
.A1(net5778),
.A2(net5779),
.ZN(net5793)
);

NAND3_X2 c5444(
.A1(net5769),
.A2(net4763),
.A3(net5773),
.ZN(net5794)
);

XOR2_X2 c5445(
.A(net5788),
.B(net5715),
.Z(net5795)
);

DFFRS_X2 c5446(
.D(net5746),
.RN(net5787),
.SN(net3843),
.CK(clk),
.Q(net5797),
.QN(net5796)
);

INV_X2 c5447(
.A(net9759),
.ZN(net5798)
);

OR3_X1 c5448(
.A1(net5798),
.A2(net2821),
.A3(net10942),
.ZN(net5799)
);

XNOR2_X1 c5449(
.A(net3789),
.B(net4781),
.ZN(net5800)
);

OR2_X4 c5450(
.A1(net5774),
.A2(net2854),
.ZN(net5801)
);

MUX2_X1 c5451(
.A(net5772),
.B(net5773),
.S(net5768),
.Z(net5802)
);

INV_X8 c5452(
.A(net10217),
.ZN(net5803)
);

OR2_X1 c5453(
.A1(net5799),
.A2(net5772),
.ZN(net5804)
);

SDFF_X1 c5454(
.D(net5766),
.SE(net5804),
.SI(net4839),
.CK(clk),
.Q(net5806),
.QN(net5805)
);

OAI21_X4 c5455(
.A(net5801),
.B1(net5764),
.B2(net11521),
.ZN(net5807)
);

SDFF_X2 c5456(
.D(net5775),
.SE(net5787),
.SI(net5795),
.CK(clk),
.Q(net5809),
.QN(net5808)
);

DFFRS_X1 c5457(
.D(net5787),
.RN(net3810),
.SN(net5695),
.CK(clk),
.Q(net5811),
.QN(net5810)
);

MUX2_X2 c5458(
.A(net5806),
.B(net5785),
.S(net5764),
.Z(net5812)
);

NAND3_X4 c5459(
.A1(net3723),
.A2(net4819),
.A3(net5805),
.ZN(net5813)
);

OR3_X4 c5460(
.A1(net4766),
.A2(net5771),
.A3(net5751),
.ZN(net5814)
);

XNOR2_X2 c5461(
.A(net5809),
.B(net5805),
.ZN(net5815)
);

AND3_X2 c5462(
.A1(net5813),
.A2(net5719),
.A3(net5795),
.ZN(net5816)
);

DFFRS_X2 c5463(
.D(net4807),
.RN(net5807),
.SN(net5784),
.CK(clk),
.Q(net5818),
.QN(net5817)
);

INV_X16 c5464(
.A(net10093),
.ZN(net5819)
);

AND2_X4 c5465(
.A1(net4808),
.A2(net5802),
.ZN(net5820)
);

SDFF_X1 c5466(
.D(net5800),
.SE(net5808),
.SI(net5788),
.CK(clk),
.Q(net5822),
.QN(net5821)
);

NOR3_X1 c5467(
.A1(net4847),
.A2(net5716),
.A3(net5816),
.ZN(net5823)
);

OR3_X2 c5468(
.A1(net5793),
.A2(net5813),
.A3(net5795),
.ZN(net5824)
);

OAI21_X2 c5469(
.A(net5751),
.B1(net5806),
.B2(net5757),
.ZN(net5825)
);

SDFF_X2 c5470(
.D(net5812),
.SE(net4766),
.SI(net10905),
.CK(clk),
.Q(net5827),
.QN(net5826)
);

AOI22_X2 c5471(
.A1(net5783),
.A2(net5786),
.B1(net5826),
.B2(net11520),
.ZN(net5828)
);

AND2_X1 c5472(
.A1(net4810),
.A2(net5799),
.ZN(net5829)
);

OAI21_X1 c5473(
.A(net5763),
.B1(net5791),
.B2(net11034),
.ZN(net5830)
);

AOI222_X4 c5474(
.A1(net5737),
.A2(net5791),
.B1(out25),
.B2(net5753),
.C1(net10973),
.C2(net11509),
.ZN(net5831)
);

OAI33_X1 c5475(
.A1(net5829),
.A2(net5830),
.A3(net5827),
.B1(net5668),
.B2(net3691),
.B3(out25),
.ZN(net5832)
);

AOI21_X2 c5476(
.A(net5825),
.B1(net5828),
.B2(net11546),
.ZN(net5833)
);

AOI21_X1 c5477(
.A(net5798),
.B1(net5833),
.B2(net11547),
.ZN(net5834)
);

NAND2_X1 c5478(
.A1(net4918),
.A2(net2945),
.ZN(net5835)
);

INV_X32 c5479(
.A(net4888),
.ZN(net5836)
);

INV_X4 c5480(
.A(net4910),
.ZN(net5837)
);

INV_X1 c5481(
.A(net4888),
.ZN(net5838)
);

INV_X2 c5482(
.A(net4903),
.ZN(net5839)
);

INV_X8 c5483(
.A(net2945),
.ZN(net5840)
);

INV_X16 c5484(
.A(net4872),
.ZN(net5841)
);

INV_X32 c5485(
.A(net5837),
.ZN(net5842)
);

INV_X4 c5486(
.A(net3897),
.ZN(net5843)
);

DFFR_X1 c5487(
.D(net4877),
.RN(net4935),
.CK(clk),
.Q(net5845),
.QN(net5844)
);

INV_X1 c5488(
.A(net4920),
.ZN(net5846)
);

INV_X2 c5489(
.A(net5842),
.ZN(net5847)
);

INV_X8 c5490(
.A(net4939),
.ZN(net5848)
);

INV_X16 c5491(
.A(net3930),
.ZN(net5849)
);

NAND2_X2 c5492(
.A1(net4871),
.A2(net5849),
.ZN(net5850)
);

NAND2_X4 c5493(
.A1(net4870),
.A2(net5849),
.ZN(net5851)
);

INV_X32 c5494(
.A(net4930),
.ZN(net5852)
);

AND2_X2 c5495(
.A1(net4909),
.A2(net2902),
.ZN(net5853)
);

INV_X4 c5496(
.A(net3969),
.ZN(net5854)
);

INV_X1 c5497(
.A(net988),
.ZN(net5855)
);

INV_X2 c5498(
.A(net9789),
.ZN(net5856)
);

INV_X8 c5499(
.A(net4930),
.ZN(net5857)
);

INV_X16 c5500(
.A(net9788),
.ZN(net5858)
);

INV_X32 c5501(
.A(net5846),
.ZN(net5859)
);

INV_X4 c5502(
.A(net9818),
.ZN(net5860)
);

XOR2_X1 c5503(
.A(net1016),
.B(net4872),
.Z(net5861)
);

DFFR_X2 c5504(
.D(net5838),
.RN(net4928),
.CK(clk),
.Q(net5863),
.QN(net5862)
);

INV_X1 c5505(
.A(net5852),
.ZN(net5864)
);

INV_X2 c5506(
.A(net4913),
.ZN(net5865)
);

DFFS_X1 c5507(
.D(net5842),
.SN(net3904),
.CK(clk),
.Q(net5867),
.QN(net5866)
);

AOI21_X4 c5508(
.A(net5846),
.B1(net4920),
.B2(net4869),
.ZN(net5868)
);

NOR2_X1 c5509(
.A1(net5858),
.A2(net5842),
.ZN(net5869)
);

INV_X8 c5510(
.A(net4946),
.ZN(net5870)
);

OR2_X2 c5511(
.A1(net5865),
.A2(net4929),
.ZN(net5871)
);

INV_X16 c5512(
.A(net10552),
.ZN(net5872)
);

INV_X32 c5513(
.A(net3954),
.ZN(net5873)
);

INV_X4 c5514(
.A(net5867),
.ZN(net5874)
);

AND3_X1 c5515(
.A1(net5873),
.A2(net5842),
.A3(net5859),
.ZN(net5875)
);

NOR2_X4 c5516(
.A1(net3897),
.A2(net4909),
.ZN(net5876)
);

INV_X1 c5517(
.A(net5871),
.ZN(net5877)
);

INV_X2 c5518(
.A(net5844),
.ZN(net5878)
);

INV_X8 c5519(
.A(net9985),
.ZN(net5879)
);

INV_X16 c5520(
.A(net5873),
.ZN(net5880)
);

INV_X32 c5521(
.A(net5850),
.ZN(net5881)
);

NOR2_X2 c5522(
.A1(net5877),
.A2(net5857),
.ZN(net5882)
);

INV_X4 c5523(
.A(net4882),
.ZN(net5883)
);

INV_X1 c5524(
.A(net5879),
.ZN(net5884)
);

INV_X2 c5525(
.A(net9862),
.ZN(net5885)
);

XOR2_X2 c5526(
.A(net5858),
.B(net5859),
.Z(net5886)
);

XNOR2_X1 c5527(
.A(net2006),
.B(net5868),
.ZN(net5887)
);

NAND3_X1 c5528(
.A1(net5874),
.A2(net5884),
.A3(net4862),
.ZN(net5888)
);

DFFS_X2 c5529(
.D(net4877),
.SN(net5836),
.CK(clk),
.Q(net5890),
.QN(net5889)
);

INV_X8 c5530(
.A(net9884),
.ZN(net5891)
);

INV_X16 c5531(
.A(net5868),
.ZN(net5892)
);

INV_X32 c5532(
.A(net4903),
.ZN(net5893)
);

INV_X4 c5533(
.A(net5863),
.ZN(net5894)
);

INV_X1 c5534(
.A(net5860),
.ZN(net5895)
);

INV_X2 c5535(
.A(net5890),
.ZN(net5896)
);

OR2_X4 c5536(
.A1(net5886),
.A2(net5896),
.ZN(net5897)
);

DFFR_X1 c5537(
.D(net5892),
.RN(net2945),
.CK(clk),
.Q(net5899),
.QN(net5898)
);

INV_X8 c5538(
.A(net5855),
.ZN(net5900)
);

INV_X16 c5539(
.A(net5888),
.ZN(net5901)
);

INV_X32 c5540(
.A(net9935),
.ZN(net5902)
);

DFFRS_X1 c5541(
.D(net5887),
.RN(net5902),
.SN(net5870),
.CK(clk),
.Q(net5904),
.QN(net5903)
);

NOR3_X4 c5542(
.A1(net5884),
.A2(net5873),
.A3(net5902),
.ZN(net5905)
);

NOR3_X2 c5543(
.A1(net5875),
.A2(net5866),
.A3(net5874),
.ZN(net5906)
);

AND3_X4 c5544(
.A1(net5893),
.A2(net5905),
.A3(net5894),
.ZN(net5907)
);

DFFRS_X2 c5545(
.D(net5902),
.RN(net5862),
.SN(net5843),
.CK(clk),
.Q(net5909),
.QN(net5908)
);

DFFR_X2 c5546(
.D(net5840),
.RN(net5907),
.CK(clk),
.Q(net5911),
.QN(net5910)
);

OR2_X1 c5547(
.A1(net5904),
.A2(net5910),
.ZN(net5912)
);

NAND3_X2 c5548(
.A1(net5863),
.A2(net5894),
.A3(net5902),
.ZN(net5913)
);

OR3_X1 c5549(
.A1(net5905),
.A2(net5872),
.A3(net10561),
.ZN(net5914)
);

SDFFR_X2 c5550(
.D(net5907),
.RN(net5890),
.SE(net5835),
.SI(net5894),
.CK(clk),
.Q(net5916),
.QN(net5915)
);

MUX2_X1 c5551(
.A(net4878),
.B(net4945),
.S(net5910),
.Z(net5917)
);

XNOR2_X2 c5552(
.A(net5893),
.B(net10562),
.ZN(net5918)
);

OAI21_X4 c5553(
.A(net5895),
.B1(net5917),
.B2(net3968),
.ZN(net5919)
);

AOI222_X2 c5554(
.A1(net5878),
.A2(net5908),
.B1(net5889),
.B2(net5859),
.C1(net5883),
.C2(net4935),
.ZN(net5920)
);

MUX2_X2 c5555(
.A(net5885),
.B(net5915),
.S(net5913),
.Z(net5921)
);

SDFF_X1 c5556(
.D(net5917),
.SE(net3930),
.SI(net5883),
.CK(clk),
.Q(net5923),
.QN(net5922)
);

AND2_X4 c5557(
.A1(net5921),
.A2(net5871),
.ZN(net5924)
);

NAND3_X4 c5558(
.A1(net5901),
.A2(net5924),
.A3(net1016),
.ZN(net5925)
);

SDFFS_X1 c5559(
.D(net5923),
.SE(net5918),
.SI(net5921),
.SN(net5925),
.CK(clk),
.Q(net5927),
.QN(net5926)
);

NAND4_X4 c5560(
.A1(net5896),
.A2(net5922),
.A3(net5850),
.A4(net5924),
.ZN(net5928)
);

INV_X4 c5561(
.A(net4962),
.ZN(net5929)
);

INV_X1 c5562(
.A(net11049),
.ZN(net5930)
);

AND2_X1 c5563(
.A1(net5851),
.A2(net4954),
.ZN(net5931)
);

NAND2_X1 c5564(
.A1(net2081),
.A2(net5024),
.ZN(net5932)
);

INV_X2 c5565(
.A(net4923),
.ZN(net5933)
);

DFFS_X1 c5566(
.D(net5015),
.SN(net5836),
.CK(clk),
.Q(net5935),
.QN(net5934)
);

NAND2_X2 c5567(
.A1(net5836),
.A2(net11103),
.ZN(net5936)
);

OR3_X4 c5568(
.A1(net5018),
.A2(net5861),
.A3(net4969),
.ZN(net5937)
);

NAND2_X4 c5569(
.A1(net5853),
.A2(net4974),
.ZN(net5938)
);

AND2_X2 c5570(
.A1(net4897),
.A2(net5934),
.ZN(net5939)
);

XOR2_X1 c5571(
.A(net3982),
.B(net4902),
.Z(net5940)
);

NOR2_X1 c5572(
.A1(net5927),
.A2(net2081),
.ZN(net5941)
);

INV_X8 c5573(
.A(net9690),
.ZN(net5942)
);

OR2_X2 c5574(
.A1(net4995),
.A2(net5872),
.ZN(net5943)
);

NOR2_X4 c5575(
.A1(net3955),
.A2(net4936),
.ZN(net5944)
);

INV_X16 c5576(
.A(net5022),
.ZN(net5945)
);

NOR2_X2 c5577(
.A1(net3991),
.A2(net5018),
.ZN(net5946)
);

XOR2_X2 c5578(
.A(net4908),
.B(net5903),
.Z(net5947)
);

INV_X32 c5579(
.A(net11011),
.ZN(net5948)
);

INV_X4 c5580(
.A(net9690),
.ZN(net5949)
);

XNOR2_X1 c5581(
.A(net4908),
.B(net10581),
.ZN(net5950)
);

OR2_X4 c5582(
.A1(net5918),
.A2(net5851),
.ZN(net5951)
);

INV_X1 c5583(
.A(net5881),
.ZN(net5952)
);

AND3_X2 c5584(
.A1(net5951),
.A2(net3991),
.A3(net4949),
.ZN(net5953)
);

INV_X2 c5585(
.A(net10383),
.ZN(net5954)
);

INV_X8 c5586(
.A(net4969),
.ZN(net5955)
);

INV_X16 c5587(
.A(net10502),
.ZN(net5956)
);

NOR3_X1 c5588(
.A1(net5841),
.A2(net5836),
.A3(net1922),
.ZN(net5957)
);

INV_X32 c5589(
.A(net5909),
.ZN(net5958)
);

INV_X4 c5590(
.A(net942),
.ZN(net5959)
);

INV_X1 c5591(
.A(net9883),
.ZN(net5960)
);

INV_X2 c5592(
.A(net3054),
.ZN(net5961)
);

INV_X8 c5593(
.A(net10158),
.ZN(net5962)
);

DFFS_X2 c5594(
.D(net5954),
.SN(net3038),
.CK(clk),
.Q(net5964),
.QN(net5963)
);

OR2_X1 c5595(
.A1(net4908),
.A2(net2902),
.ZN(net5965)
);

XNOR2_X2 c5596(
.A(net4983),
.B(net4962),
.ZN(net5966)
);

AND2_X4 c5597(
.A1(net5939),
.A2(net5962),
.ZN(net5967)
);

AND2_X1 c5598(
.A1(net5964),
.A2(net5939),
.ZN(net5968)
);

INV_X16 c5599(
.A(net5930),
.ZN(net5969)
);

INV_X32 c5600(
.A(net9863),
.ZN(net5970)
);

INV_X4 c5601(
.A(net10504),
.ZN(net5971)
);

NAND2_X1 c5602(
.A1(net5959),
.A2(net10889),
.ZN(net5972)
);

NAND2_X2 c5603(
.A1(net5960),
.A2(net4996),
.ZN(net5973)
);

NAND2_X4 c5604(
.A1(net5959),
.A2(net5945),
.ZN(net5974)
);

AND2_X2 c5605(
.A1(net5961),
.A2(net3054),
.ZN(net5975)
);

INV_X1 c5606(
.A(net5958),
.ZN(net5976)
);

INV_X2 c5607(
.A(net10056),
.ZN(net5977)
);

XOR2_X1 c5608(
.A(net4937),
.B(net5955),
.Z(net5978)
);

SDFF_X2 c5609(
.D(net5963),
.SE(net5975),
.SI(net5002),
.CK(clk),
.Q(net5980),
.QN(net5979)
);

NOR2_X1 c5610(
.A1(net5872),
.A2(net5021),
.ZN(net5981)
);

INV_X8 c5611(
.A(net5880),
.ZN(net5982)
);

INV_X16 c5612(
.A(net5968),
.ZN(net5983)
);

OR3_X2 c5613(
.A1(net5952),
.A2(net5967),
.A3(net5940),
.ZN(net5984)
);

DFFR_X1 c5614(
.D(net5944),
.RN(net5982),
.CK(clk),
.Q(net5986),
.QN(net5985)
);

OR2_X2 c5615(
.A1(net5981),
.A2(net5036),
.ZN(net5987)
);

INV_X32 c5616(
.A(net11049),
.ZN(net5988)
);

NOR2_X4 c5617(
.A1(net5987),
.A2(net5931),
.ZN(net5989)
);

OAI21_X2 c5618(
.A(net4040),
.B1(net5981),
.B2(net5980),
.ZN(net5990)
);

NOR2_X2 c5619(
.A1(net5989),
.A2(net5987),
.ZN(net5991)
);

OAI211_X2 c5620(
.A(net4974),
.B(net5952),
.C1(net5926),
.C2(net153),
.ZN(net5992)
);

OAI21_X1 c5621(
.A(net5969),
.B1(net5974),
.B2(net4953),
.ZN(net5993)
);

INV_X4 c5622(
.A(net10073),
.ZN(net5994)
);

XOR2_X2 c5623(
.A(net5971),
.B(net5962),
.Z(net5995)
);

XNOR2_X1 c5624(
.A(net5970),
.B(net5952),
.ZN(net5996)
);

AOI21_X2 c5625(
.A(net5931),
.B1(net5974),
.B2(net10731),
.ZN(net5997)
);

OR2_X4 c5626(
.A1(net5972),
.A2(net5974),
.ZN(net5998)
);

SDFFS_X2 c5627(
.D(net5991),
.SE(net5946),
.SI(net5980),
.SN(net5925),
.CK(clk),
.Q(net6000),
.QN(net5999)
);

OR2_X1 c5628(
.A1(net5993),
.A2(net4992),
.ZN(net6001)
);

INV_X1 c5629(
.A(net11010),
.ZN(net6002)
);

AOI21_X1 c5630(
.A(net5928),
.B1(net5987),
.B2(net11008),
.ZN(net6003)
);

XNOR2_X2 c5631(
.A(net5976),
.B(net4024),
.ZN(net6004)
);

AND2_X4 c5632(
.A1(net5982),
.A2(net4935),
.ZN(net6005)
);

OR4_X2 c5633(
.A1(net5997),
.A2(net5960),
.A3(net3054),
.A4(net5975),
.ZN(net6006)
);

AOI21_X4 c5634(
.A(net6002),
.B1(net6000),
.B2(net10924),
.ZN(net6007)
);

DFFRS_X1 c5635(
.D(net5836),
.RN(net5958),
.SN(net10888),
.CK(clk),
.Q(net6009),
.QN(net6008)
);

INV_X2 c5636(
.A(net10388),
.ZN(net6010)
);

DFFRS_X2 c5637(
.D(net6008),
.RN(net5938),
.SN(net11011),
.CK(clk),
.Q(net6012),
.QN(net6011)
);

AND3_X1 c5638(
.A1(net6004),
.A2(net5983),
.A3(net4975),
.ZN(net6013)
);

NAND3_X1 c5639(
.A1(net6009),
.A2(net4937),
.A3(net5881),
.ZN(net6014)
);

AND2_X1 c5640(
.A1(net6014),
.A2(net6002),
.ZN(net6015)
);

NOR3_X4 c5641(
.A1(net5995),
.A2(net6000),
.A3(net6014),
.ZN(net6016)
);

SDFFR_X1 c5642(
.D(net6007),
.RN(net5997),
.SE(net3904),
.SI(net6014),
.CK(clk),
.Q(net6018),
.QN(net6017)
);

OAI222_X1 c5643(
.A1(net6016),
.A2(net3038),
.B1(net5938),
.B2(net5975),
.C1(net6014),
.C2(net5856),
.ZN(net6019)
);

INV_X8 c5644(
.A(net4996),
.ZN(net6020)
);

INV_X16 c5645(
.A(net4050),
.ZN(net6021)
);

NAND2_X1 c5646(
.A1(net3902),
.A2(net3054),
.ZN(net6022)
);

NAND2_X2 c5647(
.A1(net4997),
.A2(net5941),
.ZN(net6023)
);

INV_X32 c5648(
.A(net9865),
.ZN(net6024)
);

INV_X4 c5649(
.A(net9758),
.ZN(net6025)
);

INV_X1 c5650(
.A(net11551),
.ZN(net6026)
);

INV_X2 c5651(
.A(net4881),
.ZN(net6027)
);

INV_X8 c5652(
.A(net4024),
.ZN(net6028)
);

NOR3_X2 c5653(
.A1(net5021),
.A2(net6026),
.A3(net5119),
.ZN(net6029)
);

AOI211_X1 c5654(
.A(net5119),
.B(net4996),
.C1(net6023),
.C2(net4140),
.ZN(net6030)
);

NAND2_X4 c5655(
.A1(net5977),
.A2(net6029),
.ZN(net6031)
);

AND2_X2 c5656(
.A1(net5986),
.A2(net4935),
.ZN(net6032)
);

INV_X16 c5657(
.A(net9757),
.ZN(net6033)
);

INV_X32 c5658(
.A(net6023),
.ZN(net6034)
);

XOR2_X1 c5659(
.A(net4142),
.B(net11551),
.Z(net6035)
);

INV_X4 c5660(
.A(net9837),
.ZN(net6036)
);

INV_X1 c5661(
.A(net5023),
.ZN(net6037)
);

NOR2_X1 c5662(
.A1(net6029),
.A2(net6033),
.ZN(net6038)
);

OR2_X2 c5663(
.A1(net5973),
.A2(net5903),
.ZN(net6039)
);

INV_X2 c5664(
.A(net6033),
.ZN(net6040)
);

INV_X8 c5665(
.A(net5941),
.ZN(net6041)
);

INV_X16 c5666(
.A(net10041),
.ZN(net6042)
);

NOR2_X4 c5667(
.A1(net3161),
.A2(net5107),
.ZN(net6043)
);

NAND4_X2 c5668(
.A1(net6041),
.A2(net6023),
.A3(net6029),
.A4(net6026),
.ZN(net6044)
);

OR4_X4 c5669(
.A1(net6023),
.A2(net5985),
.A3(net5942),
.A4(net6033),
.ZN(net6045)
);

NOR2_X2 c5670(
.A1(net6034),
.A2(net4988),
.ZN(net6046)
);

INV_X32 c5671(
.A(net10140),
.ZN(net6047)
);

XOR2_X2 c5672(
.A(net6037),
.B(net6026),
.Z(net6048)
);

XNOR2_X1 c5673(
.A(net4935),
.B(net3054),
.ZN(net6049)
);

INV_X4 c5674(
.A(net4956),
.ZN(net6050)
);

INV_X1 c5675(
.A(net11002),
.ZN(net6051)
);

OR2_X4 c5676(
.A1(net6031),
.A2(net6022),
.ZN(net6052)
);

OR2_X1 c5677(
.A1(net6048),
.A2(net3054),
.ZN(net6053)
);

AND3_X4 c5678(
.A1(net5071),
.A2(net4085),
.A3(net5962),
.ZN(net6054)
);

INV_X2 c5679(
.A(net6043),
.ZN(net6055)
);

INV_X8 c5680(
.A(net10902),
.ZN(net6056)
);

INV_X16 c5681(
.A(net11177),
.ZN(net6057)
);

INV_X32 c5682(
.A(net10045),
.ZN(net6058)
);

INV_X4 c5683(
.A(net6046),
.ZN(net6059)
);

XNOR2_X2 c5684(
.A(net6022),
.B(net6037),
.ZN(net6060)
);

INV_X1 c5685(
.A(net5845),
.ZN(net6061)
);

NAND3_X2 c5686(
.A1(net5119),
.A2(net5107),
.A3(net10747),
.ZN(net6062)
);

INV_X2 c5687(
.A(net9921),
.ZN(net6063)
);

INV_X8 c5688(
.A(net10204),
.ZN(net6064)
);

OR3_X1 c5689(
.A1(net6024),
.A2(net6063),
.A3(net4999),
.ZN(net6065)
);

INV_X16 c5690(
.A(net5966),
.ZN(net6066)
);

AND2_X4 c5691(
.A1(net6038),
.A2(net5946),
.ZN(net6067)
);

INV_X32 c5692(
.A(net10580),
.ZN(net6068)
);

AND2_X1 c5693(
.A1(net6055),
.A2(net6026),
.ZN(net6069)
);

INV_X4 c5694(
.A(net6061),
.ZN(net6070)
);

NAND2_X1 c5695(
.A1(net5983),
.A2(net6033),
.ZN(net6071)
);

MUX2_X1 c5696(
.A(net6057),
.B(net5057),
.S(net11550),
.Z(net6072)
);

OAI21_X4 c5697(
.A(net6063),
.B1(net6070),
.B2(net5052),
.ZN(net6073)
);

NAND2_X2 c5698(
.A1(net6051),
.A2(net5052),
.ZN(net6074)
);

NAND2_X4 c5699(
.A1(net6039),
.A2(net6020),
.ZN(net6075)
);

INV_X1 c5700(
.A(net6056),
.ZN(net6076)
);

AND2_X2 c5701(
.A1(net6064),
.A2(net6015),
.ZN(net6077)
);

INV_X2 c5702(
.A(net5121),
.ZN(net6078)
);

XOR2_X1 c5703(
.A(net6044),
.B(net6077),
.Z(net6079)
);

NOR2_X1 c5704(
.A1(net6074),
.A2(net6022),
.ZN(net6080)
);

OR2_X2 c5705(
.A1(net4988),
.A2(net6077),
.ZN(net6081)
);

MUX2_X2 c5706(
.A(net6070),
.B(net4140),
.S(net6077),
.Z(net6082)
);

INV_X8 c5707(
.A(net11132),
.ZN(net6083)
);

OAI22_X2 c5708(
.A1(net5089),
.A2(net5876),
.B1(net5941),
.B2(net5119),
.ZN(net6084)
);

NOR2_X4 c5709(
.A1(net6073),
.A2(net4973),
.ZN(net6085)
);

INV_X16 c5710(
.A(net10090),
.ZN(net6086)
);

INV_X32 c5711(
.A(net6086),
.ZN(net6087)
);

INV_X4 c5712(
.A(net10050),
.ZN(net6088)
);

NOR2_X2 c5713(
.A1(net6082),
.A2(net5100),
.ZN(net6089)
);

XOR2_X2 c5714(
.A(net5956),
.B(net6031),
.Z(net6090)
);

INV_X1 c5715(
.A(net11378),
.ZN(net6091)
);

NAND3_X4 c5716(
.A1(net5082),
.A2(net6090),
.A3(net6082),
.ZN(net6092)
);

XNOR2_X1 c5717(
.A(net6088),
.B(net6090),
.ZN(net6093)
);

SDFF_X1 c5718(
.D(net6079),
.SE(net6060),
.SI(net6091),
.CK(clk),
.Q(net6095),
.QN(net6094)
);

OR3_X4 c5719(
.A1(net6040),
.A2(net6042),
.A3(net6029),
.ZN(net6096)
);

SDFF_X2 c5720(
.D(net6085),
.SE(net6060),
.SI(net6021),
.CK(clk),
.Q(net6098),
.QN(net6097)
);

AND3_X2 c5721(
.A1(net6083),
.A2(net6029),
.A3(net5119),
.ZN(net6099)
);

OR2_X4 c5722(
.A1(net6091),
.A2(net11489),
.ZN(net6100)
);

OR2_X1 c5723(
.A1(net6099),
.A2(net10609),
.ZN(net6101)
);

XNOR2_X2 c5724(
.A(net6063),
.B(net10968),
.ZN(net6102)
);

NOR3_X1 c5725(
.A1(net6078),
.A2(net6079),
.A3(net6102),
.ZN(net6103)
);

DFFRS_X1 c5726(
.D(net6102),
.RN(net6103),
.SN(net6093),
.CK(clk),
.Q(net6105),
.QN(net6104)
);

OR3_X2 c5727(
.A1(net5895),
.A2(net4997),
.A3(net6072),
.ZN(net6106)
);

SDFFR_X2 c5728(
.D(net5127),
.RN(net5913),
.SE(net4207),
.SI(net3054),
.CK(clk),
.Q(net6108),
.QN(net6107)
);

INV_X2 c5729(
.A(net6047),
.ZN(net6109)
);

INV_X8 c5730(
.A(net11284),
.ZN(net6110)
);

INV_X16 c5731(
.A(net6077),
.ZN(net6111)
);

AND2_X4 c5732(
.A1(net6015),
.A2(net5177),
.ZN(net6112)
);

INV_X32 c5733(
.A(net5949),
.ZN(net6113)
);

INV_X4 c5734(
.A(net3258),
.ZN(net6114)
);

AND2_X1 c5735(
.A1(net1254),
.A2(net5174),
.ZN(net6115)
);

INV_X1 c5736(
.A(net2203),
.ZN(net6116)
);

INV_X2 c5737(
.A(net9754),
.ZN(net6117)
);

INV_X8 c5738(
.A(net9754),
.ZN(net6118)
);

NAND2_X1 c5739(
.A1(net5148),
.A2(net6100),
.ZN(net6119)
);

DFFR_X2 c5740(
.D(net2261),
.RN(net285),
.CK(clk),
.Q(net6121),
.QN(net6120)
);

INV_X16 c5741(
.A(net9922),
.ZN(net6122)
);

INV_X32 c5742(
.A(net5184),
.ZN(net6123)
);

NAND2_X2 c5743(
.A1(net5904),
.A2(net6072),
.ZN(net6124)
);

INV_X4 c5744(
.A(net6109),
.ZN(net6125)
);

NAND2_X4 c5745(
.A1(net6116),
.A2(net5110),
.ZN(net6126)
);

AND2_X2 c5746(
.A1(net5207),
.A2(net3248),
.ZN(net6127)
);

INV_X1 c5747(
.A(net5193),
.ZN(net6128)
);

AOI221_X4 c5748(
.A(net6127),
.B1(net5190),
.B2(net2142),
.C1(net4159),
.C2(net6125),
.ZN(net6129)
);

INV_X2 c5749(
.A(net5110),
.ZN(net6130)
);

INV_X8 c5750(
.A(net10194),
.ZN(net6131)
);

XOR2_X1 c5751(
.A(net4169),
.B(net6108),
.Z(net6132)
);

INV_X16 c5752(
.A(net6131),
.ZN(net6133)
);

INV_X32 c5753(
.A(net6112),
.ZN(net6134)
);

INV_X4 c5754(
.A(net2227),
.ZN(net6135)
);

NOR2_X1 c5755(
.A1(net6068),
.A2(net3223),
.ZN(net6136)
);

OR2_X2 c5756(
.A1(net6110),
.A2(net5037),
.ZN(net6137)
);

NOR2_X4 c5757(
.A1(net6126),
.A2(net5127),
.ZN(net6138)
);

NOR2_X2 c5758(
.A1(net4973),
.A2(net6126),
.ZN(net6139)
);

XOR2_X2 c5759(
.A(net6122),
.B(net5202),
.Z(net6140)
);

XNOR2_X1 c5760(
.A(net6125),
.B(net5148),
.ZN(net6141)
);

INV_X1 c5761(
.A(net10452),
.ZN(net6142)
);

OR2_X4 c5762(
.A1(net1220),
.A2(net6142),
.ZN(net6143)
);

INV_X2 c5763(
.A(net5037),
.ZN(net6144)
);

INV_X8 c5764(
.A(net9841),
.ZN(net6145)
);

DFFS_X1 c5765(
.D(net5162),
.SN(net4159),
.CK(clk),
.Q(net6147),
.QN(net6146)
);

OR2_X1 c5766(
.A1(net6133),
.A2(net6126),
.ZN(net6148)
);

INV_X16 c5767(
.A(net6145),
.ZN(net6149)
);

XNOR2_X2 c5768(
.A(net6119),
.B(net6148),
.ZN(net6150)
);

INV_X32 c5769(
.A(net6140),
.ZN(net6151)
);

INV_X4 c5770(
.A(net5144),
.ZN(net6152)
);

AND2_X4 c5771(
.A1(net6114),
.A2(net6146),
.ZN(net6153)
);

OAI21_X2 c5772(
.A(net6109),
.B1(net6069),
.B2(net6130),
.ZN(net6154)
);

OAI211_X4 c5773(
.A(net5204),
.B(net5945),
.C1(net6130),
.C2(net5999),
.ZN(net6155)
);

AND2_X1 c5774(
.A1(net5998),
.A2(net6071),
.ZN(net6156)
);

NAND2_X1 c5775(
.A1(net5861),
.A2(net6087),
.ZN(net6157)
);

INV_X1 c5776(
.A(net6157),
.ZN(net6158)
);

NAND2_X2 c5777(
.A1(net4228),
.A2(net5139),
.ZN(net6159)
);

INV_X2 c5778(
.A(net5126),
.ZN(net6160)
);

INV_X8 c5779(
.A(net6142),
.ZN(net6161)
);

NAND2_X4 c5780(
.A1(net4181),
.A2(net6123),
.ZN(net6162)
);

INV_X16 c5781(
.A(net6139),
.ZN(net6163)
);

AND2_X2 c5782(
.A1(net6123),
.A2(net6125),
.ZN(net6164)
);

INV_X32 c5783(
.A(net5187),
.ZN(net6165)
);

XOR2_X1 c5784(
.A(net6116),
.B(net5190),
.Z(net6166)
);

NOR2_X1 c5785(
.A1(net6154),
.A2(net3982),
.ZN(net6167)
);

INV_X4 c5786(
.A(net11402),
.ZN(net6168)
);

OAI211_X1 c5787(
.A(net6161),
.B(net6138),
.C1(net6107),
.C2(net6153),
.ZN(net6169)
);

OR2_X2 c5788(
.A1(net6144),
.A2(net3182),
.ZN(net6170)
);

INV_X1 c5789(
.A(net6151),
.ZN(net6171)
);

OAI21_X1 c5790(
.A(net6134),
.B1(net6166),
.B2(net6148),
.ZN(net6172)
);

NOR2_X4 c5791(
.A1(net6128),
.A2(net6138),
.ZN(net6173)
);

NOR2_X2 c5792(
.A1(net2198),
.A2(net6173),
.ZN(net6174)
);

XOR2_X2 c5793(
.A(net6162),
.B(net11474),
.Z(net6175)
);

XNOR2_X1 c5794(
.A(net6167),
.B(net6164),
.ZN(net6176)
);

INV_X2 c5795(
.A(net10277),
.ZN(net6177)
);

AOI21_X2 c5796(
.A(net6067),
.B1(net6147),
.B2(net6164),
.ZN(net6178)
);

AOI21_X1 c5797(
.A(net6173),
.B1(net6178),
.B2(net5207),
.ZN(net6179)
);

AOI21_X4 c5798(
.A(net4071),
.B1(net6163),
.B2(net6177),
.ZN(net6180)
);

OR2_X4 c5799(
.A1(net6169),
.A2(net6167),
.ZN(net6181)
);

OR2_X1 c5800(
.A1(net6111),
.A2(net6027),
.ZN(net6182)
);

NOR4_X4 c5801(
.A1(net6136),
.A2(net6172),
.A3(net6182),
.A4(net6175),
.ZN(net6183)
);

AOI221_X2 c5802(
.A(net6058),
.B1(net3182),
.B2(net5181),
.C1(net6105),
.C2(net6182),
.ZN(net6184)
);

AND3_X1 c5803(
.A1(net6137),
.A2(net6125),
.A3(net11185),
.ZN(net6185)
);

INV_X8 c5804(
.A(net10455),
.ZN(net6186)
);

NAND3_X1 c5805(
.A1(net6069),
.A2(net6186),
.A3(net11436),
.ZN(net6187)
);

XNOR2_X2 c5806(
.A(net6185),
.B(net6175),
.ZN(net6188)
);

AND2_X4 c5807(
.A1(net5101),
.A2(net11436),
.ZN(net6189)
);

AOI221_X1 c5808(
.A(net6159),
.B1(net6132),
.B2(net6182),
.C1(net3248),
.C2(net3182),
.ZN(net6190)
);

OAI221_X1 c5809(
.A(net6171),
.B1(net5110),
.B2(net6182),
.C1(net4194),
.C2(net10828),
.ZN(net6191)
);

AND2_X1 c5810(
.A1(net4276),
.A2(net5136),
.ZN(net6192)
);

NAND2_X1 c5811(
.A1(net6021),
.A2(net11467),
.ZN(net6193)
);

INV_X16 c5812(
.A(net4993),
.ZN(net6194)
);

NOR3_X4 c5813(
.A1(net5190),
.A2(net5279),
.A3(net6175),
.ZN(net6195)
);

NAND2_X2 c5814(
.A1(net5924),
.A2(net5273),
.ZN(net6196)
);

NAND2_X4 c5815(
.A1(net5929),
.A2(net5225),
.ZN(net6197)
);

INV_X32 c5816(
.A(net6045),
.ZN(net6198)
);

NOR3_X2 c5817(
.A1(net5009),
.A2(net6160),
.A3(net6071),
.ZN(net6199)
);

AND2_X2 c5818(
.A1(net6194),
.A2(net5243),
.ZN(net6200)
);

INV_X4 c5819(
.A(net11385),
.ZN(net6201)
);

INV_X1 c5820(
.A(net9644),
.ZN(net6202)
);

AND3_X4 c5821(
.A1(net5136),
.A2(net5139),
.A3(net5235),
.ZN(net6203)
);

INV_X2 c5822(
.A(net9643),
.ZN(net6204)
);

INV_X8 c5823(
.A(net11482),
.ZN(net6205)
);

XOR2_X1 c5824(
.A(net3248),
.B(net5962),
.Z(net6206)
);

INV_X16 c5825(
.A(net5273),
.ZN(net6207)
);

INV_X32 c5826(
.A(net6141),
.ZN(net6208)
);

NOR2_X1 c5827(
.A1(net6202),
.A2(net5228),
.ZN(net6209)
);

INV_X4 c5828(
.A(net6192),
.ZN(net6210)
);

INV_X1 c5829(
.A(net10230),
.ZN(net6211)
);

OR2_X2 c5830(
.A1(net5225),
.A2(net6045),
.ZN(net6212)
);

DFFS_X2 c5831(
.D(net6143),
.SN(net5277),
.CK(clk),
.Q(net6214),
.QN(net6213)
);

INV_X2 c5832(
.A(net6117),
.ZN(net6215)
);

INV_X8 c5833(
.A(net10391),
.ZN(net6216)
);

INV_X16 c5834(
.A(net11100),
.ZN(net6217)
);

INV_X32 c5835(
.A(net6147),
.ZN(net6218)
);

INV_X4 c5836(
.A(net5131),
.ZN(net6219)
);

INV_X1 c5837(
.A(net11043),
.ZN(net6220)
);

NOR2_X4 c5838(
.A1(net6025),
.A2(net6214),
.ZN(net6221)
);

NOR2_X2 c5839(
.A1(net6193),
.A2(net6215),
.ZN(net6222)
);

XOR2_X2 c5840(
.A(net5946),
.B(net6208),
.Z(net6223)
);

INV_X2 c5841(
.A(net10448),
.ZN(net6224)
);

XNOR2_X1 c5842(
.A(net5236),
.B(net2142),
.ZN(net6225)
);

OR2_X4 c5843(
.A1(net6189),
.A2(net6222),
.ZN(net6226)
);

OR2_X1 c5844(
.A1(net6200),
.A2(net6226),
.ZN(net6227)
);

XNOR2_X2 c5845(
.A(net4153),
.B(net6113),
.ZN(net6228)
);

AND2_X4 c5846(
.A1(net5216),
.A2(net5924),
.ZN(net6229)
);

AND2_X1 c5847(
.A1(net5269),
.A2(net6153),
.ZN(net6230)
);

NAND2_X1 c5848(
.A1(net4312),
.A2(net3248),
.ZN(net6231)
);

NAND2_X2 c5849(
.A1(net3296),
.A2(net6192),
.ZN(net6232)
);

NAND2_X4 c5850(
.A1(net6156),
.A2(net5181),
.ZN(net6233)
);

AND2_X2 c5851(
.A1(net4194),
.A2(net5131),
.ZN(net6234)
);

DFFRS_X2 c5852(
.D(net6199),
.RN(net6217),
.SN(net6231),
.CK(clk),
.Q(net6236),
.QN(net6235)
);

XOR2_X1 c5853(
.A(net6228),
.B(net6141),
.Z(net6237)
);

NAND3_X2 c5854(
.A1(net6203),
.A2(net6198),
.A3(net6228),
.ZN(net6238)
);

NOR2_X1 c5855(
.A1(net6207),
.A2(net6228),
.ZN(net6239)
);

OR3_X1 c5856(
.A1(net6204),
.A2(net6232),
.A3(net6234),
.ZN(net6240)
);

OR2_X2 c5857(
.A1(net6206),
.A2(net6234),
.ZN(net6241)
);

INV_X8 c5858(
.A(net10307),
.ZN(net6242)
);

NOR2_X4 c5859(
.A1(net6205),
.A2(net6235),
.ZN(net6243)
);

INV_X16 c5860(
.A(net6027),
.ZN(net6244)
);

INV_X32 c5861(
.A(net6215),
.ZN(net6245)
);

NOR2_X2 c5862(
.A1(net6225),
.A2(net6224),
.ZN(net6246)
);

XOR2_X2 c5863(
.A(net4206),
.B(net6175),
.Z(net6247)
);

MUX2_X1 c5864(
.A(net6247),
.B(net5296),
.S(net6223),
.Z(net6248)
);

XNOR2_X1 c5865(
.A(net6220),
.B(net6194),
.ZN(net6249)
);

SDFF_X1 c5866(
.D(net6246),
.SE(net6212),
.SI(net6240),
.CK(clk),
.Q(net6251),
.QN(net6250)
);

OR2_X4 c5867(
.A1(net6245),
.A2(net6239),
.ZN(net6252)
);

OR2_X1 c5868(
.A1(net6222),
.A2(net4194),
.ZN(net6253)
);

XNOR2_X2 c5869(
.A(net6226),
.B(net6214),
.ZN(net6254)
);

OAI21_X4 c5870(
.A(net6188),
.B1(net6252),
.B2(net6220),
.ZN(net6255)
);

MUX2_X2 c5871(
.A(net6198),
.B(net6236),
.S(net5287),
.Z(net6256)
);

NAND3_X4 c5872(
.A1(net6231),
.A2(net6250),
.A3(net6241),
.ZN(net6257)
);

AND2_X4 c5873(
.A1(net6210),
.A2(net6249),
.ZN(net6258)
);

OR3_X4 c5874(
.A1(net6242),
.A2(net6227),
.A3(net6216),
.ZN(net6259)
);

AND3_X2 c5875(
.A1(net6241),
.A2(net6245),
.A3(net4282),
.ZN(net6260)
);

NOR3_X1 c5876(
.A1(net6249),
.A2(net6219),
.A3(net6259),
.ZN(net6261)
);

OR3_X2 c5877(
.A1(net6244),
.A2(net6236),
.A3(net6205),
.ZN(net6262)
);

OAI21_X2 c5878(
.A(net6118),
.B1(net6262),
.B2(net6245),
.ZN(net6263)
);

INV_X4 c5879(
.A(net11486),
.ZN(net6264)
);

OAI21_X1 c5880(
.A(net4156),
.B1(net6235),
.B2(net5287),
.ZN(net6265)
);

AOI21_X2 c5881(
.A(net6258),
.B1(net6158),
.B2(net11208),
.ZN(net6266)
);

AOI21_X1 c5882(
.A(net6234),
.B1(net6266),
.B2(net11100),
.ZN(net6267)
);

AND2_X1 c5883(
.A1(net6254),
.A2(net6232),
.ZN(net6268)
);

OAI221_X4 c5884(
.A(net6158),
.B1(net6260),
.B2(net6265),
.C1(net6268),
.C2(net6093),
.ZN(net6269)
);

SDFF_X2 c5885(
.D(net4059),
.SE(net6252),
.SI(net6263),
.CK(clk),
.Q(net6271),
.QN(net6270)
);

AOI21_X4 c5886(
.A(net6243),
.B1(net6254),
.B2(net11283),
.ZN(net6272)
);

AND3_X1 c5887(
.A1(net5107),
.A2(net6266),
.A3(net6268),
.ZN(net6273)
);

NAND3_X1 c5888(
.A1(net6267),
.A2(net6240),
.A3(net6264),
.ZN(net6274)
);

NOR3_X4 c5889(
.A1(net4173),
.A2(net6274),
.A3(net6265),
.ZN(net6275)
);

NOR3_X2 c5890(
.A1(net6272),
.A2(net6273),
.A3(net6265),
.ZN(net6276)
);

SDFFRS_X2 c5891(
.D(net5208),
.RN(net6264),
.SE(net5225),
.SI(net6276),
.SN(net6259),
.CK(clk),
.Q(net6278),
.QN(net6277)
);

AND3_X4 c5892(
.A1(net6278),
.A2(net6276),
.A3(net11171),
.ZN(net6279)
);

INV_X1 c5893(
.A(net11283),
.ZN(net6280)
);

NAND2_X1 c5894(
.A1(net6160),
.A2(net1412),
.ZN(net6281)
);

INV_X2 c5895(
.A(net1400),
.ZN(net6282)
);

INV_X8 c5896(
.A(net9853),
.ZN(net6283)
);

INV_X16 c5897(
.A(net9796),
.ZN(net6284)
);

INV_X32 c5898(
.A(net5287),
.ZN(net6285)
);

INV_X4 c5899(
.A(net6219),
.ZN(net6286)
);

NAND2_X2 c5900(
.A1(net5312),
.A2(net6260),
.ZN(net6287)
);

NAND3_X2 c5901(
.A1(net6283),
.A2(net6224),
.A3(net6229),
.ZN(net6288)
);

DFFRS_X1 c5902(
.D(net6285),
.RN(net6172),
.SN(net6281),
.CK(clk),
.Q(net6290),
.QN(net6289)
);

INV_X1 c5903(
.A(net6268),
.ZN(net6291)
);

NAND2_X4 c5904(
.A1(net5371),
.A2(net6093),
.ZN(net6292)
);

AND2_X2 c5905(
.A1(net6268),
.A2(net10802),
.ZN(net6293)
);

INV_X2 c5906(
.A(net5296),
.ZN(net6294)
);

OR3_X1 c5907(
.A1(net5362),
.A2(net4322),
.A3(net4374),
.ZN(net6295)
);

INV_X8 c5908(
.A(net9795),
.ZN(net6296)
);

DFFR_X1 c5909(
.D(net6209),
.RN(net6296),
.CK(clk),
.Q(net6298),
.QN(net6297)
);

INV_X16 c5910(
.A(net11399),
.ZN(net6299)
);

INV_X32 c5911(
.A(net9825),
.ZN(net6300)
);

XOR2_X1 c5912(
.A(net6296),
.B(net1254),
.Z(net6301)
);

INV_X4 c5913(
.A(net10209),
.ZN(net6302)
);

INV_X1 c5914(
.A(net5307),
.ZN(net6303)
);

INV_X2 c5915(
.A(net5894),
.ZN(net6304)
);

DFFR_X2 c5916(
.D(net5379),
.RN(net6292),
.CK(clk),
.Q(net6306),
.QN(net6305)
);

INV_X8 c5917(
.A(net6230),
.ZN(net6307)
);

NOR2_X1 c5918(
.A1(net5310),
.A2(net11399),
.ZN(net6308)
);

OR2_X2 c5919(
.A1(net5194),
.A2(net6280),
.ZN(net6309)
);

NOR2_X4 c5920(
.A1(net6299),
.A2(net6219),
.ZN(net6310)
);

INV_X16 c5921(
.A(net9873),
.ZN(net6311)
);

NOR2_X2 c5922(
.A1(net6284),
.A2(net5304),
.ZN(net6312)
);

MUX2_X1 c5923(
.A(net6300),
.B(net5307),
.S(net6093),
.Z(net6313)
);

OAI21_X4 c5924(
.A(net6310),
.B1(net6283),
.B2(net6305),
.ZN(net6314)
);

DFFS_X1 c5925(
.D(net5277),
.SN(net6298),
.CK(clk),
.Q(net6316),
.QN(net6315)
);

XOR2_X2 c5926(
.A(net5284),
.B(net6162),
.Z(net6317)
);

XNOR2_X1 c5927(
.A(net6297),
.B(net10606),
.ZN(net6318)
);

OR2_X4 c5928(
.A1(net6286),
.A2(net6295),
.ZN(net6319)
);

INV_X32 c5929(
.A(net4346),
.ZN(net6320)
);

OR2_X1 c5930(
.A1(net4374),
.A2(net6318),
.ZN(net6321)
);

DFFS_X2 c5931(
.D(net6287),
.SN(net6280),
.CK(clk),
.Q(net6323),
.QN(net6322)
);

XNOR2_X2 c5932(
.A(net5370),
.B(net4205),
.ZN(net6324)
);

AND2_X4 c5933(
.A1(net6295),
.A2(net4401),
.ZN(net6325)
);

NOR4_X2 c5934(
.A1(net6304),
.A2(net6306),
.A3(net5364),
.A4(net6260),
.ZN(net6326)
);

AOI211_X4 c5935(
.A(net6303),
.B(net6310),
.C1(net6268),
.C2(net6293),
.ZN(net6327)
);

AND2_X1 c5936(
.A1(net3258),
.A2(net6284),
.ZN(net6328)
);

INV_X4 c5937(
.A(net10148),
.ZN(net6329)
);

NAND2_X1 c5938(
.A1(net6289),
.A2(net10605),
.ZN(net6330)
);

NAND2_X2 c5939(
.A1(net4353),
.A2(net6280),
.ZN(net6331)
);

INV_X1 c5940(
.A(net6330),
.ZN(net6332)
);

MUX2_X2 c5941(
.A(net6283),
.B(net5310),
.S(net11217),
.Z(net6333)
);

NAND2_X4 c5942(
.A1(net6309),
.A2(net5258),
.ZN(net6334)
);

INV_X2 c5943(
.A(net11479),
.ZN(net6335)
);

AND2_X2 c5944(
.A1(net6317),
.A2(net5234),
.ZN(net6336)
);

XOR2_X1 c5945(
.A(net6307),
.B(net6318),
.Z(net6337)
);

INV_X8 c5946(
.A(net10422),
.ZN(net6338)
);

NOR2_X1 c5947(
.A1(net6311),
.A2(net6337),
.ZN(net6339)
);

OR2_X2 c5948(
.A1(net6321),
.A2(net6303),
.ZN(net6340)
);

NOR2_X4 c5949(
.A1(net6294),
.A2(net6340),
.ZN(net6341)
);

NOR2_X2 c5950(
.A1(net5318),
.A2(net6162),
.ZN(net6342)
);

DFFR_X1 c5951(
.D(net4366),
.RN(net6276),
.CK(clk),
.Q(net6344),
.QN(net6343)
);

XOR2_X2 c5952(
.A(net6342),
.B(net6310),
.Z(net6345)
);

XNOR2_X1 c5953(
.A(net5378),
.B(net6323),
.ZN(net6346)
);

OR2_X4 c5954(
.A1(net6332),
.A2(net6343),
.ZN(net6347)
);

OAI221_X2 c5955(
.A(net6337),
.B1(net6113),
.B2(net5371),
.C1(net6345),
.C2(net5352),
.ZN(net6348)
);

NOR4_X1 c5956(
.A1(net6224),
.A2(net6344),
.A3(net6345),
.A4(net6348),
.ZN(net6349)
);

INV_X16 c5957(
.A(net6345),
.ZN(net6350)
);

NAND3_X4 c5958(
.A1(net6291),
.A2(net6343),
.A3(net6302),
.ZN(net6351)
);

OR2_X1 c5959(
.A1(net6344),
.A2(net6286),
.ZN(net6352)
);

XNOR2_X2 c5960(
.A(net4340),
.B(net6339),
.ZN(net6353)
);

AND2_X4 c5961(
.A1(net6352),
.A2(net6320),
.ZN(net6354)
);

OAI222_X4 c5962(
.A1(net4350),
.A2(net6316),
.B1(net6348),
.B2(net5307),
.C1(net5383),
.C2(net6333),
.ZN(net6355)
);

AOI211_X2 c5963(
.A(net5948),
.B(net4405),
.C1(net6309),
.C2(net6162),
.ZN(net6356)
);

AND2_X1 c5964(
.A1(net5230),
.A2(net6305),
.ZN(net6357)
);

OR3_X4 c5965(
.A1(net6327),
.A2(net6309),
.A3(net6345),
.ZN(net6358)
);

AND3_X2 c5966(
.A1(net6338),
.A2(net6356),
.A3(net6354),
.ZN(net6359)
);

AOI22_X1 c5967(
.A1(net6350),
.A2(net6303),
.B1(net6348),
.B2(net5351),
.ZN(net6360)
);

NOR3_X1 c5968(
.A1(net6349),
.A2(net6358),
.A3(net5362),
.ZN(net6361)
);

NAND2_X1 c5969(
.A1(net6325),
.A2(net11440),
.ZN(net6362)
);

NAND2_X2 c5970(
.A1(net6353),
.A2(net6339),
.ZN(net6363)
);

OR3_X2 c5971(
.A1(net6351),
.A2(net6362),
.A3(net10982),
.ZN(net6364)
);

NAND2_X4 c5972(
.A1(net6280),
.A2(net6363),
.ZN(net6365)
);

OAI21_X2 c5973(
.A(net6359),
.B1(net6340),
.B2(net6358),
.ZN(net6366)
);

OAI21_X1 c5974(
.A(net6362),
.B1(net6347),
.B2(net6356),
.ZN(net6367)
);

AOI221_X4 c5975(
.A(net6348),
.B1(net3432),
.B2(net6367),
.C1(net6263),
.C2(net11348),
.ZN(net6368)
);

AND2_X2 c5976(
.A1(net5166),
.A2(net6351),
.ZN(net6369)
);

INV_X32 c5977(
.A(net9974),
.ZN(net6370)
);

INV_X4 c5978(
.A(net6314),
.ZN(net6371)
);

INV_X1 c5979(
.A(net9696),
.ZN(net6372)
);

XOR2_X1 c5980(
.A(net5402),
.B(net6298),
.Z(net6373)
);

NOR2_X1 c5981(
.A1(net6335),
.A2(net6322),
.ZN(net6374)
);

OR2_X2 c5982(
.A1(net6339),
.A2(net6281),
.ZN(net6375)
);

INV_X2 c5983(
.A(net6281),
.ZN(net6376)
);

NOR2_X4 c5984(
.A1(net5351),
.A2(net10923),
.ZN(net6377)
);

INV_X8 c5985(
.A(net10169),
.ZN(net6378)
);

INV_X16 c5986(
.A(net6375),
.ZN(net6379)
);

INV_X32 c5987(
.A(net5412),
.ZN(net6380)
);

NOR2_X2 c5988(
.A1(net6282),
.A2(net5389),
.ZN(net6381)
);

INV_X4 c5989(
.A(net5470),
.ZN(net6382)
);

INV_X1 c5990(
.A(net6373),
.ZN(net6383)
);

XOR2_X2 c5991(
.A(net6316),
.B(net6351),
.Z(net6384)
);

AOI21_X2 c5992(
.A(net6348),
.B1(net6382),
.B2(net5423),
.ZN(net6385)
);

XNOR2_X1 c5993(
.A(net5446),
.B(net6374),
.ZN(net6386)
);

INV_X2 c5994(
.A(net6372),
.ZN(net6387)
);

OR2_X4 c5995(
.A1(net5962),
.A2(net5334),
.ZN(net6388)
);

OR2_X1 c5996(
.A1(net5391),
.A2(net6153),
.ZN(net6389)
);

XNOR2_X2 c5997(
.A(net5405),
.B(net6260),
.ZN(net6390)
);

INV_X8 c5998(
.A(net6260),
.ZN(net6391)
);

AOI21_X1 c5999(
.A(net6351),
.B1(net6333),
.B2(net5234),
.ZN(net6392)
);

INV_X16 c6000(
.A(net5476),
.ZN(net6393)
);

DFFRS_X2 c6001(
.D(net5965),
.RN(net6393),
.SN(net5408),
.CK(clk),
.Q(net6395),
.QN(net6394)
);

AND2_X4 c6002(
.A1(net6381),
.A2(net5321),
.ZN(net6396)
);

INV_X32 c6003(
.A(net10325),
.ZN(net6397)
);

AND2_X1 c6004(
.A1(net4423),
.A2(net6383),
.ZN(net6398)
);

NAND2_X1 c6005(
.A1(net2509),
.A2(net4451),
.ZN(net6399)
);

INV_X4 c6006(
.A(net9696),
.ZN(net6400)
);

NAND2_X2 c6007(
.A1(net6323),
.A2(net5414),
.ZN(net6401)
);

NAND2_X4 c6008(
.A1(net6374),
.A2(net6383),
.ZN(net6402)
);

AND2_X2 c6009(
.A1(net6367),
.A2(net4413),
.ZN(net6403)
);

INV_X1 c6010(
.A(net10790),
.ZN(net6404)
);

INV_X2 c6011(
.A(net10404),
.ZN(net6405)
);

XOR2_X1 c6012(
.A(net6153),
.B(net6403),
.Z(net6406)
);

INV_X8 c6013(
.A(net6401),
.ZN(net6407)
);

NOR2_X1 c6014(
.A1(net6400),
.A2(net4423),
.ZN(net6408)
);

OR2_X2 c6015(
.A1(net6370),
.A2(net5962),
.ZN(net6409)
);

NOR2_X4 c6016(
.A1(net6402),
.A2(net6278),
.ZN(net6410)
);

AND4_X4 c6017(
.A1(net6376),
.A2(net5224),
.A3(net5231),
.A4(net6302),
.ZN(net6411)
);

NOR2_X2 c6018(
.A1(net4479),
.A2(net6367),
.ZN(net6412)
);

XOR2_X2 c6019(
.A(net6341),
.B(net6348),
.Z(net6413)
);

XNOR2_X1 c6020(
.A(net6408),
.B(net5321),
.ZN(net6414)
);

OR2_X4 c6021(
.A1(net6030),
.A2(net6410),
.ZN(net6415)
);

AOI21_X4 c6022(
.A(net5334),
.B1(net5399),
.B2(net5476),
.ZN(net6416)
);

INV_X16 c6023(
.A(net10076),
.ZN(net6417)
);

AND3_X1 c6024(
.A1(net5445),
.A2(net6406),
.A3(net6218),
.ZN(net6418)
);

OR2_X1 c6025(
.A1(net6400),
.A2(net11022),
.ZN(net6419)
);

XNOR2_X2 c6026(
.A(net5334),
.B(net10789),
.ZN(net6420)
);

AND2_X4 c6027(
.A1(net6407),
.A2(net10583),
.ZN(net6421)
);

AND2_X1 c6028(
.A1(net5425),
.A2(net6367),
.ZN(net6422)
);

NAND2_X1 c6029(
.A1(net5453),
.A2(net6397),
.ZN(net6423)
);

NAND3_X1 c6030(
.A1(net6406),
.A2(net6417),
.A3(net6394),
.ZN(net6424)
);

INV_X32 c6031(
.A(net11458),
.ZN(net6425)
);

NAND2_X2 c6032(
.A1(net6422),
.A2(net6238),
.ZN(net6426)
);

INV_X4 c6033(
.A(net10251),
.ZN(net6427)
);

NAND2_X4 c6034(
.A1(net6421),
.A2(net4488),
.ZN(net6428)
);

AND2_X2 c6035(
.A1(net5899),
.A2(net5389),
.ZN(net6429)
);

SDFFS_X1 c6036(
.D(net6218),
.SE(net6425),
.SI(net6030),
.SN(net5234),
.CK(clk),
.Q(net6431),
.QN(net6430)
);

NOR3_X4 c6037(
.A1(net4451),
.A2(net6420),
.A3(net6425),
.ZN(net6432)
);

XOR2_X1 c6038(
.A(net6368),
.B(net5470),
.Z(net6433)
);

NOR2_X1 c6039(
.A1(net6398),
.A2(net6425),
.ZN(net6434)
);

OR2_X2 c6040(
.A1(net6385),
.A2(net6376),
.ZN(net6435)
);

NOR2_X4 c6041(
.A1(net6427),
.A2(net6432),
.ZN(net6436)
);

NOR2_X2 c6042(
.A1(net5422),
.A2(net6313),
.ZN(net6437)
);

INV_X1 c6043(
.A(net11184),
.ZN(net6438)
);

NOR3_X2 c6044(
.A1(net6417),
.A2(net6432),
.A3(net6423),
.ZN(net6439)
);

XOR2_X2 c6045(
.A(net6419),
.B(net6436),
.Z(net6440)
);

AND3_X4 c6046(
.A1(net6395),
.A2(net5412),
.A3(net6437),
.ZN(net6441)
);

INV_X2 c6047(
.A(net10374),
.ZN(net6442)
);

AOI221_X2 c6048(
.A(net6429),
.B1(net6436),
.B2(net6440),
.C1(net6397),
.C2(net6437),
.ZN(net6443)
);

XNOR2_X1 c6049(
.A(net6428),
.B(net6430),
.ZN(net6444)
);

OR2_X4 c6050(
.A1(net6416),
.A2(net6432),
.ZN(net6445)
);

AOI221_X1 c6051(
.A(net6412),
.B1(net5446),
.B2(net6429),
.C1(net6425),
.C2(net6440),
.ZN(net6446)
);

SDFF_X1 c6052(
.D(net6446),
.SE(net6412),
.SI(net6440),
.CK(clk),
.Q(net6448),
.QN(net6447)
);

OR2_X1 c6053(
.A1(net6436),
.A2(net6416),
.ZN(net6449)
);

SDFFRS_X1 c6054(
.D(net6403),
.RN(net6438),
.SE(net6434),
.SI(net6447),
.SN(net6333),
.CK(clk),
.Q(net6451),
.QN(net6450)
);

XNOR2_X2 c6055(
.A(net6433),
.B(net6447),
.ZN(net6452)
);

AND2_X4 c6056(
.A1(net6444),
.A2(net6398),
.ZN(net6453)
);

INV_X8 c6057(
.A(net9925),
.ZN(net6454)
);

OAI221_X1 c6058(
.A(net6424),
.B1(net6454),
.B2(net6378),
.C1(net6442),
.C2(net5413),
.ZN(net6455)
);

INV_X16 c6059(
.A(net10164),
.ZN(net6456)
);

INV_X32 c6060(
.A(net6445),
.ZN(net6457)
);

INV_X4 c6061(
.A(net6380),
.ZN(net6458)
);

AND2_X1 c6062(
.A1(net5454),
.A2(net5375),
.ZN(net6459)
);

NAND3_X2 c6063(
.A1(net4458),
.A2(net5545),
.A3(net10545),
.ZN(net6460)
);

INV_X1 c6064(
.A(net9750),
.ZN(net6461)
);

NAND2_X1 c6065(
.A1(net5321),
.A2(net5537),
.ZN(net6462)
);

INV_X2 c6066(
.A(net3448),
.ZN(net6463)
);

INV_X8 c6067(
.A(net10313),
.ZN(net6464)
);

NAND2_X2 c6068(
.A1(net6265),
.A2(net6438),
.ZN(net6465)
);

OR3_X1 c6069(
.A1(net6457),
.A2(net6465),
.A3(net6464),
.ZN(net6466)
);

NAND2_X4 c6070(
.A1(net4540),
.A2(net5228),
.ZN(net6467)
);

INV_X16 c6071(
.A(net3598),
.ZN(net6468)
);

AND2_X2 c6072(
.A1(net5508),
.A2(net5496),
.ZN(net6469)
);

INV_X32 c6073(
.A(net6456),
.ZN(net6470)
);

MUX2_X1 c6074(
.A(net5527),
.B(net4562),
.S(net6463),
.Z(net6471)
);

INV_X4 c6075(
.A(net5232),
.ZN(net6472)
);

INV_X1 c6076(
.A(net10346),
.ZN(net6473)
);

INV_X2 c6077(
.A(net10152),
.ZN(net6474)
);

XOR2_X1 c6078(
.A(net6438),
.B(net6462),
.Z(net6475)
);

INV_X8 c6079(
.A(net6379),
.ZN(net6476)
);

NOR2_X1 c6080(
.A1(net6389),
.A2(net6397),
.ZN(net6477)
);

OR2_X2 c6081(
.A1(net6477),
.A2(net5449),
.ZN(net6478)
);

NOR2_X4 c6082(
.A1(net6449),
.A2(net6418),
.ZN(net6479)
);

INV_X16 c6083(
.A(net10216),
.ZN(net6480)
);

INV_X32 c6084(
.A(net6473),
.ZN(net6481)
);

INV_X4 c6085(
.A(net10412),
.ZN(net6482)
);

INV_X1 c6086(
.A(net9749),
.ZN(net6483)
);

OAI21_X4 c6087(
.A(net4458),
.B1(net6471),
.B2(net4392),
.ZN(net6484)
);

NOR2_X2 c6088(
.A1(net5537),
.A2(net4442),
.ZN(net6485)
);

XOR2_X2 c6089(
.A(net6474),
.B(net6469),
.Z(net6486)
);

XNOR2_X1 c6090(
.A(net5424),
.B(net6485),
.ZN(net6487)
);

OR2_X4 c6091(
.A1(net5498),
.A2(net6485),
.ZN(net6488)
);

MUX2_X2 c6092(
.A(net5536),
.B(net6459),
.S(net5503),
.Z(net6489)
);

INV_X2 c6093(
.A(net10378),
.ZN(net6490)
);

OR2_X1 c6094(
.A1(net6475),
.A2(net6486),
.ZN(net6491)
);

XNOR2_X2 c6095(
.A(net6458),
.B(net6227),
.ZN(net6492)
);

AND2_X4 c6096(
.A1(net6485),
.A2(net6423),
.ZN(net6493)
);

SDFF_X2 c6097(
.D(net6420),
.SE(net6490),
.SI(net6484),
.CK(clk),
.Q(net6495),
.QN(net6494)
);

AND2_X1 c6098(
.A1(net1599),
.A2(net11353),
.ZN(net6496)
);

INV_X8 c6099(
.A(net11354),
.ZN(net6497)
);

NAND2_X1 c6100(
.A1(net6483),
.A2(net5375),
.ZN(net6498)
);

INV_X16 c6101(
.A(net10150),
.ZN(net6499)
);

NAND2_X2 c6102(
.A1(net6496),
.A2(net5228),
.ZN(net6500)
);

NAND2_X4 c6103(
.A1(net5503),
.A2(net6496),
.ZN(net6501)
);

AND2_X2 c6104(
.A1(net6404),
.A2(net5427),
.ZN(net6502)
);

NAND3_X4 c6105(
.A1(net6336),
.A2(net6485),
.A3(net10986),
.ZN(net6503)
);

DFFRS_X1 c6106(
.D(net5502),
.RN(net6483),
.SN(net6500),
.CK(clk),
.Q(net6505),
.QN(net6504)
);

XOR2_X1 c6107(
.A(net6487),
.B(net10657),
.Z(net6506)
);

NOR2_X1 c6108(
.A1(net6470),
.A2(net11353),
.ZN(net6507)
);

OR2_X2 c6109(
.A1(net2629),
.A2(net6507),
.ZN(net6508)
);

NOR2_X4 c6110(
.A1(net4573),
.A2(net6493),
.ZN(net6509)
);

NOR2_X2 c6111(
.A1(net6507),
.A2(net10803),
.ZN(net6510)
);

XOR2_X2 c6112(
.A(net6470),
.B(net5454),
.Z(net6511)
);

XNOR2_X1 c6113(
.A(net6501),
.B(net6482),
.ZN(net6512)
);

INV_X32 c6114(
.A(net10174),
.ZN(net6513)
);

OR2_X4 c6115(
.A1(net6502),
.A2(net6510),
.ZN(net6514)
);

OR2_X1 c6116(
.A1(net2582),
.A2(net6445),
.ZN(net6515)
);

OR3_X4 c6117(
.A1(net6511),
.A2(net5508),
.A3(net6162),
.ZN(net6516)
);

OAI222_X2 c6118(
.A1(net6503),
.A2(net6162),
.B1(net6475),
.B2(net5423),
.C1(net5413),
.C2(net6486),
.ZN(net6517)
);

XNOR2_X2 c6119(
.A(net6490),
.B(net6474),
.ZN(net6518)
);

DFFRS_X2 c6120(
.D(net6512),
.RN(net6459),
.SN(net5511),
.CK(clk),
.Q(net6520),
.QN(net6519)
);

NAND4_X1 c6121(
.A1(net6465),
.A2(net6518),
.A3(net6517),
.A4(net6519),
.ZN(net6521)
);

AOI222_X1 c6122(
.A1(net6518),
.A2(net6485),
.B1(net6504),
.B2(net6493),
.C1(net5556),
.C2(net6423),
.ZN(net6522)
);

AND3_X2 c6123(
.A1(net5424),
.A2(net6507),
.A3(net10823),
.ZN(net6523)
);

NOR3_X1 c6124(
.A1(net6393),
.A2(net6484),
.A3(net6510),
.ZN(net6524)
);

INV_X4 c6125(
.A(net11265),
.ZN(net6525)
);

AND2_X4 c6126(
.A1(net6510),
.A2(net6501),
.ZN(net6526)
);

OR4_X1 c6127(
.A1(net5389),
.A2(net3582),
.A3(net5557),
.A4(net11451),
.ZN(net6527)
);

OR3_X2 c6128(
.A1(net6526),
.A2(net6510),
.A3(net10656),
.ZN(net6528)
);

OAI21_X2 c6129(
.A(net6517),
.B1(net6520),
.B2(net6507),
.ZN(net6529)
);

OAI21_X1 c6130(
.A(net6526),
.B1(net4392),
.B2(net10987),
.ZN(net6530)
);

AND2_X1 c6131(
.A1(net6505),
.A2(net11081),
.ZN(net6531)
);

AOI21_X2 c6132(
.A(net6405),
.B1(net6507),
.B2(net6531),
.ZN(net6532)
);

OAI221_X4 c6133(
.A(net6093),
.B1(net6487),
.B2(net6510),
.C1(net6531),
.C2(net6462),
.ZN(net6533)
);

NAND2_X1 c6134(
.A1(net6505),
.A2(net6457),
.ZN(net6534)
);

INV_X1 c6135(
.A(net10476),
.ZN(net6535)
);

INV_X2 c6136(
.A(net10102),
.ZN(net6536)
);

AOI21_X1 c6137(
.A(net6487),
.B1(net6531),
.B2(net6510),
.ZN(net6537)
);

SDFF_X1 c6138(
.D(net6536),
.SE(net6537),
.SI(net4542),
.CK(clk),
.Q(net6539),
.QN(net6538)
);

AOI21_X4 c6139(
.A(net6387),
.B1(net6513),
.B2(net6494),
.ZN(net6540)
);

AND3_X1 c6140(
.A1(net6488),
.A2(net6539),
.A3(net6531),
.ZN(net6541)
);

SDFF_X2 c6141(
.D(net6540),
.SE(net6534),
.SI(net6531),
.CK(clk),
.Q(net6543),
.QN(net6542)
);

INV_X8 c6142(
.A(net11400),
.ZN(net6544)
);

INV_X16 c6143(
.A(net5565),
.ZN(net6545)
);

INV_X32 c6144(
.A(net10426),
.ZN(net6546)
);

INV_X4 c6145(
.A(net11484),
.ZN(net6547)
);

INV_X1 c6146(
.A(net9881),
.ZN(net6548)
);

NAND2_X2 c6147(
.A1(net5353),
.A2(net6547),
.ZN(net6549)
);

INV_X2 c6148(
.A(net5647),
.ZN(net6550)
);

NAND2_X4 c6149(
.A1(net4608),
.A2(net5574),
.ZN(net6551)
);

INV_X8 c6150(
.A(net10979),
.ZN(net6552)
);

AND2_X2 c6151(
.A1(net5427),
.A2(net10920),
.ZN(net6553)
);

INV_X16 c6152(
.A(net5511),
.ZN(net6554)
);

XOR2_X1 c6153(
.A(net5228),
.B(net6547),
.Z(net6555)
);

DFFR_X2 c6154(
.D(net5637),
.RN(net5586),
.CK(clk),
.Q(net6557),
.QN(net6556)
);

INV_X32 c6155(
.A(net9747),
.ZN(net6558)
);

NOR2_X1 c6156(
.A1(net6471),
.A2(net5557),
.ZN(net6559)
);

OR2_X2 c6157(
.A1(net6557),
.A2(net10953),
.ZN(net6560)
);

NOR2_X4 c6158(
.A1(net5576),
.A2(net4608),
.ZN(net6561)
);

NOR2_X2 c6159(
.A1(net6543),
.A2(net4488),
.ZN(net6562)
);

INV_X4 c6160(
.A(net9999),
.ZN(net6563)
);

XOR2_X2 c6161(
.A(net6018),
.B(net5562),
.Z(net6564)
);

XNOR2_X1 c6162(
.A(net5595),
.B(net4442),
.ZN(net6565)
);

OR2_X4 c6163(
.A1(net6530),
.A2(net5448),
.ZN(net6566)
);

INV_X1 c6164(
.A(net10095),
.ZN(net6567)
);

INV_X2 c6165(
.A(net9747),
.ZN(net6568)
);

OR2_X1 c6166(
.A1(net5427),
.A2(net6548),
.ZN(net6569)
);

XNOR2_X2 c6167(
.A(net6549),
.B(net5634),
.ZN(net6570)
);

AND2_X4 c6168(
.A1(net5581),
.A2(net6556),
.ZN(net6571)
);

AND2_X1 c6169(
.A1(net6562),
.A2(net6553),
.ZN(net6572)
);

NAND2_X1 c6170(
.A1(net6162),
.A2(net5601),
.ZN(net6573)
);

INV_X8 c6171(
.A(net5448),
.ZN(net6574)
);

NAND2_X2 c6172(
.A1(net4636),
.A2(net6551),
.ZN(net6575)
);

INV_X16 c6173(
.A(net11382),
.ZN(net6576)
);

INV_X32 c6174(
.A(net4442),
.ZN(net6577)
);

NAND2_X4 c6175(
.A1(net6463),
.A2(net5602),
.ZN(net6578)
);

OAI221_X2 c6176(
.A(net6546),
.B1(net6547),
.B2(net6548),
.C1(net6418),
.C2(net11400),
.ZN(net6579)
);

AND2_X2 c6177(
.A1(net3668),
.A2(net6577),
.ZN(net6580)
);

XOR2_X1 c6178(
.A(net6576),
.B(net5565),
.Z(net6581)
);

NOR2_X1 c6179(
.A1(net5612),
.A2(net4091),
.ZN(net6582)
);

OR2_X2 c6180(
.A1(net6582),
.A2(net5510),
.ZN(net6583)
);

NAND3_X1 c6181(
.A1(net6575),
.A2(net6565),
.A3(net5615),
.ZN(net6584)
);

INV_X4 c6182(
.A(net6551),
.ZN(net6585)
);

NOR2_X4 c6183(
.A1(net6580),
.A2(net4604),
.ZN(net6586)
);

NOR2_X2 c6184(
.A1(net4655),
.A2(net6584),
.ZN(net6587)
);

INV_X1 c6185(
.A(net6464),
.ZN(net6588)
);

XOR2_X2 c6186(
.A(net6568),
.B(net5353),
.Z(net6589)
);

XNOR2_X1 c6187(
.A(net3675),
.B(net6576),
.ZN(net6590)
);

NOR3_X4 c6188(
.A1(net6578),
.A2(net6543),
.A3(net6556),
.ZN(net6591)
);

NOR3_X2 c6189(
.A1(net6544),
.A2(net6567),
.A3(net11412),
.ZN(net6592)
);

OR2_X4 c6190(
.A1(net6564),
.A2(net6582),
.ZN(net6593)
);

OR2_X1 c6191(
.A1(net6577),
.A2(net6592),
.ZN(net6594)
);

XNOR2_X2 c6192(
.A(net6585),
.B(net6592),
.ZN(net6595)
);

AND2_X4 c6193(
.A1(net6461),
.A2(net5564),
.ZN(net6596)
);

AND2_X1 c6194(
.A1(net6508),
.A2(net6569),
.ZN(net6597)
);

INV_X2 c6195(
.A(net6563),
.ZN(net6598)
);

INV_X8 c6196(
.A(net10125),
.ZN(net6599)
);

NAND2_X1 c6197(
.A1(net6589),
.A2(net6571),
.ZN(net6600)
);

NAND2_X2 c6198(
.A1(net6572),
.A2(net6538),
.ZN(net6601)
);

INV_X16 c6199(
.A(net11404),
.ZN(net6602)
);

AND3_X4 c6200(
.A1(net6601),
.A2(net6602),
.A3(net6486),
.ZN(net6603)
);

NAND2_X4 c6201(
.A1(net6581),
.A2(net6602),
.ZN(net6604)
);

NAND3_X2 c6202(
.A1(net6552),
.A2(net6589),
.A3(net5637),
.ZN(net6605)
);

INV_X32 c6203(
.A(net11390),
.ZN(net6606)
);

AND2_X2 c6204(
.A1(net6588),
.A2(net6544),
.ZN(net6607)
);

XOR2_X1 c6205(
.A(net6594),
.B(net6397),
.Z(net6608)
);

OR3_X1 c6206(
.A1(net6560),
.A2(net6600),
.A3(net6578),
.ZN(net6609)
);

NOR2_X1 c6207(
.A1(net6557),
.A2(net6508),
.ZN(net6610)
);

OR2_X2 c6208(
.A1(net6597),
.A2(net6551),
.ZN(net6611)
);

NOR2_X4 c6209(
.A1(net6604),
.A2(net6585),
.ZN(net6612)
);

MUX2_X1 c6210(
.A(net6598),
.B(net6600),
.S(net6602),
.Z(net6613)
);

NOR2_X2 c6211(
.A1(net6606),
.A2(net6597),
.ZN(net6614)
);

OAI21_X4 c6212(
.A(net6613),
.B1(net6602),
.B2(net10810),
.ZN(net6615)
);

MUX2_X2 c6213(
.A(net6539),
.B(net6607),
.S(net6050),
.Z(net6616)
);

AOI222_X4 c6214(
.A1(net6584),
.A2(net6613),
.B1(net6569),
.B2(net6162),
.C1(net2605),
.C2(net5615),
.ZN(net6617)
);

NAND3_X4 c6215(
.A1(net6613),
.A2(net6615),
.A3(net6600),
.ZN(net6618)
);

OR3_X4 c6216(
.A1(net6500),
.A2(net6461),
.A3(net6592),
.ZN(net6619)
);

AND3_X2 c6217(
.A1(net6371),
.A2(net6589),
.A3(net6566),
.ZN(net6620)
);

NOR3_X1 c6218(
.A1(net6610),
.A2(net1730),
.A3(net11491),
.ZN(net6621)
);

OR3_X2 c6219(
.A1(net6595),
.A2(net6612),
.A3(net6616),
.ZN(net6622)
);

OAI33_X1 c6220(
.A1(net6618),
.A2(net6597),
.A3(net6615),
.B1(net6533),
.B2(net6607),
.B3(net6548),
.ZN(net6623)
);

AOI222_X2 c6221(
.A1(net6620),
.A2(net6565),
.B1(net6486),
.B2(net6545),
.C1(net11491),
.C2(net11552),
.ZN(net6624)
);

OAI21_X2 c6222(
.A(net6614),
.B1(net6577),
.B2(net11552),
.ZN(net6625)
);

OAI21_X1 c6223(
.A(net6621),
.B1(net6624),
.B2(net11553),
.ZN(net6626)
);

AOI21_X2 c6224(
.A(net6602),
.B1(net6625),
.B2(net11553),
.ZN(net6627)
);

AOI21_X1 c6225(
.A(net5721),
.B1(net3750),
.B2(net5705),
.ZN(net6628)
);

XOR2_X2 c6226(
.A(net2713),
.B(net6628),
.Z(net6629)
);

XNOR2_X1 c6227(
.A(net5644),
.B(net5414),
.ZN(net6630)
);

INV_X4 c6228(
.A(net10498),
.ZN(net6631)
);

INV_X1 c6229(
.A(net5699),
.ZN(net6632)
);

OR2_X4 c6230(
.A1(net4664),
.A2(net5562),
.ZN(net6633)
);

INV_X2 c6231(
.A(net9766),
.ZN(net6634)
);

OR2_X1 c6232(
.A1(net5563),
.A2(out1),
.ZN(net6635)
);

INV_X8 c6233(
.A(net11227),
.ZN(net6636)
);

INV_X16 c6234(
.A(net9833),
.ZN(net6637)
);

INV_X32 c6235(
.A(net6050),
.ZN(net6638)
);

XNOR2_X2 c6236(
.A(net6633),
.B(net6548),
.ZN(net6639)
);

AND2_X4 c6237(
.A1(net5375),
.A2(net6545),
.ZN(net6640)
);

AND2_X1 c6238(
.A1(net6565),
.A2(net5662),
.ZN(net6641)
);

NAND2_X1 c6239(
.A1(net6634),
.A2(net6632),
.ZN(net6642)
);

NAND2_X2 c6240(
.A1(net4592),
.A2(net11412),
.ZN(net6643)
);

INV_X4 c6241(
.A(net9952),
.ZN(net6644)
);

INV_X1 c6242(
.A(net3707),
.ZN(net6645)
);

NAND2_X4 c6243(
.A1(net3775),
.A2(net4742),
.ZN(net6646)
);

DFFRS_X1 c6244(
.D(net5605),
.RN(net5699),
.SN(net6462),
.CK(clk),
.Q(net6648),
.QN(net6647)
);

INV_X2 c6245(
.A(net9767),
.ZN(net6649)
);

INV_X8 c6246(
.A(net6574),
.ZN(net6650)
);

AND2_X2 c6247(
.A1(net6554),
.A2(net6632),
.ZN(net6651)
);

XOR2_X1 c6248(
.A(net6644),
.B(net4719),
.Z(net6652)
);

INV_X16 c6249(
.A(net10179),
.ZN(net6653)
);

NOR2_X1 c6250(
.A1(net5733),
.A2(net6643),
.ZN(net6654)
);

OR2_X2 c6251(
.A1(net6634),
.A2(out0),
.ZN(net6655)
);

NOR2_X4 c6252(
.A1(net6621),
.A2(net6545),
.ZN(net6656)
);

INV_X32 c6253(
.A(net10033),
.ZN(net6657)
);

NOR2_X2 c6254(
.A1(net5656),
.A2(net6644),
.ZN(net6658)
);

AOI21_X4 c6255(
.A(net6656),
.B1(net6658),
.B2(net6647),
.ZN(net6659)
);

XOR2_X2 c6256(
.A(net6647),
.B(net11451),
.Z(net6660)
);

AND3_X1 c6257(
.A1(net6659),
.A2(net6651),
.A3(net5605),
.ZN(net6661)
);

INV_X4 c6258(
.A(net6592),
.ZN(net6662)
);

XNOR2_X1 c6259(
.A(net6652),
.B(net6558),
.ZN(net6663)
);

SDFFRS_X2 c6260(
.D(net6357),
.RN(net5669),
.SE(net6639),
.SI(net6644),
.SN(net5704),
.CK(clk),
.Q(net6665),
.QN(net6664)
);

OR2_X4 c6261(
.A1(net5678),
.A2(net4702),
.ZN(net6666)
);

OR2_X1 c6262(
.A1(net5602),
.A2(net5699),
.ZN(net6667)
);

INV_X1 c6263(
.A(net6497),
.ZN(net6668)
);

XNOR2_X2 c6264(
.A(net6650),
.B(net5707),
.ZN(net6669)
);

INV_X2 c6265(
.A(net6639),
.ZN(net6670)
);

DFFRS_X2 c6266(
.D(net6663),
.RN(net6639),
.SN(net6545),
.CK(clk),
.Q(net6672),
.QN(net6671)
);

NAND3_X1 c6267(
.A1(net5683),
.A2(net3775),
.A3(net5706),
.ZN(net6673)
);

AND2_X4 c6268(
.A1(net6599),
.A2(net6635),
.ZN(net6674)
);

AND2_X1 c6269(
.A1(net6658),
.A2(net6674),
.ZN(net6675)
);

INV_X8 c6270(
.A(net9807),
.ZN(net6676)
);

INV_X16 c6271(
.A(net6571),
.ZN(net6677)
);

SDFF_X1 c6272(
.D(net5693),
.SE(net6670),
.SI(net6677),
.CK(clk),
.Q(net6679),
.QN(net6678)
);

INV_X32 c6273(
.A(net11455),
.ZN(net6680)
);

NAND2_X1 c6274(
.A1(net6666),
.A2(net6644),
.ZN(net6681)
);

INV_X4 c6275(
.A(net10096),
.ZN(net6682)
);

NAND2_X2 c6276(
.A1(net6641),
.A2(net6639),
.ZN(net6683)
);

AOI221_X4 c6277(
.A(net4595),
.B1(net6514),
.B2(net5704),
.C1(net4588),
.C2(net6548),
.ZN(net6684)
);

NAND2_X4 c6278(
.A1(net6662),
.A2(net6681),
.ZN(net6685)
);

NOR3_X4 c6279(
.A1(net4703),
.A2(net6685),
.A3(net5683),
.ZN(net6686)
);

AND2_X2 c6280(
.A1(net6667),
.A2(net6566),
.ZN(net6687)
);

XOR2_X1 c6281(
.A(net2799),
.B(net10633),
.Z(net6688)
);

NOR3_X2 c6282(
.A1(net6624),
.A2(net6687),
.A3(net5701),
.ZN(net6689)
);

INV_X1 c6283(
.A(net10214),
.ZN(net6690)
);

NOR2_X1 c6284(
.A1(net4719),
.A2(net6641),
.ZN(net6691)
);

AND3_X4 c6285(
.A1(net6691),
.A2(net6650),
.A3(net6624),
.ZN(net6692)
);

OR2_X2 c6286(
.A1(net10616),
.A2(net11341),
.ZN(net6693)
);

NOR2_X4 c6287(
.A1(net6671),
.A2(net10824),
.ZN(net6694)
);

AOI221_X2 c6288(
.A(net5692),
.B1(net6495),
.B2(net3775),
.C1(net6632),
.C2(net6569),
.ZN(net6695)
);

NOR2_X2 c6289(
.A1(net5727),
.A2(net11046),
.ZN(net6696)
);

NAND3_X2 c6290(
.A1(net6672),
.A2(net6685),
.A3(net6639),
.ZN(net6697)
);

INV_X2 c6291(
.A(net9908),
.ZN(net6698)
);

OR3_X1 c6292(
.A1(net6637),
.A2(net6678),
.A3(net11341),
.ZN(net6699)
);

INV_X8 c6293(
.A(net10372),
.ZN(net6700)
);

XOR2_X2 c6294(
.A(net6680),
.B(net6690),
.Z(net6701)
);

MUX2_X1 c6295(
.A(net6627),
.B(net6699),
.S(net6682),
.Z(net6702)
);

OAI21_X4 c6296(
.A(net6699),
.B1(net6664),
.B2(net5716),
.ZN(net6703)
);

AOI221_X1 c6297(
.A(net6653),
.B1(net6694),
.B2(net5739),
.C1(net5689),
.C2(net5729),
.ZN(net6704)
);

MUX2_X2 c6298(
.A(net4740),
.B(net6666),
.S(net11120),
.Z(net6705)
);

SDFF_X2 c6299(
.D(net6705),
.SE(net6697),
.SI(net6703),
.CK(clk),
.Q(net6707),
.QN(net6706)
);

OAI22_X1 c6300(
.A1(net6676),
.A2(net5683),
.B1(net5704),
.B2(net6663),
.ZN(net6708)
);

DFFRS_X1 c6301(
.D(net6683),
.RN(net6707),
.SN(net6694),
.CK(clk),
.Q(net6710),
.QN(net6709)
);

NAND3_X4 c6302(
.A1(net6707),
.A2(net6690),
.A3(net11447),
.ZN(net6711)
);

OR3_X4 c6303(
.A1(net6586),
.A2(net6693),
.A3(net6711),
.ZN(net6712)
);

AND3_X2 c6304(
.A1(net6704),
.A2(net6703),
.A3(net6709),
.ZN(net6713)
);

NOR3_X1 c6305(
.A1(net5662),
.A2(net6713),
.A3(net6706),
.ZN(net6714)
);

INV_X16 c6306(
.A(net10271),
.ZN(net6715)
);

OR3_X2 c6307(
.A1(net6642),
.A2(net6700),
.A3(net4704),
.ZN(net6716)
);

XNOR2_X1 c6308(
.A(net5833),
.B(net6635),
.ZN(net6717)
);

AND4_X2 c6309(
.A1(net2862),
.A2(net5730),
.A3(net5833),
.A4(net3854),
.ZN(net6718)
);

OR2_X4 c6310(
.A1(net5705),
.A2(net10631),
.ZN(net6719)
);

OR2_X1 c6311(
.A1(net5749),
.A2(net4776),
.ZN(net6720)
);

OAI21_X2 c6312(
.A(net4812),
.B1(net6701),
.B2(net5784),
.ZN(net6721)
);

XNOR2_X2 c6313(
.A(net5822),
.B(net5833),
.ZN(net6722)
);

OAI21_X1 c6314(
.A(net3855),
.B1(net4784),
.B2(net5826),
.ZN(net6723)
);

AND2_X4 c6315(
.A1(net3833),
.A2(net5821),
.ZN(net6724)
);

AND2_X1 c6316(
.A1(net5782),
.A2(net5777),
.ZN(net6725)
);

INV_X32 c6317(
.A(net9802),
.ZN(out3)
);

NAND2_X1 c6318(
.A1(net5740),
.A2(net11544),
.ZN(net6726)
);

DFFRS_X2 c6319(
.D(net6561),
.RN(net6722),
.SN(net5759),
.CK(clk),
.Q(net6728),
.QN(net6727)
);

NAND2_X2 c6320(
.A1(net6628),
.A2(net6727),
.ZN(net6729)
);

SDFF_X1 c6321(
.D(net6721),
.SE(net6725),
.SI(net6674),
.CK(clk),
.Q(net6731),
.QN(net6730)
);

AOI21_X2 c6322(
.A(net6635),
.B1(net5616),
.B2(net3859),
.ZN(net6732)
);

NAND2_X4 c6323(
.A1(net5797),
.A2(net4784),
.ZN(net6733)
);

INV_X4 c6324(
.A(net9801),
.ZN(net6734)
);

AOI21_X1 c6325(
.A(net6674),
.B1(net5705),
.B2(net5740),
.ZN(net6735)
);

AND2_X2 c6326(
.A1(net5816),
.A2(net6728),
.ZN(net6736)
);

SDFF_X2 c6327(
.D(net6723),
.SE(net6648),
.SI(net6734),
.CK(clk),
.Q(net6738),
.QN(net6737)
);

AOI21_X4 c6328(
.A(net5777),
.B1(net6635),
.B2(net4764),
.ZN(net6739)
);

XOR2_X1 c6329(
.A(net5758),
.B(net11089),
.Z(net6740)
);

DFFRS_X1 c6330(
.D(net3859),
.RN(net4837),
.SN(net6195),
.CK(clk),
.Q(net6742),
.QN(net6741)
);

AND3_X1 c6331(
.A1(net5745),
.A2(net1857),
.A3(net5708),
.ZN(net6743)
);

SDFFS_X2 c6332(
.D(net6724),
.SE(net6665),
.SI(net6743),
.SN(net5545),
.CK(clk),
.Q(net6745),
.QN(net6744)
);

NAND3_X1 c6333(
.A1(net5770),
.A2(net6737),
.A3(net6714),
.ZN(net6746)
);

NOR3_X4 c6334(
.A1(net5590),
.A2(net3878),
.A3(net6545),
.ZN(net6747)
);

NOR3_X2 c6335(
.A1(net6740),
.A2(net5832),
.A3(net2843),
.ZN(net6748)
);

NOR2_X1 c6336(
.A1(net4823),
.A2(net4846),
.ZN(net6749)
);

AND3_X4 c6337(
.A1(net6742),
.A2(net6717),
.A3(net4776),
.ZN(net6750)
);

NAND3_X2 c6338(
.A1(net6677),
.A2(net4784),
.A3(net5782),
.ZN(net6751)
);

OR2_X2 c6339(
.A1(net6462),
.A2(net6742),
.ZN(net6752)
);

AND4_X1 c6340(
.A1(net5708),
.A2(net6742),
.A3(net4764),
.A4(net6701),
.ZN(net6753)
);

OR3_X1 c6341(
.A1(net6718),
.A2(net6690),
.A3(net5753),
.ZN(net6754)
);

MUX2_X1 c6342(
.A(net5758),
.B(net5810),
.S(net5754),
.Z(net6755)
);

AOI22_X4 c6343(
.A1(net6738),
.A2(net4856),
.B1(net6749),
.B2(net5791),
.ZN(net6756)
);

OAI21_X4 c6344(
.A(net6753),
.B1(net6749),
.B2(net10777),
.ZN(net6757)
);

INV_X1 c6345(
.A(net11455),
.ZN(net6758)
);

MUX2_X2 c6346(
.A(net4776),
.B(net6674),
.S(net5759),
.Z(net6759)
);

NAND3_X4 c6347(
.A1(net6747),
.A2(net6739),
.A3(net5650),
.ZN(net6760)
);

OR3_X4 c6348(
.A1(net5794),
.A2(net6749),
.A3(net3859),
.ZN(net6761)
);

AND3_X2 c6349(
.A1(net5760),
.A2(net6740),
.A3(net11137),
.ZN(net6762)
);

INV_X2 c6350(
.A(net10027),
.ZN(net6763)
);

NOR3_X1 c6351(
.A1(net5824),
.A2(net6701),
.A3(net6732),
.ZN(net6764)
);

OR3_X2 c6352(
.A1(net5811),
.A2(net6757),
.A3(net5650),
.ZN(net6765)
);

OAI21_X2 c6353(
.A(net6669),
.B1(net6749),
.B2(net4843),
.ZN(net6766)
);

NOR2_X4 c6354(
.A1(net3820),
.A2(net6749),
.ZN(net6767)
);

OAI21_X1 c6355(
.A(net6761),
.B1(net6725),
.B2(net6762),
.ZN(net6768)
);

NOR2_X2 c6356(
.A1(net6583),
.A2(net5827),
.ZN(net6769)
);

AOI21_X2 c6357(
.A(net6761),
.B1(net6769),
.B2(net10945),
.ZN(net6770)
);

XOR2_X2 c6358(
.A(net6630),
.B(net6738),
.Z(net6771)
);

AOI21_X1 c6359(
.A(net5761),
.B1(net6669),
.B2(net10870),
.ZN(net6772)
);

OAI221_X1 c6360(
.A(net6771),
.B1(net5708),
.B2(net6607),
.C1(net6762),
.C2(net10679),
.ZN(net6773)
);

AOI21_X4 c6361(
.A(net5784),
.B1(net6753),
.B2(net5580),
.ZN(net6774)
);

AND3_X1 c6362(
.A1(net6767),
.A2(net6755),
.A3(net4704),
.ZN(net6775)
);

NAND3_X1 c6363(
.A1(net6726),
.A2(net5827),
.A3(net6741),
.ZN(net6776)
);

NOR3_X4 c6364(
.A1(net6722),
.A2(net6756),
.A3(net4844),
.ZN(net6777)
);

NOR3_X2 c6365(
.A1(net6773),
.A2(net5796),
.A3(net6669),
.ZN(net6778)
);

AND3_X4 c6366(
.A1(net6774),
.A2(net6753),
.A3(net6730),
.ZN(net6779)
);

NAND3_X2 c6367(
.A1(net6776),
.A2(net6719),
.A3(net5590),
.ZN(net6780)
);

OR3_X1 c6368(
.A1(net5819),
.A2(net6779),
.A3(net6729),
.ZN(net6781)
);

MUX2_X1 c6369(
.A(net6701),
.B(net6779),
.S(net6762),
.Z(net6782)
);

OAI22_X4 c6370(
.A1(net2844),
.A2(net5816),
.B1(net6741),
.B2(net6761),
.ZN(net6783)
);

OAI21_X4 c6371(
.A(net6763),
.B1(net6781),
.B2(net6769),
.ZN(net6784)
);

DFFRS_X2 c6372(
.D(net6781),
.RN(net5708),
.SN(net6714),
.CK(clk),
.Q(net6786),
.QN(net6785)
);

MUX2_X2 c6373(
.A(net4844),
.B(net6740),
.S(net10937),
.Z(net6787)
);

SDFF_X1 c6374(
.D(net6729),
.SE(net6764),
.SI(net6744),
.CK(clk),
.Q(net6789),
.QN(net6788)
);

NAND3_X4 c6375(
.A1(net6695),
.A2(net6761),
.A3(net4764),
.ZN(net6790)
);

OR3_X4 c6376(
.A1(net6545),
.A2(net6772),
.A3(net6779),
.ZN(net6791)
);

AND3_X2 c6377(
.A1(net6787),
.A2(net6769),
.A3(net6775),
.ZN(net6792)
);

NOR3_X1 c6378(
.A1(net6751),
.A2(net5553),
.A3(net6769),
.ZN(net6793)
);

OR3_X2 c6379(
.A1(net6775),
.A2(net6749),
.A3(net6785),
.ZN(net6794)
);

OAI21_X2 c6380(
.A(net6794),
.B1(net5748),
.B2(net10938),
.ZN(net6795)
);

SDFF_X2 c6381(
.D(net6725),
.SE(net6792),
.SI(net6774),
.CK(clk),
.Q(net6797),
.QN(net6796)
);

OAI21_X1 c6382(
.A(net5764),
.B1(net6665),
.B2(net6677),
.ZN(net6798)
);

AOI21_X2 c6383(
.A(net6786),
.B1(net6791),
.B2(net11067),
.ZN(net6799)
);

DFFRS_X1 c6384(
.D(net6797),
.RN(net6799),
.SN(net10678),
.CK(clk),
.Q(net6801),
.QN(net6800)
);

AOI22_X2 c6385(
.A1(net6791),
.A2(net6777),
.B1(net6796),
.B2(net4837),
.ZN(net6802)
);

NAND4_X4 c6386(
.A1(net6745),
.A2(net6798),
.A3(net6763),
.A4(net6732),
.ZN(net6803)
);

OAI221_X4 c6387(
.A(net6736),
.B1(net6745),
.B2(net6803),
.C1(net6694),
.C2(net11035),
.ZN(net6804)
);

OAI211_X2 c6388(
.A(net6714),
.B(net6794),
.C1(net6761),
.C2(net10753),
.ZN(net6805)
);

OR4_X2 c6389(
.A1(net6799),
.A2(net6758),
.A3(net3829),
.A4(net6803),
.ZN(net6806)
);

OAI221_X2 c6390(
.A(net4764),
.B1(net6771),
.B2(net6740),
.C1(net1731),
.C2(net10838),
.ZN(net6807)
);

INV_X8 c6391(
.A(net3936),
.ZN(net6808)
);

INV_X16 c6392(
.A(net9737),
.ZN(net6809)
);

INV_X32 c6393(
.A(net4935),
.ZN(net6810)
);

XNOR2_X1 c6394(
.A(net5869),
.B(net4910),
.ZN(net6811)
);

INV_X4 c6395(
.A(net3968),
.ZN(net6812)
);

INV_X1 c6396(
.A(net4910),
.ZN(net6813)
);

INV_X2 c6397(
.A(net3916),
.ZN(net6814)
);

DFFS_X1 c6398(
.D(net6808),
.SN(net5838),
.CK(clk),
.Q(net6816),
.QN(net6815)
);

OR2_X4 c6399(
.A1(net4894),
.A2(net5839),
.ZN(net6817)
);

INV_X8 c6400(
.A(net1009),
.ZN(net6818)
);

INV_X16 c6401(
.A(net4869),
.ZN(net6819)
);

INV_X32 c6402(
.A(net1951),
.ZN(net6820)
);

INV_X4 c6403(
.A(net5857),
.ZN(net6821)
);

INV_X1 c6404(
.A(net6819),
.ZN(net6822)
);

INV_X2 c6405(
.A(net4894),
.ZN(net6823)
);

INV_X8 c6406(
.A(net5840),
.ZN(net6824)
);

INV_X16 c6407(
.A(net3955),
.ZN(net6825)
);

INV_X32 c6408(
.A(net6814),
.ZN(net6826)
);

INV_X4 c6409(
.A(net5847),
.ZN(net6827)
);

INV_X1 c6410(
.A(net4863),
.ZN(net6828)
);

OR2_X1 c6411(
.A1(net3912),
.A2(net11549),
.ZN(net6829)
);

INV_X2 c6412(
.A(net6820),
.ZN(net6830)
);

INV_X8 c6413(
.A(net2964),
.ZN(net6831)
);

XNOR2_X2 c6414(
.A(net5870),
.B(net5857),
.ZN(net6832)
);

INV_X16 c6415(
.A(net6827),
.ZN(net6833)
);

INV_X32 c6416(
.A(net9736),
.ZN(net6834)
);

INV_X4 c6417(
.A(net9830),
.ZN(net6835)
);

AND2_X4 c6418(
.A1(net6834),
.A2(net6818),
.ZN(net6836)
);

INV_X1 c6419(
.A(net9852),
.ZN(net6837)
);

INV_X2 c6420(
.A(net6836),
.ZN(net6838)
);

AND2_X1 c6421(
.A1(net6823),
.A2(net5924),
.ZN(net6839)
);

NAND2_X1 c6422(
.A1(net3968),
.A2(net5911),
.ZN(net6840)
);

NAND2_X2 c6423(
.A1(net5891),
.A2(net3936),
.ZN(net6841)
);

NAND2_X4 c6424(
.A1(net6812),
.A2(net6815),
.ZN(net6842)
);

AND2_X2 c6425(
.A1(net6829),
.A2(net4869),
.ZN(net6843)
);

INV_X8 c6426(
.A(net6842),
.ZN(net6844)
);

INV_X16 c6427(
.A(net6818),
.ZN(net6845)
);

XOR2_X1 c6428(
.A(net6845),
.B(net6842),
.Z(net6846)
);

NOR2_X1 c6429(
.A1(net6846),
.A2(net3968),
.ZN(net6847)
);

OR2_X2 c6430(
.A1(net6843),
.A2(net6844),
.ZN(net6848)
);

INV_X32 c6431(
.A(net9851),
.ZN(net6849)
);

NOR2_X4 c6432(
.A1(net4871),
.A2(net6846),
.ZN(net6850)
);

DFFS_X2 c6433(
.D(net5914),
.SN(net5916),
.CK(clk),
.Q(net6852),
.QN(net6851)
);

INV_X4 c6434(
.A(net4913),
.ZN(net6853)
);

INV_X1 c6435(
.A(net9936),
.ZN(net6854)
);

INV_X2 c6436(
.A(net9824),
.ZN(net6855)
);

DFFRS_X2 c6437(
.D(net4863),
.RN(net6826),
.SN(net6808),
.CK(clk),
.Q(net6857),
.QN(net6856)
);

INV_X8 c6438(
.A(net10553),
.ZN(net6858)
);

INV_X16 c6439(
.A(net6855),
.ZN(net6859)
);

DFFR_X1 c6440(
.D(net6850),
.RN(net2996),
.CK(clk),
.Q(net6861),
.QN(net6860)
);

DFFR_X2 c6441(
.D(net6839),
.RN(net5905),
.CK(clk),
.Q(net6863),
.QN(net6862)
);

INV_X32 c6442(
.A(net6858),
.ZN(net6864)
);

NOR2_X2 c6443(
.A1(net6817),
.A2(net6861),
.ZN(net6865)
);

AOI21_X1 c6444(
.A(net6820),
.B1(net6855),
.B2(net6859),
.ZN(net6866)
);

XOR2_X2 c6445(
.A(net6826),
.B(net6865),
.Z(net6867)
);

XNOR2_X1 c6446(
.A(net6834),
.B(net6866),
.ZN(net6868)
);

OR2_X4 c6447(
.A1(net6830),
.A2(net6866),
.ZN(net6869)
);

AOI211_X1 c6448(
.A(net6861),
.B(net6859),
.C1(net6828),
.C2(net5924),
.ZN(net6870)
);

AOI21_X4 c6449(
.A(net5891),
.B1(net6866),
.B2(net5839),
.ZN(net6871)
);

DFFS_X1 c6450(
.D(net4909),
.SN(net6870),
.CK(clk),
.Q(net6873),
.QN(net6872)
);

DFFS_X2 c6451(
.D(net6853),
.SN(net6867),
.CK(clk),
.Q(net6875),
.QN(net6874)
);

OR2_X1 c6452(
.A1(net5916),
.A2(net6856),
.ZN(net6876)
);

XNOR2_X2 c6453(
.A(net6837),
.B(net6876),
.ZN(net6877)
);

SDFF_X1 c6454(
.D(net6813),
.SE(net6867),
.SI(net6846),
.CK(clk),
.Q(net6879),
.QN(net6878)
);

AND2_X4 c6455(
.A1(net6864),
.A2(net6878),
.ZN(net6880)
);

AND2_X1 c6456(
.A1(net6828),
.A2(net6864),
.ZN(net6881)
);

NAND2_X1 c6457(
.A1(net5869),
.A2(net6850),
.ZN(net6882)
);

NAND2_X2 c6458(
.A1(net5911),
.A2(net6880),
.ZN(net6883)
);

AND3_X1 c6459(
.A1(net6879),
.A2(net4874),
.A3(net10553),
.ZN(net6884)
);

NAND2_X4 c6460(
.A1(net6879),
.A2(net6860),
.ZN(net6885)
);

AND2_X2 c6461(
.A1(net6859),
.A2(net5919),
.ZN(net6886)
);

SDFF_X2 c6462(
.D(net6881),
.SE(net6832),
.SI(net6872),
.CK(clk),
.Q(net6888),
.QN(net6887)
);

OAI222_X1 c6463(
.A1(net6871),
.A2(net6833),
.B1(net6887),
.B2(net6808),
.C1(net6870),
.C2(net5924),
.ZN(net6889)
);

NAND3_X1 c6464(
.A1(net6825),
.A2(net6828),
.A3(net6877),
.ZN(net6890)
);

NOR3_X4 c6465(
.A1(net6880),
.A2(net5859),
.A3(net6883),
.ZN(net6891)
);

NOR3_X2 c6466(
.A1(net6854),
.A2(net6887),
.A3(net5839),
.ZN(net6892)
);

AND3_X4 c6467(
.A1(net6869),
.A2(net6836),
.A3(net6862),
.ZN(net6893)
);

NAND3_X2 c6468(
.A1(net6893),
.A2(net6890),
.A3(net11555),
.ZN(net6894)
);

OAI222_X4 c6469(
.A1(net6865),
.A2(net6894),
.B1(net6870),
.B2(net6872),
.C1(net5924),
.C2(net6812),
.ZN(net6895)
);

DFFRS_X1 c6470(
.D(net6821),
.RN(net6892),
.SN(net11557),
.CK(clk),
.Q(net6897),
.QN(net6896)
);

NAND4_X2 c6471(
.A1(net6892),
.A2(net6877),
.A3(net6890),
.A4(net11555),
.ZN(net6898)
);

OR3_X1 c6472(
.A1(net6894),
.A2(net6890),
.A3(net11556),
.ZN(net6899)
);

OR4_X4 c6473(
.A1(net6897),
.A2(net6884),
.A3(net11554),
.A4(net11556),
.ZN(net6900)
);

INV_X4 c6474(
.A(net6890),
.ZN(net6901)
);

INV_X1 c6475(
.A(net9691),
.ZN(net6902)
);

INV_X2 c6476(
.A(net5019),
.ZN(net6903)
);

INV_X8 c6477(
.A(net5988),
.ZN(net6904)
);

MUX2_X1 c6478(
.A(net5930),
.B(net5012),
.S(net3955),
.Z(net6905)
);

INV_X16 c6479(
.A(net4914),
.ZN(net6906)
);

INV_X32 c6480(
.A(net6014),
.ZN(net6907)
);

INV_X4 c6481(
.A(net4954),
.ZN(net6908)
);

INV_X1 c6482(
.A(net9692),
.ZN(net6909)
);

SDFFR_X1 c6483(
.D(net6896),
.RN(net6014),
.SE(net5883),
.SI(net4038),
.CK(clk),
.Q(net6911),
.QN(net6910)
);

INV_X2 c6484(
.A(net6843),
.ZN(net6912)
);

INV_X8 c6485(
.A(net10503),
.ZN(net6913)
);

INV_X16 c6486(
.A(net6903),
.ZN(net6914)
);

XOR2_X1 c6487(
.A(net6818),
.B(net6868),
.Z(net6915)
);

NOR2_X1 c6488(
.A1(net4975),
.A2(net5885),
.ZN(net6916)
);

INV_X32 c6489(
.A(net6002),
.ZN(net6917)
);

INV_X4 c6490(
.A(net6812),
.ZN(net6918)
);

INV_X1 c6491(
.A(net5990),
.ZN(net6919)
);

INV_X2 c6492(
.A(net6907),
.ZN(net6920)
);

INV_X8 c6493(
.A(net6915),
.ZN(net6921)
);

INV_X16 c6494(
.A(net6902),
.ZN(net6922)
);

INV_X32 c6495(
.A(net6906),
.ZN(net6923)
);

INV_X4 c6496(
.A(net6913),
.ZN(net6924)
);

OR2_X2 c6497(
.A1(net5859),
.A2(net5849),
.ZN(net6925)
);

INV_X1 c6498(
.A(net6904),
.ZN(net6926)
);

INV_X2 c6499(
.A(net6849),
.ZN(net6927)
);

NOR2_X4 c6500(
.A1(net5002),
.A2(net5955),
.ZN(net6928)
);

NOR2_X2 c6501(
.A1(net6925),
.A2(net5934),
.ZN(net6929)
);

OAI21_X4 c6502(
.A(net6824),
.B1(net6902),
.B2(net6900),
.ZN(net6930)
);

INV_X8 c6503(
.A(net6920),
.ZN(net6931)
);

INV_X16 c6504(
.A(net6909),
.ZN(net6932)
);

INV_X32 c6505(
.A(net6900),
.ZN(net6933)
);

MUX2_X2 c6506(
.A(net6877),
.B(net4984),
.S(net6917),
.Z(net6934)
);

XOR2_X2 c6507(
.A(net6912),
.B(net5859),
.Z(net6935)
);

INV_X4 c6508(
.A(net6857),
.ZN(net6936)
);

NAND3_X4 c6509(
.A1(net6918),
.A2(net6934),
.A3(net6930),
.ZN(net6937)
);

INV_X1 c6510(
.A(net6923),
.ZN(net6938)
);

XNOR2_X1 c6511(
.A(net3936),
.B(net4949),
.ZN(net6939)
);

INV_X2 c6512(
.A(net9891),
.ZN(net6940)
);

OR3_X4 c6513(
.A1(net6907),
.A2(net6925),
.A3(net6921),
.ZN(net6941)
);

OAI22_X2 c6514(
.A1(net6931),
.A2(net2995),
.B1(net5955),
.B2(net6932),
.ZN(net6942)
);

INV_X8 c6515(
.A(net6919),
.ZN(net6943)
);

OR2_X4 c6516(
.A1(net6937),
.A2(net6928),
.ZN(net6944)
);

INV_X16 c6517(
.A(net6905),
.ZN(net6945)
);

OR2_X1 c6518(
.A1(net1009),
.A2(net10617),
.ZN(net6946)
);

INV_X32 c6519(
.A(net6918),
.ZN(net6947)
);

XNOR2_X2 c6520(
.A(net4869),
.B(net6932),
.ZN(net6948)
);

AND2_X4 c6521(
.A1(net4949),
.A2(net6920),
.ZN(net6949)
);

INV_X4 c6522(
.A(net11072),
.ZN(net6950)
);

INV_X1 c6523(
.A(net10456),
.ZN(net6951)
);

AND3_X2 c6524(
.A1(net6949),
.A2(net5937),
.A3(net6948),
.ZN(net6952)
);

INV_X2 c6525(
.A(net6940),
.ZN(net6953)
);

NOR3_X1 c6526(
.A1(net6816),
.A2(net4993),
.A3(net6950),
.ZN(net6954)
);

AND2_X1 c6527(
.A1(net6868),
.A2(net10816),
.ZN(net6955)
);

NAND2_X1 c6528(
.A1(net5931),
.A2(net6932),
.ZN(net6956)
);

NAND2_X2 c6529(
.A1(net6933),
.A2(net6927),
.ZN(net6957)
);

INV_X8 c6530(
.A(net10311),
.ZN(net6958)
);

NAND2_X4 c6531(
.A1(net6932),
.A2(net6950),
.ZN(net6959)
);

SDFFR_X2 c6532(
.D(net6958),
.RN(net6942),
.SE(net6957),
.SI(net2964),
.CK(clk),
.Q(net6961),
.QN(net6960)
);

AND2_X2 c6533(
.A1(net6957),
.A2(net11557),
.ZN(net6962)
);

INV_X16 c6534(
.A(net6911),
.ZN(net6963)
);

XOR2_X1 c6535(
.A(net6946),
.B(net6962),
.Z(net6964)
);

INV_X32 c6536(
.A(net6950),
.ZN(net6965)
);

NOR2_X1 c6537(
.A1(net6962),
.A2(net4914),
.ZN(net6966)
);

OR2_X2 c6538(
.A1(net6938),
.A2(net6964),
.ZN(net6967)
);

NOR2_X4 c6539(
.A1(net6954),
.A2(net6849),
.ZN(net6968)
);

OAI211_X4 c6540(
.A(net6955),
.B(net6961),
.C1(net6912),
.C2(net6967),
.ZN(net6969)
);

AOI221_X4 c6541(
.A(net6964),
.B1(net6920),
.B2(net6950),
.C1(net6960),
.C2(net6967),
.ZN(net6970)
);

OR3_X2 c6542(
.A1(net6947),
.A2(net5935),
.A3(net6968),
.ZN(net6971)
);

INV_X4 c6543(
.A(net10053),
.ZN(net6972)
);

AOI221_X2 c6544(
.A(net6970),
.B1(net6966),
.B2(net6915),
.C1(net6967),
.C2(net6011),
.ZN(net6973)
);

DFFRS_X2 c6545(
.D(net6971),
.RN(net4949),
.SN(net6928),
.CK(clk),
.Q(net6975),
.QN(net6974)
);

OAI21_X2 c6546(
.A(net6951),
.B1(net6974),
.B2(net6959),
.ZN(net6976)
);

OAI21_X1 c6547(
.A(net5925),
.B1(net6901),
.B2(net10618),
.ZN(net6977)
);

INV_X1 c6548(
.A(net10074),
.ZN(net6978)
);

NOR2_X2 c6549(
.A1(net5996),
.A2(net6963),
.ZN(net6979)
);

XOR2_X2 c6550(
.A(net6975),
.B(net6903),
.Z(net6980)
);

XNOR2_X1 c6551(
.A(net6966),
.B(net10836),
.ZN(net6981)
);

AOI21_X2 c6552(
.A(net6926),
.B1(net6949),
.B2(net6936),
.ZN(net6982)
);

DFFR_X1 c6553(
.D(net6982),
.RN(net10730),
.CK(clk),
.Q(net6984),
.QN(net6983)
);

OR2_X4 c6554(
.A1(net6976),
.A2(net6983),
.ZN(net6985)
);

AOI221_X1 c6555(
.A(net6959),
.B1(net6978),
.B2(net6982),
.C1(net6936),
.C2(net6976),
.ZN(net6986)
);

OAI222_X2 c6556(
.A1(net6978),
.A2(net6932),
.B1(net6976),
.B2(net6985),
.C1(net6980),
.C2(net4999),
.ZN(net6987)
);

INV_X2 c6557(
.A(net6059),
.ZN(net6988)
);

INV_X8 c6558(
.A(net4902),
.ZN(net6989)
);

INV_X16 c6559(
.A(net11337),
.ZN(net6990)
);

INV_X32 c6560(
.A(net6922),
.ZN(net6991)
);

INV_X4 c6561(
.A(net10652),
.ZN(net6992)
);

OR2_X1 c6562(
.A1(net6831),
.A2(net6967),
.ZN(net6993)
);

XNOR2_X2 c6563(
.A(net6953),
.B(net6936),
.ZN(net6994)
);

AND2_X4 c6564(
.A1(net6979),
.A2(net4935),
.ZN(net6995)
);

AND2_X1 c6565(
.A1(net6956),
.A2(net6087),
.ZN(net6996)
);

INV_X1 c6566(
.A(net6075),
.ZN(net6997)
);

INV_X2 c6567(
.A(net9792),
.ZN(net6998)
);

NAND2_X1 c6568(
.A1(net5114),
.A2(net6998),
.ZN(net6999)
);

INV_X8 c6569(
.A(net11332),
.ZN(net7000)
);

INV_X16 c6570(
.A(net6997),
.ZN(net7001)
);

NAND2_X2 c6571(
.A1(net6988),
.A2(net6994),
.ZN(net7002)
);

INV_X32 c6572(
.A(net5955),
.ZN(net7003)
);

NAND2_X4 c6573(
.A1(net7003),
.A2(net10785),
.ZN(net7004)
);

AND2_X2 c6574(
.A1(net5942),
.A2(net3129),
.ZN(net7005)
);

AOI21_X1 c6575(
.A(net7005),
.B1(net7003),
.B2(net5117),
.ZN(net7006)
);

XOR2_X1 c6576(
.A(net6095),
.B(net6928),
.Z(net7007)
);

INV_X4 c6577(
.A(net5124),
.ZN(net7008)
);

AOI21_X4 c6578(
.A(net7006),
.B1(net6961),
.B2(net6989),
.ZN(net7009)
);

INV_X1 c6579(
.A(net9791),
.ZN(net7010)
);

AND3_X1 c6580(
.A1(net5117),
.A2(net7003),
.A3(net6908),
.ZN(net7011)
);

DFFR_X2 c6581(
.D(net6993),
.RN(net11248),
.CK(clk),
.Q(net7013),
.QN(net7012)
);

NAND3_X1 c6582(
.A1(net2902),
.A2(net3976),
.A3(net6968),
.ZN(net7014)
);

INV_X2 c6583(
.A(net6066),
.ZN(net7015)
);

NOR2_X1 c6584(
.A1(net4014),
.A2(net6100),
.ZN(net7016)
);

OR2_X2 c6585(
.A1(net6957),
.A2(net6956),
.ZN(net7017)
);

INV_X8 c6586(
.A(net10166),
.ZN(net7018)
);

NOR2_X4 c6587(
.A1(net6968),
.A2(net4014),
.ZN(net7019)
);

NOR2_X2 c6588(
.A1(net6090),
.A2(net7016),
.ZN(net7020)
);

INV_X16 c6589(
.A(net9823),
.ZN(net7021)
);

INV_X32 c6590(
.A(net7001),
.ZN(net7022)
);

XOR2_X2 c6591(
.A(net6020),
.B(net6097),
.Z(net7023)
);

SDFF_X1 c6592(
.D(net6028),
.SE(net6967),
.SI(net5955),
.CK(clk),
.Q(net7025),
.QN(net7024)
);

XNOR2_X1 c6593(
.A(net6930),
.B(net6994),
.ZN(net7026)
);

OR2_X4 c6594(
.A1(net7025),
.A2(net7000),
.ZN(net7027)
);

NOR3_X4 c6595(
.A1(net6065),
.A2(net6985),
.A3(net2902),
.ZN(net7028)
);

INV_X4 c6596(
.A(net11477),
.ZN(net7029)
);

OR2_X1 c6597(
.A1(net6943),
.A2(net7022),
.ZN(net7030)
);

INV_X1 c6598(
.A(net6948),
.ZN(net7031)
);

NOR3_X2 c6599(
.A1(net6099),
.A2(net6996),
.A3(net7024),
.ZN(net7032)
);

AND3_X4 c6600(
.A1(net7023),
.A2(net6994),
.A3(net11248),
.ZN(net7033)
);

INV_X2 c6601(
.A(net10049),
.ZN(net7034)
);

NAND3_X2 c6602(
.A1(net7018),
.A2(net6090),
.A3(net6987),
.ZN(net7035)
);

XNOR2_X2 c6603(
.A(net7011),
.B(net10577),
.ZN(net7036)
);

AND2_X4 c6604(
.A1(net6981),
.A2(net7004),
.ZN(net7037)
);

SDFF_X2 c6605(
.D(net6996),
.SE(net6998),
.SI(net7031),
.CK(clk),
.Q(net7039),
.QN(net7038)
);

INV_X8 c6606(
.A(net7003),
.ZN(net7040)
);

INV_X16 c6607(
.A(net11378),
.ZN(net7041)
);

INV_X32 c6608(
.A(net9803),
.ZN(net7042)
);

AND2_X1 c6609(
.A1(net7030),
.A2(net7026),
.ZN(net7043)
);

NAND2_X1 c6610(
.A1(net7033),
.A2(net7041),
.ZN(net7044)
);

INV_X4 c6611(
.A(net7026),
.ZN(net7045)
);

OR3_X1 c6612(
.A1(net6809),
.A2(net7038),
.A3(net7041),
.ZN(net7046)
);

INV_X1 c6613(
.A(net7035),
.ZN(net7047)
);

NAND2_X2 c6614(
.A1(net7018),
.A2(net10831),
.ZN(net7048)
);

NAND2_X4 c6615(
.A1(net6991),
.A2(net6094),
.ZN(net7049)
);

MUX2_X1 c6616(
.A(net7047),
.B(net4092),
.S(net7016),
.Z(net7050)
);

INV_X2 c6617(
.A(net11332),
.ZN(net7051)
);

OAI21_X4 c6618(
.A(net6091),
.B1(net7025),
.B2(net6042),
.ZN(net7052)
);

MUX2_X2 c6619(
.A(net7046),
.B(net7026),
.S(net7041),
.Z(net7053)
);

AND2_X2 c6620(
.A1(net6995),
.A2(net7049),
.ZN(net7054)
);

XOR2_X1 c6621(
.A(net7044),
.B(net6963),
.Z(net7055)
);

NOR2_X1 c6622(
.A1(net7049),
.A2(net7035),
.ZN(net7056)
);

OR2_X2 c6623(
.A1(net7031),
.A2(net6095),
.ZN(net7057)
);

OAI211_X1 c6624(
.A(net7027),
.B(net7050),
.C1(net6944),
.C2(net6870),
.ZN(net7058)
);

INV_X8 c6625(
.A(net10187),
.ZN(net7059)
);

INV_X16 c6626(
.A(net10206),
.ZN(net7060)
);

NAND3_X4 c6627(
.A1(net7043),
.A2(net7046),
.A3(net7005),
.ZN(net7061)
);

INV_X32 c6628(
.A(net10167),
.ZN(net7062)
);

DFFS_X1 c6629(
.D(net7054),
.SN(net7039),
.CK(clk),
.Q(net7064),
.QN(net7063)
);

INV_X4 c6630(
.A(net10326),
.ZN(net7065)
);

OR3_X4 c6631(
.A1(net7000),
.A2(net7064),
.A3(net5978),
.ZN(net7066)
);

AND3_X2 c6632(
.A1(net7020),
.A2(net7045),
.A3(net7052),
.ZN(net7067)
);

NOR2_X4 c6633(
.A1(net5047),
.A2(net7067),
.ZN(net7068)
);

INV_X1 c6634(
.A(net10128),
.ZN(net7069)
);

NOR3_X1 c6635(
.A1(net7060),
.A2(net7055),
.A3(net5975),
.ZN(net7070)
);

NOR2_X2 c6636(
.A1(net7069),
.A2(net7034),
.ZN(net7071)
);

DFFRS_X1 c6637(
.D(net7071),
.RN(net7036),
.SN(net7021),
.CK(clk),
.Q(net7073),
.QN(net7072)
);

XOR2_X2 c6638(
.A(net7045),
.B(net7073),
.Z(net7074)
);

AOI222_X1 c6639(
.A1(net7065),
.A2(net7061),
.B1(net7071),
.B2(net7072),
.C1(net7074),
.C2(net7012),
.ZN(net7075)
);

INV_X2 c6640(
.ZN(net7076)
);

XNOR2_X1 c6641(
.A(net6135),
.B(net6148),
.ZN(net7077)
);

OR2_X4 c6642(
.A1(net7010),
.A2(net6177),
.ZN(net7078)
);

OR2_X1 c6643(
.A1(net6130),
.A2(net7056),
.ZN(net7079)
);

XNOR2_X2 c6644(
.A(net7029),
.B(net11474),
.ZN(net7080)
);

AND2_X4 c6645(
.A1(net6101),
.A2(net6840),
.ZN(net7081)
);

AND2_X1 c6646(
.A1(net6168),
.A2(net6100),
.ZN(net7082)
);

NAND2_X1 c6647(
.A1(net5202),
.A2(net6987),
.ZN(net7083)
);

INV_X8 c6648(
.A(net11475),
.ZN(net7084)
);

NAND2_X2 c6649(
.A1(net5174),
.A2(net6124),
.ZN(net7085)
);

INV_X16 c6650(
.A(net6992),
.ZN(net7086)
);

DFFS_X2 c6651(
.D(net7077),
.SN(net6106),
.CK(clk),
.Q(net7088),
.QN(net7087)
);

INV_X32 c6652(
.A(net3223),
.ZN(net7089)
);

NAND2_X4 c6653(
.A1(net6081),
.A2(net4201),
.ZN(net7090)
);

INV_X4 c6654(
.A(net9973),
.ZN(net7091)
);

OR3_X2 c6655(
.A1(net5052),
.A2(net7067),
.A3(net3182),
.ZN(net7092)
);

AND2_X2 c6656(
.A1(net6165),
.A2(net11201),
.ZN(net7093)
);

XOR2_X1 c6657(
.A(net6148),
.B(net7079),
.Z(net7094)
);

DFFRS_X2 c6658(
.D(net6945),
.RN(net6944),
.SN(net6100),
.CK(clk),
.Q(net7096),
.QN(net7095)
);

NOR2_X1 c6659(
.A1(net7086),
.A2(net6120),
.ZN(net7097)
);

OR2_X2 c6660(
.A1(net5146),
.A2(net7011),
.ZN(net7098)
);

NOR2_X4 c6661(
.A1(net6866),
.A2(net6990),
.ZN(net7099)
);

NOR2_X2 c6662(
.A1(net6105),
.A2(net11313),
.ZN(net7100)
);

XOR2_X2 c6663(
.A(net6944),
.B(net6808),
.Z(net7101)
);

INV_X1 c6664(
.A(net11475),
.ZN(net7102)
);

INV_X2 c6665(
.A(net10122),
.ZN(net7103)
);

OAI21_X2 c6666(
.A(net6990),
.B1(net7098),
.B2(net7029),
.ZN(net7104)
);

INV_X8 c6667(
.A(net11184),
.ZN(net7105)
);

INV_X16 c6668(
.A(net6138),
.ZN(net7106)
);

XNOR2_X1 c6669(
.A(net3228),
.B(net4159),
.ZN(net7107)
);

INV_X32 c6670(
.A(net11402),
.ZN(net7108)
);

OR2_X4 c6671(
.A1(net7067),
.A2(net5174),
.ZN(net7109)
);

OR2_X1 c6672(
.A1(net6944),
.A2(net10852),
.ZN(net7110)
);

XNOR2_X2 c6673(
.A(net6087),
.B(net6965),
.ZN(net7111)
);

AND2_X4 c6674(
.A1(net7091),
.A2(net7105),
.ZN(net7112)
);

AND2_X1 c6675(
.A1(net7102),
.A2(net6168),
.ZN(net7113)
);

NAND2_X1 c6676(
.A1(net7073),
.A2(net6115),
.ZN(net7114)
);

OAI21_X1 c6677(
.A(net7022),
.B1(net7078),
.B2(net7108),
.ZN(net7115)
);

NAND2_X2 c6678(
.A1(net5849),
.A2(net7098),
.ZN(net7116)
);

NAND2_X4 c6679(
.A1(net6072),
.A2(net7081),
.ZN(net7117)
);

AOI21_X2 c6680(
.A(net6108),
.B1(net6138),
.B2(net7019),
.ZN(net7118)
);

INV_X4 c6681(
.A(net10067),
.ZN(net7119)
);

AOI21_X1 c6682(
.A(net7106),
.B1(net7082),
.B2(net7072),
.ZN(net7120)
);

AND2_X2 c6683(
.A1(net6106),
.A2(net5052),
.ZN(net7121)
);

XOR2_X1 c6684(
.A(net6035),
.B(net7080),
.Z(net7122)
);

AOI21_X4 c6685(
.A(net7089),
.B1(net6990),
.B2(net10919),
.ZN(net7123)
);

INV_X1 c6686(
.A(net10244),
.ZN(net7124)
);

NOR2_X1 c6687(
.A1(net7021),
.A2(net991),
.ZN(net7125)
);

DFFR_X1 c6688(
.D(net6965),
.RN(net7050),
.CK(clk),
.Q(net7127),
.QN(net7126)
);

INV_X2 c6689(
.A(net9972),
.ZN(net7128)
);

OR2_X2 c6690(
.A1(net7119),
.A2(net7107),
.ZN(net7129)
);

SDFF_X1 c6691(
.D(net7128),
.SE(net7122),
.SI(net11549),
.CK(clk),
.Q(net7131),
.QN(net7130)
);

NOR2_X4 c6692(
.A1(net7007),
.A2(net7063),
.ZN(net7132)
);

NOR2_X2 c6693(
.A1(net7131),
.A2(net7087),
.ZN(net7133)
);

XOR2_X2 c6694(
.A(net7108),
.B(net10734),
.Z(net7134)
);

XNOR2_X1 c6695(
.A(net7008),
.B(net7132),
.ZN(net7135)
);

OR2_X4 c6696(
.A1(net7123),
.A2(net11414),
.ZN(net7136)
);

OR2_X1 c6697(
.A1(net7134),
.A2(net7083),
.ZN(net7137)
);

SDFFS_X1 c6698(
.D(net6132),
.SE(net7128),
.SI(net4201),
.SN(net5181),
.CK(clk),
.Q(net7139),
.QN(net7138)
);

XNOR2_X2 c6699(
.A(net7121),
.B(net7139),
.ZN(net7140)
);

AND2_X4 c6700(
.A1(net7133),
.A2(net10859),
.ZN(net7141)
);

AND3_X1 c6701(
.A1(net7125),
.A2(net7082),
.A3(net10829),
.ZN(net7142)
);

AND2_X1 c6702(
.A1(net6182),
.A2(net7123),
.ZN(net7143)
);

NAND2_X1 c6703(
.A1(net7097),
.A2(net6098),
.ZN(net7144)
);

NAND3_X1 c6704(
.A1(net7015),
.A2(net7140),
.A3(net7122),
.ZN(net7145)
);

NAND2_X2 c6705(
.A1(net6124),
.A2(net7117),
.ZN(net7146)
);

NAND2_X4 c6706(
.A1(net7138),
.A2(net10896),
.ZN(net7147)
);

AND2_X2 c6707(
.A1(net7146),
.A2(net4992),
.ZN(net7148)
);

XOR2_X1 c6708(
.A(net7147),
.B(net6168),
.Z(net7149)
);

NOR2_X1 c6709(
.A1(net7076),
.A2(net5209),
.ZN(net7150)
);

OR2_X2 c6710(
.A1(net5974),
.A2(net7144),
.ZN(net7151)
);

NOR4_X4 c6711(
.A1(net7115),
.A2(net7144),
.A3(net7123),
.A4(net6168),
.ZN(net7152)
);

NOR2_X4 c6712(
.A1(net7125),
.A2(net7076),
.ZN(net7153)
);

SDFF_X2 c6713(
.D(net7153),
.SE(net7107),
.SI(net7132),
.CK(clk),
.Q(net7155),
.QN(net7154)
);

NOR3_X4 c6714(
.A1(net6121),
.A2(net7096),
.A3(net11461),
.ZN(net7156)
);

NOR2_X2 c6715(
.A1(net4159),
.A2(net7123),
.ZN(net7157)
);

NOR3_X2 c6716(
.A1(net7133),
.A2(net7157),
.A3(net11461),
.ZN(net7158)
);

AND3_X4 c6717(
.A1(net7156),
.A2(net7124),
.A3(net10918),
.ZN(net7159)
);

XOR2_X2 c6718(
.A(net7085),
.B(net7073),
.Z(net7160)
);

XNOR2_X1 c6719(
.A(net5978),
.B(net7156),
.ZN(net7161)
);

NAND3_X2 c6720(
.A1(net7157),
.A2(net7142),
.A3(net7151),
.ZN(net7162)
);

AOI222_X4 c6721(
.A1(net7156),
.A2(net7130),
.B1(net7037),
.B2(net7123),
.C1(net5975),
.C2(net10735),
.ZN(net7163)
);

OR2_X4 c6722(
.A1(net7161),
.A2(net11014),
.ZN(net7164)
);

INV_X8 c6723(
.A(net7111),
.ZN(net7165)
);

INV_X16 c6724(
.A(net7164),
.ZN(net7166)
);

OR2_X1 c6725(
.A1(net7100),
.A2(net5279),
.ZN(net7167)
);

NOR4_X2 c6726(
.A1(net7042),
.A2(net7074),
.A3(net5279),
.A4(net6262),
.ZN(net7168)
);

XNOR2_X2 c6727(
.A(net7151),
.B(net6273),
.ZN(net7169)
);

INV_X32 c6728(
.A(net7064),
.ZN(net7170)
);

SDFFS_X2 c6729(
.D(net6071),
.SE(net5222),
.SI(net7169),
.SN(net11405),
.CK(clk),
.Q(net7172),
.QN(net7171)
);

DFFRS_X1 c6730(
.D(net6256),
.RN(net7140),
.SN(net6195),
.CK(clk),
.Q(net7174),
.QN(net7173)
);

AND2_X4 c6731(
.A1(net6221),
.A2(net7042),
.ZN(net7175)
);

AND2_X1 c6732(
.A1(net7056),
.A2(net6273),
.ZN(net7176)
);

INV_X4 c6733(
.A(net5243),
.ZN(net7177)
);

INV_X1 c6734(
.A(net10247),
.ZN(net7178)
);

NAND2_X1 c6735(
.A1(net5935),
.A2(net7169),
.ZN(net7179)
);

INV_X2 c6736(
.A(net7139),
.ZN(net7180)
);

NAND2_X2 c6737(
.A1(net6251),
.A2(net5180),
.ZN(net7181)
);

INV_X8 c6738(
.A(net7140),
.ZN(net7182)
);

INV_X16 c6739(
.A(net9665),
.ZN(net7183)
);

INV_X32 c6740(
.A(net10500),
.ZN(net7184)
);

NAND2_X4 c6741(
.A1(net7177),
.A2(net7095),
.ZN(net7185)
);

AND2_X2 c6742(
.A1(net5279),
.A2(net6257),
.ZN(net7186)
);

DFFR_X2 c6743(
.D(net7128),
.RN(net7169),
.CK(clk),
.Q(net7188),
.QN(net7187)
);

OR3_X1 c6744(
.A1(net7136),
.A2(net7172),
.A3(net5101),
.ZN(net7189)
);

XOR2_X1 c6745(
.A(net6987),
.B(net11543),
.Z(net7190)
);

INV_X4 c6746(
.A(net11435),
.ZN(net7191)
);

INV_X1 c6747(
.A(net10020),
.ZN(net7192)
);

NOR2_X1 c6748(
.A1(net6263),
.A2(net11209),
.ZN(net7193)
);

OR2_X2 c6749(
.A1(net6248),
.A2(net7172),
.ZN(net7194)
);

MUX2_X1 c6750(
.A(net7099),
.B(net6208),
.S(net7173),
.Z(net7195)
);

INV_X2 c6751(
.A(net7144),
.ZN(net7196)
);

NOR2_X4 c6752(
.A1(net7180),
.A2(net11505),
.ZN(net7197)
);

INV_X8 c6753(
.A(net10390),
.ZN(net7198)
);

INV_X16 c6754(
.A(net10447),
.ZN(net7199)
);

INV_X32 c6755(
.A(net7188),
.ZN(net7200)
);

NOR2_X2 c6756(
.A1(net7185),
.A2(net6221),
.ZN(net7201)
);

INV_X4 c6757(
.A(net6125),
.ZN(net7202)
);

XOR2_X2 c6758(
.A(net7096),
.B(net7196),
.Z(net7203)
);

INV_X1 c6759(
.A(net11351),
.ZN(net7204)
);

XNOR2_X1 c6760(
.A(net7202),
.B(net7195),
.ZN(net7205)
);

INV_X2 c6761(
.A(net7198),
.ZN(net7206)
);

OR2_X4 c6762(
.A1(net4250),
.A2(net1130),
.ZN(net7207)
);

INV_X8 c6763(
.A(net6000),
.ZN(net7208)
);

INV_X16 c6764(
.A(net7207),
.ZN(net7209)
);

INV_X32 c6765(
.A(net4282),
.ZN(net7210)
);

INV_X4 c6766(
.A(net7152),
.ZN(net7211)
);

OR2_X1 c6767(
.A1(net7193),
.A2(net7198),
.ZN(net7212)
);

DFFRS_X2 c6768(
.D(net7200),
.RN(net7196),
.SN(net7169),
.CK(clk),
.Q(net7214),
.QN(net7213)
);

XNOR2_X2 c6769(
.A(net6253),
.B(net3912),
.ZN(net7215)
);

AND2_X4 c6770(
.A1(net7199),
.A2(net6187),
.ZN(net7216)
);

AND2_X1 c6771(
.A1(net7205),
.A2(net7083),
.ZN(net7217)
);

NAND2_X1 c6772(
.A1(net6262),
.A2(net7127),
.ZN(net7218)
);

NAND2_X2 c6773(
.A1(net7215),
.A2(net6125),
.ZN(net7219)
);

OAI21_X4 c6774(
.A(net7191),
.B1(net6270),
.B2(net7063),
.ZN(net7220)
);

INV_X1 c6775(
.A(net5181),
.ZN(net7221)
);

INV_X2 c6776(
.A(net9665),
.ZN(net7222)
);

MUX2_X2 c6777(
.A(net7204),
.B(net7167),
.S(net7182),
.Z(net7223)
);

NAND3_X4 c6778(
.A1(net7216),
.A2(net7215),
.A3(net7151),
.ZN(net7224)
);

NAND2_X4 c6779(
.A1(net7221),
.A2(net7080),
.ZN(net7225)
);

AND2_X2 c6780(
.A1(net7056),
.A2(net11021),
.ZN(net7226)
);

XOR2_X1 c6781(
.A(net7165),
.B(net10670),
.Z(net7227)
);

NOR2_X1 c6782(
.A1(net6223),
.A2(net7221),
.ZN(net7228)
);

INV_X8 c6783(
.A(net9944),
.ZN(net7229)
);

INV_X16 c6784(
.A(net11333),
.ZN(net7230)
);

INV_X32 c6785(
.A(net7194),
.ZN(net7231)
);

OR2_X2 c6786(
.A1(net7209),
.A2(net5224),
.ZN(net7232)
);

SDFF_X1 c6787(
.D(net7201),
.SE(net7187),
.SI(net7167),
.CK(clk),
.Q(net7234),
.QN(net7233)
);

INV_X4 c6788(
.A(net10043),
.ZN(net7235)
);

INV_X1 c6789(
.A(net9895),
.ZN(net7236)
);

OR3_X4 c6790(
.A1(net7203),
.A2(net7226),
.A3(net5935),
.ZN(net7237)
);

NOR2_X4 c6791(
.A1(net7221),
.A2(net10750),
.ZN(net7238)
);

AND3_X2 c6792(
.A1(net7210),
.A2(net7217),
.A3(net5200),
.ZN(net7239)
);

NOR2_X2 c6793(
.A1(net7230),
.A2(net7165),
.ZN(net7240)
);

INV_X2 c6794(
.A(net10475),
.ZN(net7241)
);

SDFFRS_X1 c6795(
.D(net7224),
.RN(net7240),
.SE(net7230),
.SI(net7172),
.SN(net7169),
.CK(clk),
.Q(net7243),
.QN(net7242)
);

INV_X8 c6796(
.A(net9803),
.ZN(net7244)
);

OAI33_X1 c6797(
.A1(net7240),
.A2(net7239),
.A3(net7218),
.B1(net5924),
.B2(net5234),
.B3(net7169),
.ZN(net7245)
);

AOI211_X4 c6798(
.A(net6211),
.B(net7202),
.C1(net7221),
.C2(net11558),
.ZN(net7246)
);

XOR2_X2 c6799(
.A(net6237),
.B(net7228),
.Z(net7247)
);

NOR3_X1 c6800(
.A1(net7192),
.A2(net7244),
.A3(net7240),
.ZN(net7248)
);

XNOR2_X1 c6801(
.A(net7231),
.B(net7234),
.ZN(net7249)
);

OR3_X2 c6802(
.A1(net6271),
.A2(net7249),
.A3(net7247),
.ZN(net7250)
);

OAI21_X2 c6803(
.A(net7248),
.B1(net7242),
.B2(net7244),
.ZN(net7251)
);

OAI21_X1 c6804(
.A(net7212),
.B1(net7248),
.B2(net7214),
.ZN(net7252)
);

AOI222_X2 c6805(
.A1(net7236),
.A2(net7208),
.B1(net7252),
.B2(net7251),
.C1(net7213),
.C2(net7124),
.ZN(net7253)
);

INV_X16 c6806(
.A(net6021),
.ZN(net7254)
);

OR2_X4 c6807(
.A1(net6329),
.A2(net7235),
.ZN(net7255)
);

INV_X32 c6808(
.A(net4328),
.ZN(net7256)
);

INV_X4 c6809(
.A(net10207),
.ZN(net7257)
);

INV_X1 c6810(
.A(net9716),
.ZN(net7258)
);

OR2_X1 c6811(
.A1(net4369),
.A2(net7173),
.ZN(net7259)
);

XNOR2_X2 c6812(
.A(net6258),
.B(net6021),
.ZN(net7260)
);

INV_X2 c6813(
.A(net6347),
.ZN(net7261)
);

INV_X8 c6814(
.A(net6100),
.ZN(net7262)
);

INV_X16 c6815(
.A(net7261),
.ZN(net7263)
);

INV_X32 c6816(
.A(net6113),
.ZN(net7264)
);

AND2_X4 c6817(
.A1(net7262),
.A2(net6318),
.ZN(net7265)
);

INV_X4 c6818(
.A(net9715),
.ZN(net7266)
);

AOI21_X2 c6819(
.A(net7258),
.B1(net6290),
.B2(net6319),
.ZN(net7267)
);

INV_X1 c6820(
.A(net11383),
.ZN(net7268)
);

INV_X2 c6821(
.A(net7263),
.ZN(net7269)
);

INV_X8 c6822(
.A(net5313),
.ZN(net7270)
);

INV_X16 c6823(
.A(net7265),
.ZN(net7271)
);

INV_X32 c6824(
.A(net7234),
.ZN(net7272)
);

AOI21_X1 c6825(
.A(net3155),
.B1(net7259),
.B2(net6297),
.ZN(net7273)
);

INV_X4 c6826(
.A(net7181),
.ZN(net7274)
);

INV_X1 c6827(
.A(net7243),
.ZN(net7275)
);

AND2_X1 c6828(
.A1(net7256),
.A2(net7247),
.ZN(net7276)
);

INV_X2 c6829(
.A(net4401),
.ZN(net7277)
);

AOI21_X4 c6830(
.A(net7222),
.B1(net7168),
.B2(net7238),
.ZN(net7278)
);

INV_X8 c6831(
.A(net10430),
.ZN(net7279)
);

NAND2_X1 c6832(
.A1(net7268),
.A2(net6354),
.ZN(net7280)
);

INV_X16 c6833(
.A(net6346),
.ZN(net7281)
);

NAND2_X2 c6834(
.A1(net7244),
.A2(net7258),
.ZN(net7282)
);

NAND2_X4 c6835(
.A1(net7270),
.A2(net6346),
.ZN(net7283)
);

INV_X32 c6836(
.A(net7275),
.ZN(net7284)
);

AND2_X2 c6837(
.A1(net7195),
.A2(net7038),
.ZN(net7285)
);

INV_X4 c6838(
.A(net4085),
.ZN(net7286)
);

INV_X1 c6839(
.A(net6318),
.ZN(net7287)
);

INV_X2 c6840(
.A(net6312),
.ZN(net7288)
);

XOR2_X1 c6841(
.A(net7257),
.B(net11305),
.Z(net7289)
);

NOR2_X1 c6842(
.A1(net5356),
.A2(net7233),
.ZN(net7290)
);

INV_X8 c6843(
.A(net7255),
.ZN(net7291)
);

INV_X16 c6844(
.A(net3432),
.ZN(net7292)
);

OR2_X2 c6845(
.A1(net7292),
.A2(net7244),
.ZN(net7293)
);

INV_X32 c6846(
.A(net9955),
.ZN(net7294)
);

NOR2_X4 c6847(
.A1(net7218),
.A2(net6264),
.ZN(net7295)
);

NOR2_X2 c6848(
.A1(net7266),
.A2(net7265),
.ZN(net7296)
);

OAI221_X1 c6849(
.A(net5200),
.B1(net7243),
.B2(net7233),
.C1(net7171),
.C2(net7213),
.ZN(net7297)
);

XOR2_X2 c6850(
.A(net7168),
.B(net7214),
.Z(net7298)
);

SDFF_X2 c6851(
.D(net4364),
.SE(net6259),
.SI(net7274),
.CK(clk),
.Q(net7300),
.QN(net7299)
);

XNOR2_X1 c6852(
.A(net7276),
.B(net7265),
.ZN(net7301)
);

DFFRS_X1 c6853(
.D(net7174),
.RN(net6264),
.SN(net7273),
.CK(clk),
.Q(net7303),
.QN(net7302)
);

OR2_X4 c6854(
.A1(net7274),
.A2(net7288),
.ZN(net7304)
);

AND3_X1 c6855(
.A1(net7259),
.A2(net7169),
.A3(net7266),
.ZN(net7305)
);

INV_X4 c6856(
.A(net10671),
.ZN(net7306)
);

NAND3_X1 c6857(
.A1(net7297),
.A2(net6333),
.A3(net7277),
.ZN(net7307)
);

INV_X1 c6858(
.A(net7271),
.ZN(net7308)
);

OR2_X1 c6859(
.A1(net7171),
.A2(net11343),
.ZN(net7309)
);

XNOR2_X2 c6860(
.A(net5344),
.B(net7247),
.ZN(net7310)
);

AND2_X4 c6861(
.A1(net7080),
.A2(net6302),
.ZN(net7311)
);

AND2_X1 c6862(
.A1(net7294),
.A2(net4084),
.ZN(net7312)
);

OAI221_X4 c6863(
.A(net7272),
.B1(net5356),
.B2(net7309),
.C1(net7252),
.C2(net7213),
.ZN(net7313)
);

NOR3_X4 c6864(
.A1(net7132),
.A2(net7311),
.A3(net7287),
.ZN(net7314)
);

INV_X2 c6865(
.A(net9872),
.ZN(net7315)
);

NOR3_X2 c6866(
.A1(net7289),
.A2(net7218),
.A3(net6263),
.ZN(net7316)
);

AND3_X4 c6867(
.A1(net7311),
.A2(net7288),
.A3(net5313),
.ZN(net7317)
);

NAND2_X1 c6868(
.A1(net7306),
.A2(net11240),
.ZN(net7318)
);

NAND2_X2 c6869(
.A1(net7293),
.A2(net7074),
.ZN(net7319)
);

NAND2_X4 c6870(
.A1(net4399),
.A2(net6347),
.ZN(net7320)
);

AND2_X2 c6871(
.A1(net7311),
.A2(net10639),
.ZN(net7321)
);

XOR2_X1 c6872(
.A(net7285),
.B(net7319),
.Z(net7322)
);

NOR2_X1 c6873(
.A1(net7313),
.A2(net11438),
.ZN(net7323)
);

OR2_X2 c6874(
.A1(net7301),
.A2(net7296),
.ZN(net7324)
);

INV_X8 c6875(
.A(net11216),
.ZN(net7325)
);

NAND3_X2 c6876(
.A1(net7325),
.A2(net7124),
.A3(net7112),
.ZN(net7326)
);

OR3_X1 c6877(
.A1(net6356),
.A2(net7326),
.A3(net7263),
.ZN(net7327)
);

NOR2_X4 c6878(
.A1(net7318),
.A2(net7174),
.ZN(net7328)
);

INV_X16 c6879(
.A(net11087),
.ZN(net7329)
);

MUX2_X1 c6880(
.A(net7284),
.B(net7324),
.S(net7329),
.Z(net7330)
);

OAI21_X4 c6881(
.A(net6319),
.B1(net7326),
.B2(net7312),
.ZN(net7331)
);

NOR4_X1 c6882(
.A1(net7254),
.A2(net7321),
.A3(net7326),
.A4(net7312),
.ZN(net7332)
);

NOR2_X2 c6883(
.A1(net7316),
.A2(net7311),
.ZN(net7333)
);

MUX2_X2 c6884(
.A(net7333),
.B(net7320),
.S(net7331),
.Z(net7334)
);

AOI211_X2 c6885(
.A(net7039),
.B(net7277),
.C1(net7331),
.C2(net7311),
.ZN(net7335)
);

AOI22_X1 c6886(
.A1(net7328),
.A2(net7326),
.B1(net7331),
.B2(net7288),
.ZN(net7336)
);

OAI221_X2 c6887(
.A(net7335),
.B1(net7197),
.B2(net7326),
.C1(net6365),
.C2(net7296),
.ZN(net7337)
);

AOI221_X4 c6888(
.A(net7334),
.B1(net7112),
.B2(net7299),
.C1(net10719),
.C2(net11433),
.ZN(net7338)
);

XOR2_X2 c6889(
.A(net6177),
.B(net7252),
.Z(net7339)
);

XNOR2_X1 c6890(
.A(net5113),
.B(net6177),
.ZN(net7340)
);

OR2_X4 c6891(
.A1(net5399),
.A2(net5467),
.ZN(net7341)
);

OR2_X1 c6892(
.A1(net6431),
.A2(net2380),
.ZN(net7342)
);

INV_X32 c6893(
.A(net6071),
.ZN(net7343)
);

XNOR2_X2 c6894(
.A(net7279),
.B(net6386),
.ZN(net7344)
);

INV_X4 c6895(
.A(net6440),
.ZN(net7345)
);

AND2_X4 c6896(
.A1(net3520),
.A2(net7296),
.ZN(net7346)
);

AND2_X1 c6897(
.A1(net7247),
.A2(net7196),
.ZN(net7347)
);

NAND2_X1 c6898(
.A1(net6313),
.A2(net6354),
.ZN(net7348)
);

NAND2_X2 c6899(
.A1(net7346),
.A2(net7277),
.ZN(net7349)
);

NAND2_X4 c6900(
.A1(net6448),
.A2(net6440),
.ZN(net7350)
);

AND2_X2 c6901(
.A1(net6263),
.A2(net6306),
.ZN(net7351)
);

XOR2_X1 c6902(
.A(net7340),
.B(net6439),
.Z(net7352)
);

NOR2_X1 c6903(
.A1(net7317),
.A2(net7112),
.ZN(net7353)
);

NAND3_X4 c6904(
.A1(net7344),
.A2(net7334),
.A3(net6450),
.ZN(net7354)
);

OR2_X2 c6905(
.A1(net7310),
.A2(net7352),
.ZN(net7355)
);

INV_X1 c6906(
.A(net7347),
.ZN(net7356)
);

INV_X2 c6907(
.A(net10373),
.ZN(net7357)
);

NOR2_X4 c6908(
.A1(net7196),
.A2(net7344),
.ZN(net7358)
);

NOR2_X2 c6909(
.A1(net7112),
.A2(net7356),
.ZN(net7359)
);

INV_X8 c6910(
.A(net9781),
.ZN(net7360)
);

XOR2_X2 c6911(
.A(net7352),
.B(net7303),
.Z(net7361)
);

INV_X16 c6912(
.A(net11401),
.ZN(net7362)
);

XNOR2_X1 c6913(
.A(net7135),
.B(net11306),
.ZN(net7363)
);

OR2_X4 c6914(
.A1(net5468),
.A2(net6257),
.ZN(net7364)
);

OR2_X1 c6915(
.A1(net6386),
.A2(net6448),
.ZN(net7365)
);

OR3_X4 c6916(
.A1(net7238),
.A2(net6451),
.A3(net7352),
.ZN(net7366)
);

INV_X32 c6917(
.A(net10087),
.ZN(net7367)
);

XNOR2_X2 c6918(
.A(net7169),
.B(net6440),
.ZN(net7368)
);

AND2_X4 c6919(
.A1(net7343),
.A2(net6365),
.ZN(net7369)
);

AND2_X1 c6920(
.A1(net6383),
.A2(net7352),
.ZN(net7370)
);

INV_X4 c6921(
.A(net9926),
.ZN(net7371)
);

NAND2_X1 c6922(
.A1(net7362),
.A2(net10582),
.ZN(net7372)
);

NAND2_X2 c6923(
.A1(net6852),
.A2(net7362),
.ZN(net7373)
);

INV_X1 c6924(
.A(net10279),
.ZN(net7374)
);

NAND2_X4 c6925(
.A1(net6883),
.A2(net7358),
.ZN(net7375)
);

SDFFR_X1 c6926(
.D(net7361),
.RN(net7371),
.SE(net6369),
.SI(net6354),
.CK(clk),
.Q(net7377),
.QN(net7376)
);

AND2_X2 c6927(
.A1(net7365),
.A2(net6442),
.ZN(net7378)
);

XOR2_X1 c6928(
.A(net7374),
.B(net6440),
.Z(net7379)
);

AND3_X2 c6929(
.A1(net6425),
.A2(net7351),
.A3(net7372),
.ZN(net7380)
);

NOR2_X1 c6930(
.A1(net7349),
.A2(net7332),
.ZN(net7381)
);

OR2_X2 c6931(
.A1(net6396),
.A2(net7371),
.ZN(net7382)
);

NOR2_X4 c6932(
.A1(net6442),
.A2(net7287),
.ZN(net7383)
);

NOR2_X2 c6933(
.A1(net7367),
.A2(net7371),
.ZN(net7384)
);

INV_X2 c6934(
.A(net9950),
.ZN(net7385)
);

XOR2_X2 c6935(
.A(net7358),
.B(net7385),
.Z(net7386)
);

INV_X8 c6936(
.A(net11458),
.ZN(net7387)
);

XNOR2_X1 c6937(
.A(net7383),
.B(net7269),
.ZN(net7388)
);

OR2_X4 c6938(
.A1(net7303),
.A2(net7312),
.ZN(net7389)
);

INV_X16 c6939(
.A(net10438),
.ZN(net7390)
);

OAI222_X1 c6940(
.A1(net7384),
.A2(net7390),
.B1(net6407),
.B2(net6263),
.C1(net7356),
.C2(net6050),
.ZN(net7391)
);

OR2_X1 c6941(
.A1(net7387),
.A2(net7286),
.ZN(net7392)
);

INV_X32 c6942(
.A(net9983),
.ZN(net7393)
);

NOR3_X1 c6943(
.A1(net7375),
.A2(net7377),
.A3(net11444),
.ZN(net7394)
);

XNOR2_X2 c6944(
.A(net7394),
.B(net7390),
.ZN(net7395)
);

AND2_X4 c6945(
.A1(net7389),
.A2(net11305),
.ZN(net7396)
);

AND2_X1 c6946(
.A1(net5463),
.A2(net7352),
.ZN(net7397)
);

NAND2_X1 c6947(
.A1(net7286),
.A2(net7344),
.ZN(net7398)
);

INV_X4 c6948(
.A(net11092),
.ZN(net7399)
);

NAND2_X2 c6949(
.A1(net7373),
.A2(net7351),
.ZN(net7400)
);

NAND2_X4 c6950(
.A1(net7396),
.A2(net6177),
.ZN(net7401)
);

OR3_X2 c6951(
.A1(net7386),
.A2(net7389),
.A3(net7401),
.ZN(net7402)
);

DFFRS_X2 c6952(
.D(net5444),
.RN(net7400),
.SN(net7280),
.CK(clk),
.Q(net7404),
.QN(net7403)
);

INV_X1 c6953(
.A(net9780),
.ZN(net7405)
);

AND4_X4 c6954(
.A1(net7362),
.A2(net6302),
.A3(net6442),
.A4(net7363),
.ZN(net7406)
);

AOI221_X2 c6955(
.A(net7384),
.B1(net7400),
.B2(net7356),
.C1(net7405),
.C2(net11444),
.ZN(net7407)
);

AND2_X2 c6956(
.A1(net7380),
.A2(net7403),
.ZN(net7408)
);

XOR2_X1 c6957(
.A(net7371),
.B(net7402),
.Z(net7409)
);

OAI21_X2 c6958(
.A(net7304),
.B1(net6364),
.B2(net7407),
.ZN(net7410)
);

SDFF_X1 c6959(
.D(net7364),
.SE(net7363),
.SI(net7394),
.CK(clk),
.Q(net7412),
.QN(net7411)
);

SDFF_X2 c6960(
.D(net7407),
.SE(net7411),
.SI(net5351),
.CK(clk),
.Q(net7414),
.QN(net7413)
);

OAI222_X4 c6961(
.A1(net7408),
.A2(net7398),
.B1(net7407),
.B2(net5351),
.C1(net7413),
.C2(net7169),
.ZN(net7415)
);

OAI21_X1 c6962(
.A(net5180),
.B1(net7401),
.B2(net11481),
.ZN(net7416)
);

AOI21_X2 c6963(
.A(net5408),
.B1(net7385),
.B2(net11480),
.ZN(net7417)
);

AOI21_X1 c6964(
.A(net7417),
.B1(net7399),
.B2(net7406),
.ZN(net7418)
);

AOI21_X4 c6965(
.A(net7404),
.B1(net7407),
.B2(net7299),
.ZN(net7419)
);

AND3_X1 c6966(
.A1(net7381),
.A2(net7334),
.A3(net7405),
.ZN(net7420)
);

NAND3_X1 c6967(
.A1(net7375),
.A2(net7360),
.A3(net11480),
.ZN(net7421)
);

NOR3_X4 c6968(
.A1(net7406),
.A2(net7412),
.A3(net7421),
.ZN(net7422)
);

NAND4_X1 c6969(
.A1(net7355),
.A2(net7401),
.A3(net7356),
.A4(net11090),
.ZN(net7423)
);

OAI222_X2 c6970(
.A1(net4413),
.A2(net7412),
.B1(net5224),
.B2(net7344),
.C1(net7413),
.C2(net7376),
.ZN(net7424)
);

OR4_X1 c6971(
.A1(net7385),
.A2(net7391),
.A3(net5393),
.A4(net6397),
.ZN(net7425)
);

DFFRS_X1 c6972(
.D(net4583),
.RN(net6365),
.SN(net7013),
.CK(clk),
.Q(net7427),
.QN(net7426)
);

NOR3_X2 c6973(
.A1(net7378),
.A2(net3586),
.A3(net7189),
.ZN(net7428)
);

NOR2_X1 c6974(
.A1(net6468),
.A2(net5179),
.ZN(net7429)
);

INV_X2 c6975(
.A(net6520),
.ZN(net7430)
);

INV_X8 c6976(
.A(net7260),
.ZN(net7431)
);

INV_X16 c6977(
.A(net9702),
.ZN(net7432)
);

INV_X32 c6978(
.A(net9702),
.ZN(net7433)
);

INV_X4 c6979(
.A(net10215),
.ZN(net7434)
);

OR2_X2 c6980(
.A1(net3548),
.A2(net7269),
.ZN(net7435)
);

INV_X1 c6981(
.A(net7135),
.ZN(net7436)
);

NOR2_X4 c6982(
.A1(net7280),
.A2(net11415),
.ZN(net7437)
);

INV_X2 c6983(
.A(net11416),
.ZN(net7438)
);

DFFRS_X2 c6984(
.D(net6257),
.RN(net7246),
.SN(net6541),
.CK(clk),
.Q(net7440),
.QN(net7439)
);

INV_X8 c6985(
.A(net9938),
.ZN(net7441)
);

INV_X16 c6986(
.A(net9978),
.ZN(net7442)
);

SDFF_X1 c6987(
.D(net7246),
.SE(net6476),
.SI(net6050),
.CK(clk),
.Q(net7444),
.QN(net7443)
);

INV_X32 c6988(
.A(net10290),
.ZN(net7445)
);

INV_X4 c6989(
.A(net11333),
.ZN(net7446)
);

NOR2_X2 c6990(
.A1(net6378),
.A2(net7434),
.ZN(net7447)
);

XOR2_X2 c6991(
.A(net6480),
.B(net7443),
.Z(net7448)
);

INV_X1 c6992(
.A(net7315),
.ZN(net7449)
);

INV_X2 c6993(
.A(net11442),
.ZN(net7450)
);

INV_X8 c6994(
.A(net6499),
.ZN(net7451)
);

XNOR2_X1 c6995(
.A(net7388),
.B(net6305),
.ZN(net7452)
);

OR2_X4 c6996(
.A1(net6410),
.A2(net7433),
.ZN(net7453)
);

INV_X16 c6997(
.A(net7392),
.ZN(net7454)
);

OR2_X1 c6998(
.A1(net7453),
.A2(net5552),
.ZN(net7455)
);

XNOR2_X2 c6999(
.A(net5388),
.B(net7447),
.ZN(net7456)
);

AND2_X4 c7000(
.A1(net7438),
.A2(net6494),
.ZN(net7457)
);

AND3_X4 c7001(
.A1(net6535),
.A2(net7457),
.A3(net7219),
.ZN(net7458)
);

AND2_X1 c7002(
.A1(net7283),
.A2(net7433),
.ZN(net7459)
);

NAND2_X1 c7003(
.A1(net7456),
.A2(net6519),
.ZN(net7460)
);

NAND2_X2 c7004(
.A1(net6409),
.A2(net7452),
.ZN(net7461)
);

INV_X32 c7005(
.A(net9819),
.ZN(net7462)
);

INV_X4 c7006(
.A(net10103),
.ZN(net7463)
);

NAND2_X4 c7007(
.A1(net6523),
.A2(net7442),
.ZN(net7464)
);

AND2_X2 c7008(
.A1(net7461),
.A2(net7443),
.ZN(net7465)
);

NAND3_X2 c7009(
.A1(net7462),
.A2(net7375),
.A3(net7464),
.ZN(net7466)
);

INV_X1 c7010(
.A(net6435),
.ZN(net7467)
);

XOR2_X1 c7011(
.A(net7189),
.B(net7315),
.Z(net7468)
);

NOR2_X1 c7012(
.A1(net7353),
.A2(net7445),
.ZN(net7469)
);

OR2_X2 c7013(
.A1(net7463),
.A2(net6486),
.ZN(net7470)
);

DFFS_X1 c7014(
.D(net7313),
.SN(net7363),
.CK(clk),
.Q(net7472),
.QN(net7471)
);

NOR2_X4 c7015(
.A1(net7360),
.A2(net7439),
.ZN(net7473)
);

OR3_X1 c7016(
.A1(net7473),
.A2(net7458),
.A3(net5388),
.ZN(net7474)
);

MUX2_X1 c7017(
.A(net7446),
.B(net7474),
.S(net7448),
.Z(net7475)
);

INV_X2 c7018(
.A(net9964),
.ZN(net7476)
);

NOR2_X2 c7019(
.A1(net1562),
.A2(net6297),
.ZN(net7477)
);

OAI21_X4 c7020(
.A(net7472),
.B1(net7462),
.B2(net5388),
.ZN(net7478)
);

XOR2_X2 c7021(
.A(net7468),
.B(net6507),
.Z(net7479)
);

INV_X8 c7022(
.A(net9939),
.ZN(net7480)
);

XNOR2_X1 c7023(
.A(net7469),
.B(net6476),
.ZN(net7481)
);

DFFS_X2 c7024(
.D(net7345),
.SN(net7471),
.CK(clk),
.Q(net7483),
.QN(net7482)
);

MUX2_X2 c7025(
.A(net6515),
.B(net7477),
.S(net7479),
.Z(net7484)
);

OR2_X4 c7026(
.A1(net6435),
.A2(net11429),
.ZN(net7485)
);

OR2_X1 c7027(
.A1(net5180),
.A2(net4322),
.ZN(net7486)
);

XNOR2_X2 c7028(
.A(net4542),
.B(net7475),
.ZN(net7487)
);

SDFF_X2 c7029(
.D(net7485),
.SE(net7444),
.SI(net7451),
.CK(clk),
.Q(net7489),
.QN(net7488)
);

INV_X16 c7030(
.A(net11151),
.ZN(net7490)
);

AND2_X4 c7031(
.A1(net7490),
.A2(net7445),
.ZN(net7491)
);

INV_X32 c7032(
.A(net7433),
.ZN(net7492)
);

AOI222_X1 c7033(
.A1(net7474),
.A2(net7241),
.B1(net6435),
.B2(net7363),
.C1(net7413),
.C2(net7445),
.ZN(net7493)
);

AND2_X1 c7034(
.A1(net7491),
.A2(net7479),
.ZN(net7494)
);

NAND2_X1 c7035(
.A1(net6493),
.A2(net7474),
.ZN(net7495)
);

NAND3_X4 c7036(
.A1(net7470),
.A2(net7440),
.A3(net11415),
.ZN(net7496)
);

NAND2_X2 c7037(
.A1(net7478),
.A2(net6410),
.ZN(net7497)
);

OR3_X4 c7038(
.A1(net2605),
.A2(net6486),
.A3(net7440),
.ZN(net7498)
);

NAND2_X4 c7039(
.A1(net7497),
.A2(net6495),
.ZN(net7499)
);

AND2_X2 c7040(
.A1(net7480),
.A2(net7246),
.ZN(net7500)
);

AND3_X2 c7041(
.A1(net7389),
.A2(net5388),
.A3(net6480),
.ZN(net7501)
);

XOR2_X1 c7042(
.A(net7486),
.B(net7496),
.Z(net7502)
);

NOR2_X1 c7043(
.A1(net7500),
.A2(net7499),
.ZN(net7503)
);

OR2_X2 c7044(
.A1(net7241),
.A2(net5540),
.ZN(net7504)
);

NOR3_X1 c7045(
.A1(net3446),
.A2(net7356),
.A3(net7457),
.ZN(net7505)
);

NOR2_X4 c7046(
.A1(net7492),
.A2(net7497),
.ZN(net7506)
);

INV_X4 c7047(
.A(net10173),
.ZN(net7507)
);

NOR2_X2 c7048(
.A1(net7496),
.A2(net7486),
.ZN(net7508)
);

INV_X1 c7049(
.A(net10149),
.ZN(net7509)
);

INV_X2 c7050(
.A(net11430),
.ZN(net7510)
);

DFFRS_X1 c7051(
.D(net7502),
.RN(net7487),
.SN(net7477),
.CK(clk),
.Q(net7512),
.QN(net7511)
);

DFFRS_X2 c7052(
.D(net3586),
.RN(net7241),
.SN(net7451),
.CK(clk),
.Q(net7514),
.QN(net7513)
);

OR3_X2 c7053(
.A1(net7510),
.A2(net7507),
.A3(net7513),
.ZN(net7515)
);

OAI21_X2 c7054(
.A(net7515),
.B1(net7485),
.B2(net7511),
.ZN(net7516)
);

INV_X8 c7055(
.A(net10037),
.ZN(net7517)
);

XOR2_X2 c7056(
.A(net2589),
.B(net5616),
.Z(net7518)
);

XNOR2_X1 c7057(
.A(net7377),
.B(net4652),
.ZN(net7519)
);

INV_X16 c7058(
.A(net9660),
.ZN(net7520)
);

OR2_X4 c7059(
.A1(net3645),
.A2(net6469),
.ZN(net7521)
);

INV_X32 c7060(
.A(net9963),
.ZN(net7522)
);

INV_X4 c7061(
.A(net10031),
.ZN(net7523)
);

OAI22_X1 c7062(
.A1(net7518),
.A2(net7475),
.B1(net7197),
.B2(net5545),
.ZN(net7524)
);

OR2_X1 c7063(
.A1(net6591),
.A2(net6615),
.ZN(net7525)
);

SDFF_X1 c7064(
.D(net5627),
.SE(net6591),
.SI(net7432),
.CK(clk),
.Q(net7527),
.QN(net7526)
);

XNOR2_X2 c7065(
.A(net6609),
.B(net7377),
.ZN(net7528)
);

AND2_X4 c7066(
.A1(net7503),
.A2(net5640),
.ZN(net7529)
);

AND2_X1 c7067(
.A1(net7479),
.A2(net7426),
.ZN(net7530)
);

SDFF_X2 c7068(
.D(net4612),
.SE(net7519),
.SI(net6548),
.CK(clk),
.Q(net7532),
.QN(net7531)
);

INV_X1 c7069(
.A(net10026),
.ZN(net7533)
);

INV_X2 c7070(
.A(net11469),
.ZN(net7534)
);

NAND2_X1 c7071(
.A1(net1637),
.A2(net7531),
.ZN(net7535)
);

NAND2_X2 c7072(
.A1(net4652),
.A2(net6397),
.ZN(net7536)
);

INV_X8 c7073(
.A(net11381),
.ZN(net7537)
);

NAND2_X4 c7074(
.A1(net6590),
.A2(net7460),
.ZN(net7538)
);

AND2_X2 c7075(
.A1(net7464),
.A2(net7267),
.ZN(net7539)
);

SDFFRS_X2 c7076(
.D(net6593),
.RN(net4542),
.SE(net6525),
.SI(net6212),
.SN(net3627),
.CK(clk),
.Q(net7541),
.QN(net7540)
);

SDFFR_X2 c7077(
.D(net7534),
.RN(net6559),
.SE(net5627),
.SI(net7535),
.CK(clk),
.Q(net7543),
.QN(net7542)
);

XOR2_X1 c7078(
.A(net7450),
.B(net7455),
.Z(net7544)
);

OAI21_X1 c7079(
.A(net7522),
.B1(net7526),
.B2(net7455),
.ZN(net7545)
);

INV_X16 c7080(
.A(net9965),
.ZN(net7546)
);

NOR2_X1 c7081(
.A1(net638),
.A2(net7464),
.ZN(net7547)
);

OR2_X2 c7082(
.A1(net6567),
.A2(net7377),
.ZN(net7548)
);

NOR2_X4 c7083(
.A1(net5522),
.A2(net7470),
.ZN(net7549)
);

NOR2_X2 c7084(
.A1(net7401),
.A2(net7267),
.ZN(net7550)
);

INV_X32 c7085(
.A(net10160),
.ZN(net7551)
);

XOR2_X2 c7086(
.A(net7267),
.B(net7401),
.Z(net7552)
);

AOI21_X2 c7087(
.A(net5641),
.B1(net6548),
.B2(net7533),
.ZN(net7553)
);

AND4_X2 c7088(
.A1(net6587),
.A2(net1732),
.A3(net7540),
.A4(net7535),
.ZN(net7554)
);

INV_X4 c7089(
.A(net10489),
.ZN(net7555)
);

AOI222_X4 c7090(
.A1(net5553),
.A2(net7543),
.B1(net6567),
.B2(net6611),
.C1(net7546),
.C2(net6609),
.ZN(net7556)
);

AOI21_X1 c7091(
.A(net7529),
.B1(net5522),
.B2(net7522),
.ZN(net7557)
);

XNOR2_X1 c7092(
.A(net7552),
.B(net7414),
.ZN(net7558)
);

OR2_X4 c7093(
.A1(net7470),
.A2(net7518),
.ZN(net7559)
);

OR2_X1 c7094(
.A1(net6596),
.A2(net7542),
.ZN(net7560)
);

INV_X1 c7095(
.A(net10457),
.ZN(net7561)
);

XNOR2_X2 c7096(
.A(net7553),
.B(net7501),
.ZN(net7562)
);

AND2_X4 c7097(
.A1(net7454),
.A2(net6611),
.ZN(net7563)
);

INV_X2 c7098(
.A(net10161),
.ZN(net7564)
);

AND2_X1 c7099(
.A1(net7537),
.A2(net7553),
.ZN(net7565)
);

INV_X8 c7100(
.A(net11384),
.ZN(net7566)
);

DFFRS_X1 c7101(
.D(net6626),
.RN(net7550),
.SN(net7560),
.CK(clk),
.Q(net7568),
.QN(net7567)
);

NAND2_X1 c7102(
.A1(net5552),
.A2(net7550),
.ZN(net7569)
);

NAND2_X2 c7103(
.A1(net7548),
.A2(net7559),
.ZN(net7570)
);

NAND2_X4 c7104(
.A1(net7564),
.A2(net7569),
.ZN(net7571)
);

AND2_X2 c7105(
.A1(net7528),
.A2(net7570),
.ZN(net7572)
);

XOR2_X1 c7106(
.A(net6611),
.B(net7504),
.Z(net7573)
);

NOR2_X1 c7107(
.A1(net7572),
.A2(net7571),
.ZN(net7574)
);

AOI21_X4 c7108(
.A(net7567),
.B1(net6553),
.B2(net10956),
.ZN(net7575)
);

OR2_X2 c7109(
.A1(net7550),
.A2(net7565),
.ZN(net7576)
);

NOR2_X4 c7110(
.A1(net6547),
.A2(net7566),
.ZN(net7577)
);

NOR2_X2 c7111(
.A1(net7573),
.A2(net10572),
.ZN(net7578)
);

XOR2_X2 c7112(
.A(net7565),
.B(net7445),
.Z(net7579)
);

XNOR2_X1 c7113(
.A(net7570),
.B(net7568),
.ZN(net7580)
);

OR2_X4 c7114(
.A1(net7575),
.A2(net6611),
.ZN(net7581)
);

OR2_X1 c7115(
.A1(net7476),
.A2(net7545),
.ZN(net7582)
);

AND4_X1 c7116(
.A1(net7527),
.A2(net7577),
.A3(net4604),
.A4(net7413),
.ZN(net7583)
);

AND3_X1 c7117(
.A1(net7457),
.A2(net6486),
.A3(net7559),
.ZN(net7584)
);

XNOR2_X2 c7118(
.A(net711),
.B(net7421),
.ZN(net7585)
);

AND2_X4 c7119(
.A1(net7547),
.A2(net7566),
.ZN(net7586)
);

NAND3_X1 c7120(
.A1(net7585),
.A2(net7553),
.A3(net7581),
.ZN(net7587)
);

DFFRS_X2 c7121(
.D(net4534),
.RN(net7550),
.SN(net7587),
.CK(clk),
.Q(net7589),
.QN(net7588)
);

NOR3_X4 c7122(
.A1(net7576),
.A2(out25),
.A3(net7575),
.ZN(net7590)
);

AND2_X1 c7123(
.A1(net7375),
.A2(net4598),
.ZN(net7591)
);

NOR3_X2 c7124(
.A1(net7584),
.A2(net7589),
.A3(net7582),
.ZN(net7592)
);

NAND2_X1 c7125(
.A1(net7579),
.A2(net7566),
.ZN(net7593)
);

AND3_X4 c7126(
.A1(net7395),
.A2(net7580),
.A3(net7585),
.ZN(net7594)
);

NAND2_X2 c7127(
.A1(net7593),
.A2(net7592),
.ZN(net7595)
);

NAND3_X2 c7128(
.A1(net7273),
.A2(net7595),
.A3(net7585),
.ZN(net7596)
);

OR3_X1 c7129(
.A1(net7581),
.A2(net7572),
.A3(net7585),
.ZN(net7597)
);

MUX2_X1 c7130(
.A(net7431),
.B(net7518),
.S(net7506),
.Z(net7598)
);

SDFF_X1 c7131(
.D(net7594),
.SE(net7575),
.SI(net6533),
.CK(clk),
.Q(net7600),
.QN(net7599)
);

OAI21_X4 c7132(
.A(net7586),
.B1(net7529),
.B2(net7598),
.ZN(net7601)
);

AOI22_X4 c7133(
.A1(net7523),
.A2(net7535),
.B1(net5522),
.B2(net4523),
.ZN(net7602)
);

SDFF_X2 c7134(
.D(net7598),
.SE(net7593),
.SI(net7599),
.CK(clk),
.Q(net7604),
.QN(net7603)
);

OAI33_X1 c7135(
.A1(net7573),
.A2(net7600),
.A3(net7575),
.B1(net6611),
.B2(net7577),
.B3(net7578),
.ZN(net7605)
);

MUX2_X2 c7136(
.A(net10978),
.B(net11373),
.S(net11563),
.Z(net7606)
);

INV_X16 c7137(
.A(net9659),
.ZN(net7607)
);

NAND2_X4 c7138(
.A1(net7341),
.A2(net6694),
.ZN(net7608)
);

AND2_X2 c7139(
.A1(net7525),
.A2(net6569),
.ZN(net7609)
);

XOR2_X1 c7140(
.A(net6649),
.B(net7269),
.Z(net7610)
);

NOR2_X1 c7141(
.A1(net7604),
.A2(net3749),
.ZN(net7611)
);

OR2_X2 c7142(
.A1(net2777),
.A2(net7583),
.ZN(net7612)
);

NOR2_X4 c7143(
.A1(net7520),
.A2(net6711),
.ZN(net7613)
);

INV_X32 c7144(
.A(net9836),
.ZN(net7614)
);

NOR2_X2 c7145(
.A1(net4322),
.A2(net6694),
.ZN(net7615)
);

XOR2_X2 c7146(
.A(net6688),
.B(net6668),
.Z(net7616)
);

INV_X4 c7147(
.A(net9670),
.ZN(net7617)
);

XNOR2_X1 c7148(
.A(net6569),
.B(net7546),
.ZN(net7618)
);

OR2_X4 c7149(
.A1(net7538),
.A2(net7591),
.ZN(net7619)
);

OR2_X1 c7150(
.A1(net6696),
.A2(net7615),
.ZN(net7620)
);

XNOR2_X2 c7151(
.A(net7583),
.B(net7603),
.ZN(net7621)
);

AND2_X4 c7152(
.A1(net7610),
.A2(net7614),
.ZN(net7622)
);

NAND3_X4 c7153(
.A1(net4729),
.A2(net6050),
.A3(net11563),
.ZN(net7623)
);

OR3_X4 c7154(
.A1(net7615),
.A2(net7448),
.A3(net3742),
.ZN(net7624)
);

AND2_X1 c7155(
.A1(net7506),
.A2(net4742),
.ZN(net7625)
);

AOI221_X1 c7156(
.A(net2751),
.B1(net5702),
.B2(net2713),
.C1(net6689),
.C2(net3691),
.ZN(net7626)
);

NAND2_X1 c7157(
.A1(net6654),
.A2(net6548),
.ZN(net7627)
);

NAND2_X2 c7158(
.A1(net5689),
.A2(net720),
.ZN(net7628)
);

NAND2_X4 c7159(
.A1(net4742),
.A2(net7615),
.ZN(net7629)
);

AND2_X2 c7160(
.A1(net6698),
.A2(net6569),
.ZN(net7630)
);

INV_X1 c7161(
.A(net9669),
.ZN(net7631)
);

XOR2_X1 c7162(
.A(net4524),
.B(net4704),
.Z(net7632)
);

NOR2_X1 c7163(
.A1(net6660),
.A2(net7609),
.ZN(net7633)
);

OR2_X2 c7164(
.A1(net7614),
.A2(net7618),
.ZN(net7634)
);

NOR2_X4 c7165(
.A1(net7620),
.A2(net7615),
.ZN(net7635)
);

NOR2_X2 c7166(
.A1(net7427),
.A2(net7609),
.ZN(net7636)
);

XOR2_X2 c7167(
.A(net7532),
.B(net5689),
.Z(net7637)
);

INV_X2 c7168(
.A(net9979),
.ZN(net7638)
);

XNOR2_X1 c7169(
.A(net7609),
.B(net3742),
.ZN(net7639)
);

AND3_X2 c7170(
.A1(net7569),
.A2(net7520),
.A3(net11562),
.ZN(net7640)
);

OR2_X4 c7171(
.A1(net7635),
.A2(net7538),
.ZN(net7641)
);

NOR3_X1 c7172(
.A1(net5694),
.A2(net4729),
.A3(net7608),
.ZN(net7642)
);

OR3_X2 c7173(
.A1(net7495),
.A2(net7621),
.A3(net7609),
.ZN(net7643)
);

OAI21_X2 c7174(
.A(net7621),
.B1(net7506),
.B2(net7488),
.ZN(net7644)
);

OR2_X1 c7175(
.A1(net7636),
.A2(net6689),
.ZN(net7645)
);

OAI21_X1 c7176(
.A(net7632),
.B1(net7621),
.B2(net5706),
.ZN(net7646)
);

XNOR2_X2 c7177(
.A(net7612),
.B(net7577),
.ZN(net7647)
);

DFFRS_X1 c7178(
.D(net7622),
.RN(net7640),
.SN(net5739),
.CK(clk),
.Q(net7649),
.QN(net7648)
);

DFFRS_X2 c7179(
.D(net6710),
.RN(net6654),
.SN(net6689),
.CK(clk),
.Q(net7651),
.QN(net7650)
);

AND2_X4 c7180(
.A1(net7639),
.A2(net10654),
.ZN(net7652)
);

AOI21_X2 c7181(
.A(net7489),
.B1(net5646),
.B2(net6558),
.ZN(net7653)
);

SDFF_X1 c7182(
.D(net6570),
.SE(net7636),
.SI(net5676),
.CK(clk),
.Q(net7655),
.QN(net7654)
);

AOI21_X1 c7183(
.A(net7653),
.B1(net7648),
.B2(net11389),
.ZN(net7656)
);

INV_X8 c7184(
.A(net10309),
.ZN(net7657)
);

AOI21_X4 c7185(
.A(net7619),
.B1(net7559),
.B2(net6569),
.ZN(net7658)
);

AND2_X1 c7186(
.A1(net7629),
.A2(net7616),
.ZN(net7659)
);

AND3_X1 c7187(
.A1(net6632),
.A2(net7654),
.A3(net7640),
.ZN(net7660)
);

NAND3_X1 c7188(
.A1(net6631),
.A2(net7655),
.A3(net7630),
.ZN(net7661)
);

NAND2_X1 c7189(
.A1(net4720),
.A2(net7648),
.ZN(net7662)
);

NOR3_X4 c7190(
.A1(net7639),
.A2(net7662),
.A3(net5669),
.ZN(net7663)
);

NAND2_X2 c7191(
.A1(net7539),
.A2(net7611),
.ZN(net7664)
);

NOR3_X2 c7192(
.A1(net7655),
.A2(net6636),
.A3(net7650),
.ZN(net7665)
);

NAND2_X4 c7193(
.A1(net7665),
.A2(net7624),
.ZN(net7666)
);

AND2_X2 c7194(
.A1(net7652),
.A2(net7631),
.ZN(net7667)
);

OAI221_X1 c7195(
.A(net7623),
.B1(net7608),
.B2(net7578),
.C1(net4741),
.C2(net7633),
.ZN(net7668)
);

SDFF_X2 c7196(
.D(net5586),
.SE(net7662),
.SI(net7578),
.CK(clk),
.Q(net7670),
.QN(net7669)
);

XOR2_X1 c7197(
.A(net7657),
.B(net7659),
.Z(net7671)
);

AND3_X4 c7198(
.A1(net7671),
.A2(net7577),
.A3(net10837),
.ZN(net7672)
);

NAND3_X2 c7199(
.A1(net7630),
.A2(net7616),
.A3(net6682),
.ZN(net7673)
);

NOR2_X1 c7200(
.A1(net7644),
.A2(net7666),
.ZN(net7674)
);

OR2_X2 c7201(
.A1(net7647),
.A2(net7670),
.ZN(net7675)
);

INV_X16 c7202(
.A(net9953),
.ZN(net7676)
);

NOR2_X4 c7203(
.A1(net7671),
.A2(net7670),
.ZN(net7677)
);

OR3_X1 c7204(
.A1(net7666),
.A2(net6679),
.A3(net10653),
.ZN(net7678)
);

MUX2_X1 c7205(
.A(net5688),
.B(net7677),
.S(net7578),
.Z(net7679)
);

AOI222_X2 c7206(
.A1(net7555),
.A2(net6711),
.B1(net7673),
.B2(net7654),
.C1(net7559),
.C2(net7669),
.ZN(net7680)
);

OAI21_X4 c7207(
.A(net6615),
.B1(net7633),
.B2(net10862),
.ZN(net7681)
);

INV_X32 c7208(
.A(net11227),
.ZN(net7682)
);

MUX2_X2 c7209(
.A(net7637),
.B(net7578),
.S(net7641),
.Z(net7683)
);

OAI22_X4 c7210(
.A1(net7680),
.A2(net7615),
.B1(net7673),
.B2(net11226),
.ZN(net7684)
);

SDFFRS_X1 c7211(
.D(net2799),
.RN(net7630),
.SE(net7673),
.SI(net5553),
.SN(net11205),
.CK(clk),
.Q(net7686),
.QN(net7685)
);

NOR2_X2 c7212(
.A1(net5574),
.A2(net4720),
.ZN(net7687)
);

NAND3_X4 c7213(
.A1(net5646),
.A2(net7651),
.A3(net7532),
.ZN(net7688)
);

XOR2_X2 c7214(
.A(net7681),
.B(net7678),
.Z(net7689)
);

OR3_X4 c7215(
.A1(net7687),
.A2(net7662),
.A3(net10741),
.ZN(net7690)
);

AND3_X2 c7216(
.A1(net5707),
.A2(net7651),
.A3(net7639),
.ZN(net7691)
);

XNOR2_X1 c7217(
.A(net7613),
.B(net7675),
.ZN(net7692)
);

OR2_X4 c7218(
.A1(net7691),
.A2(net11088),
.ZN(net7693)
);

OAI222_X1 c7219(
.A1(net7656),
.A2(net6646),
.B1(net7630),
.B2(net6694),
.C1(net7693),
.C2(net7673),
.ZN(net7694)
);

NOR3_X1 c7220(
.A1(net7625),
.A2(net7650),
.A3(net11145),
.ZN(net7695)
);

OR3_X2 c7221(
.A1(net5803),
.A2(net7686),
.A3(net7638),
.ZN(out19)
);

DFFRS_X1 c7222(
.D(net4846),
.RN(net6803),
.SN(net7634),
.CK(clk),
.Q(net7697),
.QN(net7696)
);

OR2_X1 c7223(
.A1(net6690),
.A2(net7634),
.ZN(net7698)
);

OAI21_X2 c7224(
.A(net3876),
.B1(net5623),
.B2(net5759),
.ZN(net7699)
);

OAI21_X1 c7225(
.A(net7545),
.B1(net6743),
.B2(net5730),
.ZN(net7700)
);

AOI21_X2 c7226(
.A(net6782),
.B1(net7676),
.B2(net6772),
.ZN(net7701)
);

AOI21_X1 c7227(
.A(net1857),
.B1(net7618),
.B2(net5792),
.ZN(net7702)
);

AOI21_X4 c7228(
.A(net4704),
.B1(net7700),
.B2(net6732),
.ZN(net7703)
);

DFFRS_X2 c7229(
.D(net5818),
.RN(net7641),
.SN(net7269),
.CK(clk),
.Q(net7705),
.QN(net7704)
);

INV_X4 c7230(
.A(net9709),
.ZN(net7706)
);

AND3_X1 c7231(
.A1(net7617),
.A2(net7533),
.A3(net7638),
.ZN(net7707)
);

NAND3_X1 c7232(
.A1(net6646),
.A2(net5739),
.A3(net3497),
.ZN(net7708)
);

NOR3_X4 c7233(
.A1(net4819),
.A2(net7697),
.A3(net6743),
.ZN(net7709)
);

SDFF_X1 c7234(
.D(net6762),
.SE(net6643),
.SI(net6803),
.CK(clk),
.Q(net7711),
.QN(net7710)
);

NOR3_X2 c7235(
.A1(net6780),
.A2(net6735),
.A3(net7685),
.ZN(net7712)
);

AND3_X4 c7236(
.A1(net6743),
.A2(net7633),
.A3(net10740),
.ZN(out8)
);

NAND3_X2 c7237(
.A1(net7709),
.A2(net7685),
.A3(net6743),
.ZN(net7713)
);

OR3_X1 c7238(
.A1(net4832),
.A2(net6762),
.A3(net5716),
.ZN(net7714)
);

MUX2_X1 c7239(
.A(net3849),
.B(net7710),
.S(net4592),
.Z(net7715)
);

OAI21_X4 c7240(
.A(net6694),
.B1(net6743),
.B2(net7669),
.ZN(out9)
);

MUX2_X2 c7241(
.A(net7618),
.B(net6643),
.S(net6765),
.Z(net7716)
);

NAND3_X4 c7242(
.A1(net7432),
.A2(net5553),
.A3(net7696),
.ZN(net7717)
);

OR3_X4 c7243(
.A1(net7638),
.A2(net7617),
.A3(out9),
.ZN(net7718)
);

AND3_X2 c7244(
.A1(net7715),
.A2(net5739),
.A3(net7582),
.ZN(net7719)
);

NOR3_X1 c7245(
.A1(net5754),
.A2(net7545),
.A3(net6734),
.ZN(net7720)
);

OR3_X2 c7246(
.A1(net6752),
.A2(net2713),
.A3(net7716),
.ZN(net7721)
);

OAI21_X2 c7247(
.A(net7711),
.B1(net6733),
.B2(net5730),
.ZN(net7722)
);

XNOR2_X2 c7248(
.A(net6746),
.B(net6766),
.ZN(net7723)
);

OAI21_X1 c7249(
.A(net7698),
.B1(net6762),
.B2(net7720),
.ZN(net7724)
);

AOI21_X2 c7250(
.A(net6486),
.B1(net7546),
.B2(net6690),
.ZN(net7725)
);

SDFFRS_X2 c7251(
.D(net7624),
.RN(net7676),
.SE(net6780),
.SI(net6730),
.SN(net6788),
.CK(clk),
.Q(net7727),
.QN(net7726)
);

SDFF_X2 c7252(
.D(net5483),
.SE(net7533),
.SI(net7633),
.CK(clk),
.Q(net7729),
.QN(net7728)
);

AOI21_X1 c7253(
.A(net3692),
.B1(net7725),
.B2(net3838),
.ZN(net7730)
);

AOI21_X4 c7254(
.A(net6731),
.B1(net4853),
.B2(net4845),
.ZN(net7731)
);

AND3_X1 c7255(
.A1(net5730),
.A2(net5795),
.A3(net7696),
.ZN(net7732)
);

NAND3_X1 c7256(
.A1(net6807),
.A2(net7728),
.A3(net11164),
.ZN(net7733)
);

NOR3_X4 c7257(
.A1(net5702),
.A2(net7726),
.A3(net11099),
.ZN(net7734)
);

OAI221_X4 c7258(
.A(net7733),
.B1(net6607),
.B2(net6782),
.C1(net7582),
.C2(net6730),
.ZN(net7735)
);

NOR3_X2 c7259(
.A1(net5744),
.A2(net4792),
.A3(net7624),
.ZN(net7736)
);

AND3_X4 c7260(
.A1(net7731),
.A2(net7634),
.A3(net6646),
.ZN(net7737)
);

NAND3_X2 c7261(
.A1(net7706),
.A2(net7716),
.A3(net3828),
.ZN(net7738)
);

OR3_X1 c7262(
.A1(net7705),
.A2(net6754),
.A3(net7728),
.ZN(net7739)
);

DFFRS_X1 c7263(
.D(net7734),
.RN(net7721),
.SN(net1857),
.CK(clk),
.Q(net7741),
.QN(net7740)
);

SDFFRS_X1 c7264(
.D(net7703),
.RN(net7432),
.SE(net1599),
.SI(out9),
.SN(net5759),
.CK(clk),
.Q(net7743),
.QN(net7742)
);

MUX2_X1 c7265(
.A(net4804),
.B(net7727),
.S(net7682),
.Z(net7744)
);

OAI21_X4 c7266(
.A(net7741),
.B1(net7720),
.B2(net10992),
.ZN(net7745)
);

MUX2_X2 c7267(
.A(net7591),
.B(net7737),
.S(net7716),
.Z(net7746)
);

NAND3_X4 c7268(
.A1(net6807),
.A2(net7741),
.A3(net6754),
.ZN(net7747)
);

OR3_X4 c7269(
.A1(net2848),
.A2(net7723),
.A3(out1),
.ZN(net7748)
);

AND3_X2 c7270(
.A1(net7729),
.A2(net7746),
.A3(net7726),
.ZN(net7749)
);

NOR3_X1 c7271(
.A1(net5716),
.A2(net7744),
.A3(net4819),
.ZN(net7750)
);

INV_X1 c7272(
.A(net9708),
.ZN(net7751)
);

DFFRS_X2 c7273(
.D(net6533),
.RN(net7741),
.SN(net7729),
.CK(clk),
.Q(net7753),
.QN(net7752)
);

AND2_X4 c7274(
.A1(net7682),
.A2(net7752),
.ZN(net7754)
);

OR3_X2 c7275(
.A1(net3829),
.A2(net7702),
.A3(net7741),
.ZN(net7755)
);

OAI21_X2 c7276(
.A(net6735),
.B1(net7707),
.B2(net4803),
.ZN(net7756)
);

OAI21_X1 c7277(
.A(net7724),
.B1(net7753),
.B2(net4592),
.ZN(net7757)
);

AOI21_X2 c7278(
.A(net6648),
.B1(net5754),
.B2(net6752),
.ZN(net7758)
);

AOI21_X1 c7279(
.A(net7714),
.B1(net3838),
.B2(net6789),
.ZN(net7759)
);

AOI21_X4 c7280(
.A(net6648),
.B1(net11155),
.B2(net11160),
.ZN(net7760)
);

AND3_X1 c7281(
.A1(net7760),
.A2(net5834),
.A3(net5817),
.ZN(net7761)
);

SDFF_X1 c7282(
.D(net6731),
.SE(net2894),
.SI(net11198),
.CK(clk),
.Q(net7763),
.QN(net7762)
);

NAND3_X1 c7283(
.A1(net4853),
.A2(net6789),
.A3(out9),
.ZN(net7764)
);

SDFF_X2 c7284(
.D(net7730),
.SE(net7743),
.SI(net7762),
.CK(clk),
.Q(net7766),
.QN(net7765)
);

NOR3_X4 c7285(
.A1(net5759),
.A2(net6732),
.A3(net10724),
.ZN(net7767)
);

AND2_X1 c7286(
.A1(net7750),
.A2(net7761),
.ZN(net7768)
);

NOR3_X2 c7287(
.A1(net7766),
.A2(net7754),
.A3(net11225),
.ZN(net7769)
);

AND3_X4 c7288(
.A1(net7718),
.A2(net7763),
.A3(net10993),
.ZN(net7770)
);

NAND3_X2 c7289(
.A1(net7768),
.A2(net7770),
.A3(net7765),
.ZN(net7771)
);

AOI22_X2 c7290(
.A1(net7708),
.A2(net7747),
.B1(net7770),
.B2(net7728),
.ZN(net7772)
);

OAI221_X2 c7291(
.A(net7758),
.B1(net7765),
.B2(net7770),
.C1(out9),
.C2(net10511),
.ZN(net7773)
);

AOI221_X4 c7292(
.A(net5759),
.B1(net7729),
.B2(net7770),
.C1(net7633),
.C2(net10512),
.ZN(net7774)
);

OR3_X1 c7293(
.A1(net7769),
.A2(net6782),
.A3(net11121),
.ZN(net7775)
);

MUX2_X1 c7294(
.A(net7763),
.B(net7745),
.S(net7740),
.Z(net7776)
);

OAI21_X4 c7295(
.A(net7716),
.B1(net6195),
.B2(net11112),
.ZN(net7777)
);

MUX2_X2 c7296(
.A(net6731),
.B(net10954),
.S(net11287),
.Z(net7778)
);

NAND3_X4 c7297(
.A1(net7751),
.A2(net7704),
.A3(net11264),
.ZN(net7779)
);

OR3_X4 c7298(
.A1(net7738),
.A2(net7740),
.A3(net11241),
.ZN(net7780)
);

DFFRS_X1 c7299(
.D(net7776),
.RN(net7762),
.SN(net11545),
.CK(clk),
.Q(net7782),
.QN(net7781)
);

SDFFS_X1 c7300(
.D(net4827),
.SE(net7756),
.SI(net7733),
.SN(net7740),
.CK(clk),
.Q(net7784),
.QN(net7783)
);

OAI222_X4 c7301(
.A1(net7697),
.A2(net7783),
.B1(net6779),
.B2(net6694),
.C1(net6803),
.C2(net11165),
.ZN(net7785)
);

AND3_X2 c7302(
.A1(net7764),
.A2(net5483),
.A3(net11199),
.ZN(net7786)
);

AOI221_X2 c7303(
.A(net4804),
.B1(net6731),
.B2(net7633),
.C1(net11167),
.C2(net11288),
.ZN(net7787)
);

NAND2_X1 c7304(
.A1(net6842),
.A2(net6863),
.ZN(net7788)
);

INV_X2 c7305(
.A(net4874),
.ZN(net7789)
);

INV_X8 c7306(
.A(net6852),
.ZN(net7790)
);

INV_X16 c7307(
.A(net6835),
.ZN(net7791)
);

NAND2_X2 c7308(
.A1(net7789),
.A2(net2928),
.ZN(net7792)
);

INV_X32 c7309(
.A(net6876),
.ZN(net7793)
);

NAND2_X4 c7310(
.A1(net6892),
.A2(net5885),
.ZN(net7794)
);

AND2_X2 c7311(
.A1(net7788),
.A2(net6823),
.ZN(net7795)
);

XOR2_X1 c7312(
.A(net5899),
.B(net6819),
.Z(net7796)
);

INV_X4 c7313(
.A(net7793),
.ZN(net7797)
);

INV_X1 c7314(
.A(net6844),
.ZN(net7798)
);

NOR3_X1 c7315(
.A1(net6811),
.A2(net6810),
.A3(net7796),
.ZN(net7799)
);

INV_X2 c7316(
.A(net9739),
.ZN(net7800)
);

INV_X8 c7317(
.A(net6836),
.ZN(net7801)
);

INV_X16 c7318(
.A(net6810),
.ZN(net7802)
);

INV_X32 c7319(
.A(net5905),
.ZN(net7803)
);

INV_X4 c7320(
.A(net4902),
.ZN(net7804)
);

INV_X1 c7321(
.A(net6888),
.ZN(net7805)
);

NOR2_X1 c7322(
.A1(net5919),
.A2(net6810),
.ZN(net7806)
);

OR2_X2 c7323(
.A1(net4905),
.A2(net6867),
.ZN(net7807)
);

NOR2_X4 c7324(
.A1(net7801),
.A2(net6874),
.ZN(net7808)
);

INV_X2 c7325(
.A(net9817),
.ZN(net7809)
);

DFFRS_X2 c7326(
.D(net6875),
.RN(net5854),
.SN(net1922),
.CK(clk),
.Q(net7811),
.QN(net7810)
);

NOR2_X2 c7327(
.A1(net2928),
.A2(net4862),
.ZN(net7812)
);

INV_X8 c7328(
.A(net10548),
.ZN(net7813)
);

XOR2_X2 c7329(
.A(net6863),
.B(net4902),
.Z(net7814)
);

INV_X16 c7330(
.A(net7791),
.ZN(net7815)
);

DFFR_X1 c7331(
.D(net6811),
.RN(net6822),
.CK(clk),
.Q(net7817),
.QN(net7816)
);

INV_X32 c7332(
.A(net7813),
.ZN(net7818)
);

SDFF_X1 c7333(
.D(net7788),
.SE(net6829),
.SI(net7796),
.CK(clk),
.Q(net7820),
.QN(net7819)
);

XNOR2_X1 c7334(
.A(net7797),
.B(net7801),
.ZN(net7821)
);

OR2_X4 c7335(
.A1(net5837),
.A2(net7802),
.ZN(net7822)
);

INV_X4 c7336(
.A(net9839),
.ZN(net7823)
);

INV_X1 c7337(
.A(net9947),
.ZN(net7824)
);

OR2_X1 c7338(
.A1(net6888),
.A2(net7791),
.ZN(net7825)
);

INV_X2 c7339(
.A(net10549),
.ZN(net7826)
);

INV_X8 c7340(
.A(net7794),
.ZN(net7827)
);

INV_X16 c7341(
.A(net5870),
.ZN(net7828)
);

INV_X32 c7342(
.A(net7826),
.ZN(net7829)
);

OR3_X2 c7343(
.A1(net7813),
.A2(net7820),
.A3(net6842),
.ZN(net7830)
);

INV_X4 c7344(
.A(net7823),
.ZN(net7831)
);

INV_X1 c7345(
.A(net7794),
.ZN(net7832)
);

INV_X2 c7346(
.A(net9946),
.ZN(net7833)
);

XNOR2_X2 c7347(
.A(net7806),
.B(net6898),
.ZN(net7834)
);

AND2_X4 c7348(
.A1(net6813),
.A2(net6885),
.ZN(net7835)
);

INV_X8 c7349(
.A(net7809),
.ZN(net7836)
);

DFFR_X2 c7350(
.D(net7822),
.RN(net6851),
.CK(clk),
.Q(net7838),
.QN(net7837)
);

DFFS_X1 c7351(
.D(net7836),
.SN(net7834),
.CK(clk),
.Q(net7840),
.QN(net7839)
);

NAND4_X4 c7352(
.A1(net7840),
.A2(net7788),
.A3(net7818),
.A4(net6872),
.ZN(net7841)
);

AND2_X1 c7353(
.A1(net5857),
.A2(net7801),
.ZN(net7842)
);

OAI21_X2 c7354(
.A(net7808),
.B1(net7821),
.B2(net7839),
.ZN(net7843)
);

INV_X16 c7355(
.A(net7811),
.ZN(net7844)
);

INV_X32 c7356(
.A(net7844),
.ZN(net7845)
);

DFFS_X2 c7357(
.D(net7837),
.SN(net5883),
.CK(clk),
.Q(net7847),
.QN(net7846)
);

INV_X4 c7358(
.A(net7830),
.ZN(net7848)
);

INV_X1 c7359(
.A(net10006),
.ZN(net7849)
);

INV_X2 c7360(
.A(net7802),
.ZN(net7850)
);

OAI21_X1 c7361(
.A(net7815),
.B1(net7836),
.B2(net7843),
.ZN(net7851)
);

DFFR_X1 c7362(
.D(net7832),
.RN(net6886),
.CK(clk),
.Q(net7853),
.QN(net7852)
);

INV_X8 c7363(
.A(net9738),
.ZN(net7854)
);

NAND2_X1 c7364(
.A1(net7818),
.A2(net7835),
.ZN(net7855)
);

NAND2_X2 c7365(
.A1(net7855),
.A2(net6840),
.ZN(net7856)
);

AOI21_X2 c7366(
.A(net7855),
.B1(net7835),
.B2(net7844),
.ZN(net7857)
);

OAI222_X2 c7367(
.A1(net7857),
.A2(net7851),
.B1(net7842),
.B2(net6846),
.C1(net7792),
.C2(net7796),
.ZN(net7858)
);

OAI211_X2 c7368(
.A(net5847),
.B(net5919),
.C1(net7845),
.C2(net7836),
.ZN(net7859)
);

DFFR_X2 c7369(
.D(net7827),
.RN(net7836),
.CK(clk),
.Q(net7861),
.QN(net7860)
);

AOI21_X1 c7370(
.A(net7861),
.B1(net7825),
.B2(net11565),
.ZN(net7862)
);

AOI21_X4 c7371(
.A(net7856),
.B1(net7831),
.B2(net7810),
.ZN(net7863)
);

DFFS_X1 c7372(
.D(net7834),
.SN(net7792),
.CK(clk),
.Q(net7865),
.QN(net7864)
);

SDFF_X2 c7373(
.D(net7863),
.SE(net7856),
.SI(net11564),
.CK(clk),
.Q(net7867),
.QN(net7866)
);

SDFFRS_X2 c7374(
.D(net7841),
.RN(net7825),
.SE(net7812),
.SI(net7819),
.SN(net7836),
.CK(clk),
.Q(net7869),
.QN(net7868)
);

AND3_X1 c7375(
.A1(net7859),
.A2(net7861),
.A3(net7836),
.ZN(net7870)
);

DFFRS_X1 c7376(
.D(net7854),
.RN(net6899),
.SN(net7870),
.CK(clk),
.Q(net7872),
.QN(net7871)
);

DFFS_X2 c7377(
.D(net7865),
.SN(net7870),
.CK(clk),
.Q(net7874),
.QN(net7873)
);

NAND2_X4 c7378(
.A1(net7838),
.A2(net7871),
.ZN(net7875)
);

DFFR_X1 c7379(
.D(net7842),
.RN(net7846),
.CK(clk),
.Q(net7877),
.QN(net7876)
);

NAND3_X1 c7380(
.A1(net7826),
.A2(net7872),
.A3(net7854),
.ZN(net7878)
);

AOI222_X1 c7381(
.A1(net4929),
.A2(net7863),
.B1(net7875),
.B2(net7819),
.C1(net7836),
.C2(net949),
.ZN(net7879)
);

NOR3_X4 c7382(
.A1(net7872),
.A2(net7827),
.A3(net11566),
.ZN(net7880)
);

DFFRS_X2 c7383(
.D(net7869),
.RN(net7803),
.SN(net10746),
.CK(clk),
.Q(net7882),
.QN(net7881)
);

NOR3_X2 c7384(
.A1(net7876),
.A2(net7852),
.A3(net11567),
.ZN(net7883)
);

AND3_X4 c7385(
.A1(net7824),
.A2(net7883),
.A3(net7866),
.ZN(net7884)
);

NAND3_X2 c7386(
.A1(net7874),
.A2(net7868),
.A3(net7876),
.ZN(net7885)
);

INV_X16 c7387(
.A(net4984),
.ZN(net7886)
);

INV_X32 c7388(
.A(net6958),
.ZN(net7887)
);

INV_X4 c7389(
.A(net6901),
.ZN(net7888)
);

AND2_X2 c7390(
.A1(net4043),
.A2(net6980),
.ZN(net7889)
);

INV_X1 c7391(
.A(net9829),
.ZN(net7890)
);

INV_X2 c7392(
.A(net6829),
.ZN(net7891)
);

XOR2_X1 c7393(
.A(net6865),
.B(net7884),
.Z(net7892)
);

OR3_X1 c7394(
.A1(net7873),
.A2(net7825),
.A3(net6963),
.ZN(net7893)
);

INV_X8 c7395(
.A(net6835),
.ZN(net7894)
);

INV_X16 c7396(
.A(net9655),
.ZN(net7895)
);

INV_X32 c7397(
.A(net5937),
.ZN(net7896)
);

SDFF_X1 c7398(
.D(net7894),
.SE(net7798),
.SI(net11050),
.CK(clk),
.Q(net7898),
.QN(net7897)
);

INV_X4 c7399(
.A(net9654),
.ZN(net7899)
);

NOR2_X1 c7400(
.A1(net7865),
.A2(net5912),
.ZN(net7900)
);

INV_X1 c7401(
.A(net6018),
.ZN(net7901)
);

OR2_X2 c7402(
.A1(net7824),
.A2(net6017),
.ZN(net7902)
);

INV_X2 c7403(
.A(net949),
.ZN(net7903)
);

INV_X8 c7404(
.A(net7888),
.ZN(net7904)
);

NOR2_X4 c7405(
.A1(net7898),
.A2(net7903),
.ZN(net7905)
);

NOR2_X2 c7406(
.A1(net6010),
.A2(net6829),
.ZN(net7906)
);

INV_X16 c7407(
.A(net9891),
.ZN(net7907)
);

INV_X32 c7408(
.A(net3909),
.ZN(net7908)
);

INV_X4 c7409(
.A(net7908),
.ZN(net7909)
);

MUX2_X1 c7410(
.A(net5024),
.B(net6018),
.S(net7897),
.Z(net7910)
);

INV_X1 c7411(
.A(net10436),
.ZN(net7911)
);

INV_X2 c7412(
.A(net6924),
.ZN(net7912)
);

XOR2_X2 c7413(
.A(net7909),
.B(net5953),
.Z(net7913)
);

XNOR2_X1 c7414(
.A(net6823),
.B(net6960),
.ZN(net7914)
);

INV_X8 c7415(
.A(net10137),
.ZN(net7915)
);

INV_X16 c7416(
.A(net10040),
.ZN(net7916)
);

OAI21_X4 c7417(
.A(net7833),
.B1(net7910),
.B2(net5839),
.ZN(net7917)
);

MUX2_X2 c7418(
.A(net7901),
.B(net7903),
.S(net6819),
.Z(net7918)
);

OR2_X4 c7419(
.A1(net7891),
.A2(net7864),
.ZN(net7919)
);

INV_X32 c7420(
.A(net10462),
.ZN(net7920)
);

INV_X4 c7421(
.A(net7895),
.ZN(net7921)
);

INV_X1 c7422(
.A(net7912),
.ZN(net7922)
);

OR2_X1 c7423(
.A1(net7921),
.A2(net7889),
.ZN(net7923)
);

INV_X2 c7424(
.A(net7790),
.ZN(net7924)
);

XNOR2_X2 c7425(
.A(net7906),
.B(net6010),
.ZN(net7925)
);

NAND3_X4 c7426(
.A1(net7893),
.A2(net7790),
.A3(net7833),
.ZN(net7926)
);

INV_X8 c7427(
.A(net6819),
.ZN(net7927)
);

INV_X16 c7428(
.A(net6901),
.ZN(net7928)
);

INV_X32 c7429(
.A(net7914),
.ZN(net7929)
);

OR3_X4 c7430(
.A1(net4953),
.A2(net7886),
.A3(net7909),
.ZN(net7930)
);

INV_X4 c7431(
.A(net7902),
.ZN(net7931)
);

AND2_X4 c7432(
.A1(net7899),
.A2(net6917),
.ZN(net7932)
);

AND2_X1 c7433(
.A1(net7924),
.A2(net7930),
.ZN(net7933)
);

INV_X1 c7434(
.A(net7929),
.ZN(net7934)
);

NAND2_X1 c7435(
.A1(net7930),
.A2(net7878),
.ZN(net7935)
);

NAND2_X2 c7436(
.A1(net7890),
.A2(net6924),
.ZN(net7936)
);

AND3_X2 c7437(
.A1(net7884),
.A2(net7929),
.A3(net6980),
.ZN(net7937)
);

INV_X2 c7438(
.A(net7878),
.ZN(net7938)
);

NAND2_X4 c7439(
.A1(net7935),
.A2(net7926),
.ZN(net7939)
);

AND2_X2 c7440(
.A1(net7905),
.A2(net7934),
.ZN(net7940)
);

XOR2_X1 c7441(
.A(net6917),
.B(net7930),
.Z(net7941)
);

INV_X8 c7442(
.A(net7934),
.ZN(net7942)
);

NOR2_X1 c7443(
.A1(net7932),
.A2(net7926),
.ZN(net7943)
);

OR2_X2 c7444(
.A1(net5967),
.A2(net5945),
.ZN(net7944)
);

DFFR_X2 c7445(
.D(net7918),
.RN(net7808),
.CK(clk),
.Q(net7946),
.QN(net7945)
);

NOR2_X4 c7446(
.A1(net7929),
.A2(net7944),
.ZN(net7947)
);

NOR2_X2 c7447(
.A1(net7821),
.A2(net7942),
.ZN(net7948)
);

INV_X16 c7448(
.A(net7916),
.ZN(net7949)
);

XOR2_X2 c7449(
.A(net7943),
.B(net7937),
.Z(net7950)
);

INV_X32 c7450(
.A(net7931),
.ZN(net7951)
);

XNOR2_X1 c7451(
.A(net7950),
.B(net7896),
.ZN(net7952)
);

OR2_X4 c7452(
.A1(net7938),
.A2(net7952),
.ZN(net7953)
);

NOR3_X1 c7453(
.A1(net7887),
.A2(net7951),
.A3(net6983),
.ZN(net7954)
);

INV_X4 c7454(
.A(net10276),
.ZN(net7955)
);

SDFFS_X2 c7455(
.D(net7937),
.SE(net7945),
.SI(net7942),
.SN(net7796),
.CK(clk),
.Q(net7957),
.QN(net7956)
);

OR2_X1 c7456(
.A1(net7952),
.A2(net7942),
.ZN(net7958)
);

OR4_X2 c7457(
.A1(net7946),
.A2(net7849),
.A3(net6921),
.A4(net7903),
.ZN(net7959)
);

XNOR2_X2 c7458(
.A(net7793),
.B(net7937),
.ZN(net7960)
);

SDFF_X2 c7459(
.D(net7955),
.SE(net7958),
.SI(net7930),
.CK(clk),
.Q(net7962),
.QN(net7961)
);

OR3_X2 c7460(
.A1(net7941),
.A2(net7952),
.A3(net7944),
.ZN(net7963)
);

OAI21_X2 c7461(
.A(net7896),
.B1(net7943),
.B2(net7944),
.ZN(net7964)
);

AND2_X4 c7462(
.A1(net7947),
.A2(net7805),
.ZN(net7965)
);

AND2_X1 c7463(
.A1(net7923),
.A2(net7961),
.ZN(net7966)
);

OAI21_X1 c7464(
.A(net7910),
.B1(net7951),
.B2(net7965),
.ZN(net7967)
);

AOI21_X2 c7465(
.A(net7954),
.B1(net7946),
.B2(net7926),
.ZN(net7968)
);

NAND2_X1 c7466(
.A1(net7957),
.A2(net10966),
.ZN(net7969)
);

AOI21_X1 c7467(
.A(net147),
.B1(net7969),
.B2(net7965),
.ZN(net7970)
);

SDFFRS_X1 c7468(
.D(net7965),
.RN(net7943),
.SE(net7969),
.SI(net7970),
.SN(net6870),
.CK(clk),
.Q(net7972),
.QN(net7971)
);

AOI221_X1 c7469(
.A(net7904),
.B1(net7969),
.B2(net7970),
.C1(net7971),
.C2(net6980),
.ZN(net7973)
);

INV_X1 c7470(
.A(net9865),
.ZN(net7974)
);

INV_X2 c7471(
.A(net11392),
.ZN(net7975)
);

INV_X8 c7472(
.A(net10332),
.ZN(net7976)
);

DFFRS_X1 c7473(
.D(net7927),
.RN(net7928),
.SN(net6017),
.CK(clk),
.Q(net7978),
.QN(net7977)
);

NAND2_X2 c7474(
.A1(net7062),
.A2(net7978),
.ZN(net7979)
);

INV_X16 c7475(
.A(net7004),
.ZN(net7980)
);

INV_X32 c7476(
.A(net7861),
.ZN(net7981)
);

NAND2_X4 c7477(
.A1(net7882),
.A2(net7981),
.ZN(net7982)
);

INV_X4 c7478(
.A(net6042),
.ZN(net7983)
);

INV_X1 c7479(
.A(net7925),
.ZN(net7984)
);

INV_X2 c7480(
.A(net11132),
.ZN(net7985)
);

AND2_X2 c7481(
.A1(net6898),
.A2(net5093),
.ZN(net7986)
);

XOR2_X1 c7482(
.A(net7014),
.B(net7894),
.Z(net7987)
);

INV_X8 c7483(
.A(net9779),
.ZN(net7988)
);

INV_X16 c7484(
.A(net7883),
.ZN(net7989)
);

INV_X32 c7485(
.A(net10274),
.ZN(net7990)
);

NOR2_X1 c7486(
.A1(net7990),
.A2(net7055),
.ZN(net7991)
);

OR2_X2 c7487(
.A1(net6096),
.A2(net7981),
.ZN(net7992)
);

NOR2_X4 c7488(
.A1(net6868),
.A2(net7881),
.ZN(net7993)
);

AOI21_X4 c7489(
.A(net7922),
.B1(net5912),
.B2(net7977),
.ZN(net7994)
);

NOR2_X2 c7490(
.A1(net6062),
.A2(net7860),
.ZN(net7995)
);

XOR2_X2 c7491(
.A(net7055),
.B(net5000),
.Z(net7996)
);

XNOR2_X1 c7492(
.A(net7920),
.B(net6012),
.ZN(net7997)
);

INV_X4 c7493(
.A(net7983),
.ZN(net7998)
);

OR2_X4 c7494(
.A1(net7964),
.A2(net7982),
.ZN(net7999)
);

AND3_X1 c7495(
.A1(net7995),
.A2(net7986),
.A3(net7012),
.ZN(net8000)
);

INV_X1 c7496(
.A(net10005),
.ZN(net8001)
);

OR2_X1 c7497(
.A1(net3976),
.A2(net7997),
.ZN(net8002)
);

INV_X2 c7498(
.A(net9838),
.ZN(net8003)
);

INV_X8 c7499(
.A(net7966),
.ZN(net8004)
);

INV_X16 c7500(
.A(net10345),
.ZN(net8005)
);

XNOR2_X2 c7501(
.A(net7998),
.B(net7987),
.ZN(net8006)
);

AND2_X4 c7502(
.A1(net7951),
.A2(net7978),
.ZN(net8007)
);

INV_X32 c7503(
.A(net10188),
.ZN(net8008)
);

INV_X4 c7504(
.A(net10566),
.ZN(net8009)
);

AND2_X1 c7505(
.A1(net7974),
.A2(net6936),
.ZN(net8010)
);

NAND2_X1 c7506(
.A1(net7994),
.A2(net7052),
.ZN(net8011)
);

NAND3_X1 c7507(
.A1(net6928),
.A2(net7920),
.A3(net7052),
.ZN(net8012)
);

NOR3_X4 c7508(
.A1(net5100),
.A2(net8002),
.A3(net10651),
.ZN(net8013)
);

NAND2_X2 c7509(
.A1(net6985),
.A2(net7974),
.ZN(net8014)
);

INV_X1 c7510(
.A(net10565),
.ZN(net8015)
);

NOR3_X2 c7511(
.A1(net7992),
.A2(net8014),
.A3(net7970),
.ZN(net8016)
);

INV_X2 c7512(
.A(net7989),
.ZN(net8017)
);

AND3_X4 c7513(
.A1(net8001),
.A2(net8002),
.A3(net11377),
.ZN(net8018)
);

INV_X8 c7514(
.A(net10315),
.ZN(net8019)
);

INV_X16 c7515(
.A(net7048),
.ZN(net8020)
);

INV_X32 c7516(
.A(net11331),
.ZN(net8021)
);

NAND2_X4 c7517(
.A1(net6952),
.A2(net6928),
.ZN(net8022)
);

AND2_X2 c7518(
.A1(net6886),
.A2(net7883),
.ZN(net8023)
);

INV_X4 c7519(
.A(net8003),
.ZN(net8024)
);

NAND3_X2 c7520(
.A1(net6998),
.A2(net8016),
.A3(net7820),
.ZN(net8025)
);

XOR2_X1 c7521(
.A(net7903),
.B(net11488),
.Z(net8026)
);

INV_X1 c7522(
.A(net9779),
.ZN(net8027)
);

NOR2_X1 c7523(
.A1(net6054),
.A2(net7850),
.ZN(net8028)
);

OR3_X1 c7524(
.A1(net7862),
.A2(net7037),
.A3(net11243),
.ZN(net8029)
);

OR2_X2 c7525(
.A1(net6845),
.A2(net8019),
.ZN(net8030)
);

NOR2_X4 c7526(
.A1(net7831),
.A2(net8021),
.ZN(net8031)
);

INV_X2 c7527(
.A(net8007),
.ZN(net8032)
);

MUX2_X1 c7528(
.A(net8021),
.B(net8011),
.S(net10521),
.Z(net8033)
);

NOR2_X2 c7529(
.A1(net7991),
.A2(net8021),
.ZN(net8034)
);

AOI211_X1 c7530(
.A(net8032),
.B(net8030),
.C1(net7968),
.C2(net7860),
.ZN(net8035)
);

OAI21_X4 c7531(
.A(net7986),
.B1(net7928),
.B2(net7004),
.ZN(net8036)
);

MUX2_X2 c7532(
.A(net8010),
.B(net7986),
.S(net6993),
.Z(net8037)
);

XOR2_X2 c7533(
.A(net7944),
.B(net7981),
.Z(net8038)
);

XNOR2_X1 c7534(
.A(net8024),
.B(net11377),
.ZN(net8039)
);

INV_X8 c7535(
.A(net8033),
.ZN(net8040)
);

OR2_X4 c7536(
.A1(net8024),
.A2(net10578),
.ZN(net8041)
);

OR2_X1 c7537(
.A1(net8027),
.A2(net11243),
.ZN(net8042)
);

DFFRS_X2 c7538(
.D(net8013),
.RN(net8014),
.SN(net8016),
.CK(clk),
.Q(net8044),
.QN(net8043)
);

XNOR2_X2 c7539(
.A(net8001),
.B(net7980),
.ZN(net8045)
);

NAND3_X4 c7540(
.A1(net6049),
.A2(net8045),
.A3(net8035),
.ZN(net8046)
);

OAI221_X1 c7541(
.A(net7981),
.B1(net8023),
.B2(net5000),
.C1(net7982),
.C2(net7860),
.ZN(net8047)
);

INV_X16 c7542(
.A(net10331),
.ZN(net8048)
);

OR3_X4 c7543(
.A1(net7994),
.A2(net7980),
.A3(net11391),
.ZN(net8049)
);

AND3_X2 c7544(
.A1(net8041),
.A2(net8038),
.A3(net8031),
.ZN(net8050)
);

SDFFR_X1 c7545(
.D(net7986),
.RN(net8043),
.SE(net7041),
.SI(net10761),
.CK(clk),
.Q(net8052),
.QN(net8051)
);

NOR3_X1 c7546(
.A1(net8047),
.A2(net8044),
.A3(net5112),
.ZN(net8053)
);

INV_X32 c7547(
.A(net11392),
.ZN(net8054)
);

AND2_X4 c7548(
.A1(net8049),
.A2(net8054),
.ZN(net8055)
);

NAND4_X2 c7549(
.A1(net7993),
.A2(net8054),
.A3(net8055),
.A4(net5092),
.ZN(net8056)
);

OR3_X2 c7550(
.A1(net7849),
.A2(net7861),
.A3(net11201),
.ZN(net8057)
);

OAI221_X4 c7551(
.A(net7975),
.B1(net8056),
.B2(net8044),
.C1(net8057),
.C2(net7819),
.ZN(net8058)
);

OAI221_X2 c7552(
.A(net8048),
.B1(net8034),
.B2(net8055),
.C1(net8058),
.C2(net7982),
.ZN(net8059)
);

AND2_X1 c7553(
.A1(net7968),
.A2(net7160),
.ZN(net8060)
);

NAND2_X1 c7554(
.A1(net7029),
.A2(net7019),
.ZN(net8061)
);

NAND2_X2 c7555(
.A1(net7926),
.A2(net7988),
.ZN(net8062)
);

NAND2_X4 c7556(
.A1(net8062),
.A2(net8019),
.ZN(net8063)
);

AND2_X2 c7557(
.A1(net7862),
.A2(net7029),
.ZN(net8064)
);

XOR2_X1 c7558(
.A(net6840),
.B(net7907),
.Z(net8065)
);

NOR2_X1 c7559(
.A1(net3201),
.A2(net6104),
.ZN(net8066)
);

OR2_X2 c7560(
.A1(net8063),
.A2(net7980),
.ZN(net8067)
);

NOR2_X4 c7561(
.A1(net8061),
.A2(net8064),
.ZN(net8068)
);

NOR2_X2 c7562(
.A1(net5012),
.A2(net7150),
.ZN(net8069)
);

XOR2_X2 c7563(
.A(net8026),
.B(net6840),
.Z(net8070)
);

INV_X4 c7564(
.A(net10123),
.ZN(net8071)
);

XNOR2_X1 c7565(
.A(net8066),
.B(net8070),
.ZN(net8072)
);

OR2_X4 c7566(
.A1(net8071),
.A2(net8051),
.ZN(net8073)
);

INV_X1 c7567(
.A(net7113),
.ZN(net8074)
);

OAI21_X2 c7568(
.A(net6936),
.B1(net8060),
.B2(net7900),
.ZN(net8075)
);

OR2_X1 c7569(
.A1(net8065),
.A2(net8073),
.ZN(net8076)
);

INV_X2 c7570(
.A(net11250),
.ZN(net8077)
);

XNOR2_X2 c7571(
.A(net6967),
.B(net8021),
.ZN(net8078)
);

AND2_X4 c7572(
.A1(net7939),
.A2(net8011),
.ZN(net8079)
);

AND2_X1 c7573(
.A1(net8073),
.A2(net8061),
.ZN(net8080)
);

NAND2_X1 c7574(
.A1(net8070),
.A2(net8014),
.ZN(net8081)
);

DFFS_X1 c7575(
.D(net7092),
.SN(net7113),
.CK(clk),
.Q(net8083),
.QN(net8082)
);

INV_X8 c7576(
.A(net8075),
.ZN(net8084)
);

INV_X16 c7577(
.A(net7976),
.ZN(net8085)
);

OR4_X4 c7578(
.A1(net8019),
.A2(net7154),
.A3(net7940),
.A4(net7141),
.ZN(net8086)
);

NAND2_X2 c7579(
.A1(net8067),
.A2(net7997),
.ZN(net8087)
);

NAND2_X4 c7580(
.A1(net8083),
.A2(net8085),
.ZN(net8088)
);

AND2_X2 c7581(
.A1(net7011),
.A2(net8045),
.ZN(net8089)
);

XOR2_X1 c7582(
.A(net8068),
.B(net7997),
.Z(net8090)
);

NOR2_X1 c7583(
.A1(net8052),
.A2(net8073),
.ZN(net8091)
);

OR2_X2 c7584(
.A1(net8074),
.A2(net8050),
.ZN(net8092)
);

NOR2_X4 c7585(
.A1(net8064),
.A2(net7088),
.ZN(net8093)
);

NOR2_X2 c7586(
.A1(net8084),
.A2(net7087),
.ZN(net8094)
);

INV_X32 c7587(
.A(net8094),
.ZN(net8095)
);

OAI21_X1 c7588(
.A(net6963),
.B1(net7968),
.B2(net8091),
.ZN(net8096)
);

XOR2_X2 c7589(
.A(net8096),
.B(net7011),
.Z(net8097)
);

AOI21_X2 c7590(
.A(net5000),
.B1(net8082),
.B2(net8062),
.ZN(net8098)
);

INV_X4 c7591(
.A(net10066),
.ZN(net8099)
);

XNOR2_X1 c7592(
.A(net8017),
.B(net8085),
.ZN(net8100)
);

INV_X1 c7593(
.A(net10310),
.ZN(net8101)
);

OR2_X4 c7594(
.A1(net8088),
.A2(net8092),
.ZN(net8102)
);

SDFF_X1 c7595(
.D(net7918),
.SE(net7041),
.SI(net8062),
.CK(clk),
.Q(net8104),
.QN(net8103)
);

OR2_X1 c7596(
.A1(net7041),
.A2(net8035),
.ZN(net8105)
);

SDFF_X2 c7597(
.D(net8102),
.SE(net6963),
.SI(net8012),
.CK(clk),
.Q(net8107),
.QN(net8106)
);

OAI22_X2 c7598(
.A1(net7155),
.A2(net8101),
.B1(net8061),
.B2(net8098),
.ZN(net8108)
);

XNOR2_X2 c7599(
.A(net8034),
.B(net7113),
.ZN(net8109)
);

AND2_X4 c7600(
.A1(net7997),
.A2(net6170),
.ZN(net8110)
);

DFFS_X2 c7601(
.D(net7122),
.SN(net10522),
.CK(clk),
.Q(net8112),
.QN(net8111)
);

AND2_X1 c7602(
.A1(net8069),
.A2(net8109),
.ZN(net8113)
);

NAND2_X1 c7603(
.A1(net7940),
.A2(net8011),
.ZN(net8114)
);

INV_X2 c7604(
.A(net9900),
.ZN(net8115)
);

OAI211_X4 c7605(
.A(net8115),
.B(net5209),
.C1(net6011),
.C2(net8111),
.ZN(net8116)
);

NAND2_X2 c7606(
.A1(net8107),
.A2(net8092),
.ZN(net8117)
);

NAND2_X4 c7607(
.A1(net5209),
.A2(net5113),
.ZN(net8118)
);

AND2_X2 c7608(
.A1(net8089),
.A2(net8109),
.ZN(net8119)
);

XOR2_X1 c7609(
.A(net8086),
.B(net8106),
.Z(net8120)
);

INV_X8 c7610(
.A(net10203),
.ZN(net8121)
);

NOR2_X1 c7611(
.A1(net7936),
.A2(net5012),
.ZN(net8122)
);

OAI211_X1 c7612(
.A(net8072),
.B(net8120),
.C1(net5139),
.C2(net8058),
.ZN(net8123)
);

AOI21_X1 c7613(
.A(net6050),
.B1(net8103),
.B2(net11343),
.ZN(net8124)
);

OR2_X2 c7614(
.A1(net8124),
.A2(net8116),
.ZN(net8125)
);

NOR2_X4 c7615(
.A1(net8015),
.A2(net8085),
.ZN(net8126)
);

SDFFRS_X2 c7616(
.D(net7867),
.RN(net6967),
.SE(net7122),
.SI(net8062),
.SN(net8091),
.CK(clk),
.Q(net8128),
.QN(net8127)
);

INV_X16 c7617(
.A(net11401),
.ZN(net8129)
);

NOR2_X2 c7618(
.A1(net8129),
.A2(net8127),
.ZN(net8130)
);

DFFRS_X1 c7619(
.D(net8101),
.RN(net7122),
.SN(net8116),
.CK(clk),
.Q(net8132),
.QN(net8131)
);

AOI21_X4 c7620(
.A(net5912),
.B1(net7889),
.B2(net8109),
.ZN(net8133)
);

XOR2_X2 c7621(
.A(net8100),
.B(net8132),
.Z(net8134)
);

AND3_X1 c7622(
.A1(net7150),
.A2(net8073),
.A3(net8121),
.ZN(net8135)
);

NAND3_X1 c7623(
.A1(net8078),
.A2(net8133),
.A3(net8131),
.ZN(net8136)
);

AOI222_X4 c7624(
.A1(net8122),
.A2(net8132),
.B1(net5209),
.B2(net8091),
.C1(net7903),
.C2(net11190),
.ZN(net8137)
);

XNOR2_X1 c7625(
.A(net8121),
.B(net8135),
.ZN(net8138)
);

NOR4_X4 c7626(
.A1(net8104),
.A2(net8129),
.A3(net8102),
.A4(net8127),
.ZN(net8139)
);

NOR3_X4 c7627(
.A1(net8138),
.A2(net8135),
.A3(net11437),
.ZN(net8140)
);

INV_X32 c7628(
.A(net11250),
.ZN(net8141)
);

NOR3_X2 c7629(
.A1(net7037),
.A2(net7862),
.A3(net11190),
.ZN(net8142)
);

AND3_X4 c7630(
.A1(net8134),
.A2(net8116),
.A3(net11104),
.ZN(net8143)
);

NOR4_X2 c7631(
.A1(net8133),
.A2(net8130),
.A3(net7078),
.A4(net11105),
.ZN(net8144)
);

OR2_X4 c7632(
.A1(net8114),
.A2(net8143),
.ZN(net8145)
);

NAND3_X2 c7633(
.A1(net8137),
.A2(net8145),
.A3(net8133),
.ZN(net8146)
);

OAI33_X1 c7634(
.A1(net8112),
.A2(net8113),
.A3(net8109),
.B1(net8116),
.B2(net8091),
.B3(net11413),
.ZN(net8147)
);

OR3_X1 c7635(
.A1(net8145),
.A2(net7137),
.A3(net8113),
.ZN(net8148)
);

OR2_X1 c7636(
.A1(net8141),
.A2(net6883),
.ZN(net8149)
);

XNOR2_X2 c7637(
.A(net6187),
.B(net8002),
.ZN(net8150)
);

MUX2_X1 c7638(
.A(net8135),
.B(net7206),
.S(net7915),
.Z(net8151)
);

AND2_X4 c7639(
.A1(net7093),
.A2(net8116),
.ZN(net8152)
);

AOI211_X4 c7640(
.A(net6987),
.B(net5139),
.C1(net6208),
.C2(net6240),
.ZN(net8153)
);

INV_X4 c7641(
.A(net8116),
.ZN(net8154)
);

AND2_X1 c7642(
.A1(net7959),
.A2(net8153),
.ZN(net8155)
);

INV_X1 c7643(
.A(net11459),
.ZN(net8156)
);

NAND2_X1 c7644(
.A1(net7220),
.A2(net8141),
.ZN(net8157)
);

INV_X2 c7645(
.A(net9678),
.ZN(net8158)
);

OAI21_X4 c7646(
.A(net8144),
.B1(net7172),
.B2(net11306),
.ZN(net8159)
);

NAND2_X2 c7647(
.A1(net8135),
.A2(net10815),
.ZN(net8160)
);

NAND2_X4 c7648(
.A1(net7984),
.A2(net8149),
.ZN(net8161)
);

AND2_X2 c7649(
.A1(net6240),
.A2(net10851),
.ZN(net8162)
);

XOR2_X1 c7650(
.A(net8158),
.B(net6165),
.Z(net8163)
);

NOR2_X1 c7651(
.A1(net7178),
.A2(net7175),
.ZN(net8164)
);

OR2_X2 c7652(
.A1(net2276),
.A2(net8085),
.ZN(net8165)
);

INV_X8 c7653(
.A(net8164),
.ZN(net8166)
);

NOR2_X4 c7654(
.A1(net8162),
.A2(net7957),
.ZN(net8167)
);

INV_X16 c7655(
.A(net10229),
.ZN(net8168)
);

NOR2_X2 c7656(
.A1(net8156),
.A2(net7915),
.ZN(net8169)
);

MUX2_X2 c7657(
.A(net7166),
.B(net8110),
.S(net7889),
.Z(net8170)
);

INV_X32 c7658(
.A(net5139),
.ZN(net8171)
);

INV_X4 c7659(
.A(net9945),
.ZN(net8172)
);

INV_X1 c7660(
.A(net11379),
.ZN(net8173)
);

XOR2_X2 c7661(
.A(net6208),
.B(net8045),
.Z(net8174)
);

XNOR2_X1 c7662(
.A(net4322),
.B(net10743),
.ZN(net8175)
);

INV_X2 c7663(
.A(net10418),
.ZN(net8176)
);

OR2_X4 c7664(
.A1(net7252),
.A2(net10912),
.ZN(net8177)
);

OR2_X1 c7665(
.A1(net8163),
.A2(net7900),
.ZN(net8178)
);

DFFR_X1 c7666(
.D(net8042),
.RN(net7253),
.CK(clk),
.Q(net8180),
.QN(net8179)
);

XNOR2_X2 c7667(
.A(net7088),
.B(net8179),
.ZN(net8181)
);

AND2_X4 c7668(
.A1(net8092),
.A2(net7206),
.ZN(net8182)
);

NAND3_X4 c7669(
.A1(net8167),
.A2(net5234),
.A3(net7176),
.ZN(net8183)
);

AND2_X1 c7670(
.A1(net8175),
.A2(net2276),
.ZN(net8184)
);

NAND2_X1 c7671(
.A1(net8040),
.A2(net7251),
.ZN(net8185)
);

OR3_X4 c7672(
.A1(net8170),
.A2(net6165),
.A3(net8178),
.ZN(net8186)
);

NAND2_X2 c7673(
.A1(net8184),
.A2(net7229),
.ZN(net8187)
);

INV_X8 c7674(
.A(net10395),
.ZN(net8188)
);

INV_X16 c7675(
.A(net11351),
.ZN(net8189)
);

NAND2_X4 c7676(
.A1(net7225),
.A2(net8170),
.ZN(net8190)
);

AND3_X2 c7677(
.A1(net8178),
.A2(net8128),
.A3(net8130),
.ZN(net8191)
);

DFFR_X2 c7678(
.D(net8160),
.RN(net7214),
.CK(clk),
.Q(net8193),
.QN(net8192)
);

AND2_X2 c7679(
.A1(net7251),
.A2(net7235),
.ZN(out13)
);

XOR2_X1 c7680(
.A(net8181),
.B(net4904),
.Z(net8194)
);

NOR2_X1 c7681(
.A1(net5282),
.A2(net2276),
.ZN(net8195)
);

OR2_X2 c7682(
.A1(net8189),
.A2(net8195),
.ZN(net8196)
);

NOR2_X4 c7683(
.A1(net8085),
.A2(net8193),
.ZN(net8197)
);

NOR2_X2 c7684(
.A1(net8188),
.A2(net6987),
.ZN(net8198)
);

INV_X32 c7685(
.A(net10042),
.ZN(net8199)
);

DFFS_X1 c7686(
.D(net8182),
.SN(net7911),
.CK(clk),
.Q(net8201),
.QN(net8200)
);

INV_X4 c7687(
.A(net10397),
.ZN(net8202)
);

AOI221_X4 c7688(
.A(net4283),
.B1(net8024),
.B2(net8199),
.C1(net8149),
.C2(net8166),
.ZN(net8203)
);

DFFRS_X2 c7689(
.D(net7796),
.RN(net8196),
.SN(net8195),
.CK(clk),
.Q(net8205),
.QN(net8204)
);

NOR3_X1 c7690(
.A1(net8176),
.A2(net8171),
.A3(net8149),
.ZN(net8206)
);

AOI221_X2 c7691(
.A(net8199),
.B1(net7165),
.B2(net8178),
.C1(out13),
.C2(net8091),
.ZN(net8207)
);

INV_X1 c7692(
.A(net9894),
.ZN(net8208)
);

XOR2_X2 c7693(
.A(net8194),
.B(net8156),
.Z(net8209)
);

XNOR2_X1 c7694(
.A(net8185),
.B(net7175),
.ZN(net8210)
);

INV_X2 c7695(
.A(net10144),
.ZN(net8211)
);

OR2_X4 c7696(
.A1(net8205),
.A2(net8157),
.ZN(net8212)
);

OR3_X2 c7697(
.A1(net7206),
.A2(net8210),
.A3(net8204),
.ZN(net8213)
);

OR2_X1 c7698(
.A1(net8198),
.A2(net7251),
.ZN(net8214)
);

XNOR2_X2 c7699(
.A(net8214),
.B(net8205),
.ZN(net8215)
);

OAI21_X2 c7700(
.A(net8090),
.B1(net8215),
.B2(net6993),
.ZN(net8216)
);

INV_X8 c7701(
.A(net9899),
.ZN(net8217)
);

INV_X16 c7702(
.A(net9677),
.ZN(net8218)
);

OAI21_X1 c7703(
.A(net8203),
.B1(net8198),
.B2(net8212),
.ZN(net8219)
);

AOI21_X2 c7704(
.A(net8168),
.B1(net8079),
.B2(net8197),
.ZN(net8220)
);

AOI21_X1 c7705(
.A(net5222),
.B1(net8213),
.B2(net8150),
.ZN(net8221)
);

AND2_X4 c7706(
.A1(net8211),
.A2(net2276),
.ZN(net8222)
);

AOI21_X4 c7707(
.A(net8209),
.B1(net8202),
.B2(net8194),
.ZN(net8223)
);

AND2_X1 c7708(
.A1(net8218),
.A2(net10518),
.ZN(net8224)
);

AND3_X1 c7709(
.A1(net8197),
.A2(net7228),
.A3(net8223),
.ZN(net8225)
);

NAND3_X1 c7710(
.A1(net7229),
.A2(net8199),
.A3(net8223),
.ZN(net8226)
);

AOI222_X2 c7711(
.A1(net8195),
.A2(net8190),
.B1(net8226),
.B2(net8215),
.C1(net7214),
.C2(net7252),
.ZN(net8227)
);

NOR3_X4 c7712(
.A1(net7960),
.A2(net8219),
.A3(net11570),
.ZN(net8228)
);

NOR3_X2 c7713(
.A1(net8220),
.A2(net8224),
.A3(net8223),
.ZN(net8229)
);

AND3_X4 c7714(
.A1(net8226),
.A2(net8218),
.A3(net8228),
.ZN(net8230)
);

NAND3_X2 c7715(
.A1(net8208),
.A2(net7229),
.A3(net10517),
.ZN(net8231)
);

SDFF_X1 c7716(
.D(net8154),
.SE(net8199),
.SI(net8187),
.CK(clk),
.Q(net8233),
.QN(net8232)
);

OR3_X1 c7717(
.A1(net8191),
.A2(net8233),
.A3(net8090),
.ZN(net8234)
);

OAI222_X1 c7718(
.A1(net8218),
.A2(net8223),
.B1(net8198),
.B2(net8232),
.C1(net7252),
.C2(out13),
.ZN(net8235)
);

INV_X32 c7719(
.A(net5235),
.ZN(net8236)
);

NAND2_X1 c7720(
.A1(net8039),
.A2(net7141),
.ZN(net8237)
);

NAND2_X2 c7721(
.A1(net6293),
.A2(net10770),
.ZN(net8238)
);

NAND2_X4 c7722(
.A1(net7291),
.A2(net7124),
.ZN(net8239)
);

INV_X4 c7723(
.A(net6290),
.ZN(net8240)
);

INV_X1 c7724(
.A(net9744),
.ZN(net8241)
);

AND2_X2 c7725(
.A1(net6012),
.A2(net6293),
.ZN(net8242)
);

XOR2_X1 c7726(
.A(net8020),
.B(net6257),
.Z(net8243)
);

NOR4_X1 c7727(
.A1(net7141),
.A2(net5894),
.A3(net7281),
.A4(net8207),
.ZN(net8244)
);

INV_X2 c7728(
.A(net10088),
.ZN(net8245)
);

NOR2_X1 c7729(
.A1(net7281),
.A2(net7124),
.ZN(net8246)
);

INV_X8 c7730(
.A(net8225),
.ZN(net8247)
);

DFFS_X2 c7731(
.D(net7338),
.SN(net6328),
.CK(clk),
.Q(net8249),
.QN(net8248)
);

OAI222_X4 c7732(
.A1(net8132),
.A2(net7911),
.B1(net7309),
.B2(net7903),
.C1(net7171),
.C2(net8024),
.ZN(net8250)
);

INV_X16 c7733(
.A(net8031),
.ZN(net8251)
);

OR2_X2 c7734(
.A1(net8180),
.A2(net7309),
.ZN(net8252)
);

MUX2_X1 c7735(
.A(net7329),
.B(net7252),
.S(net11366),
.Z(net8253)
);

NOR2_X4 c7736(
.A1(net8245),
.A2(net8242),
.ZN(net8254)
);

INV_X32 c7737(
.A(net9956),
.ZN(net8255)
);

INV_X4 c7738(
.A(net7282),
.ZN(net8256)
);

NOR2_X2 c7739(
.A1(net6328),
.A2(net7124),
.ZN(net8257)
);

INV_X1 c7740(
.A(net9923),
.ZN(net8258)
);

XOR2_X2 c7741(
.A(net8005),
.B(net7277),
.Z(net8259)
);

XNOR2_X1 c7742(
.A(net8011),
.B(net8098),
.ZN(net8260)
);

OR2_X4 c7743(
.A1(net6293),
.A2(net5924),
.ZN(net8261)
);

OR2_X1 c7744(
.A1(net8110),
.A2(net6165),
.ZN(net8262)
);

XNOR2_X2 c7745(
.A(net7336),
.B(net8059),
.ZN(net8263)
);

AND2_X4 c7746(
.A1(net8258),
.A2(net7141),
.ZN(net8264)
);

INV_X2 c7747(
.A(net10286),
.ZN(net8265)
);

INV_X8 c7748(
.A(net9975),
.ZN(net8266)
);

AND2_X1 c7749(
.A1(net8239),
.A2(net8059),
.ZN(net8267)
);

SDFF_X2 c7750(
.D(net8253),
.SE(net7336),
.SI(net8264),
.CK(clk),
.Q(net8269),
.QN(net8268)
);

SDFFR_X2 c7751(
.D(net8263),
.RN(net8002),
.SE(net8127),
.SI(net7171),
.CK(clk),
.Q(net8271),
.QN(net8270)
);

INV_X16 c7752(
.A(net11437),
.ZN(net8272)
);

INV_X32 c7753(
.A(net9924),
.ZN(net8273)
);

DFFR_X1 c7754(
.D(net8254),
.RN(net8157),
.CK(clk),
.Q(net8275),
.QN(net8274)
);

NAND2_X1 c7755(
.A1(net1399),
.A2(net8256),
.ZN(net8276)
);

NAND2_X2 c7756(
.A1(net8262),
.A2(net8240),
.ZN(net8277)
);

INV_X4 c7757(
.A(net11384),
.ZN(net8278)
);

INV_X1 c7758(
.A(net7214),
.ZN(net8279)
);

INV_X2 c7759(
.A(net11383),
.ZN(net8280)
);

INV_X8 c7760(
.A(net8173),
.ZN(net8281)
);

NAND2_X4 c7761(
.A1(net8269),
.A2(net8279),
.ZN(net8282)
);

AND2_X2 c7762(
.A1(net5913),
.A2(net8256),
.ZN(net8283)
);

XOR2_X1 c7763(
.A(net7124),
.B(net8039),
.Z(net8284)
);

NOR2_X1 c7764(
.A1(net6984),
.A2(net8270),
.ZN(net8285)
);

OR2_X2 c7765(
.A1(net8247),
.A2(net8275),
.ZN(net8286)
);

INV_X16 c7766(
.A(net7321),
.ZN(net8287)
);

NOR2_X4 c7767(
.A1(net7172),
.A2(out13),
.ZN(net8288)
);

AOI211_X2 c7768(
.A(net7308),
.B(net8242),
.C1(net8279),
.C2(net8284),
.ZN(net8289)
);

NOR2_X2 c7769(
.A1(net7165),
.A2(net8153),
.ZN(net8290)
);

XOR2_X2 c7770(
.A(net8287),
.B(net11366),
.Z(net8291)
);

XNOR2_X1 c7771(
.A(net8282),
.B(net7252),
.ZN(net8292)
);

INV_X32 c7772(
.A(net10168),
.ZN(net8293)
);

AOI221_X1 c7773(
.A(net7327),
.B1(net8240),
.B2(net8262),
.C1(net7288),
.C2(net8279),
.ZN(net8294)
);

OR2_X4 c7774(
.A1(net8293),
.A2(net8268),
.ZN(net8295)
);

OAI21_X4 c7775(
.A(net8271),
.B1(net8130),
.B2(net8295),
.ZN(net8296)
);

MUX2_X2 c7776(
.A(net8242),
.B(net8293),
.S(net8200),
.Z(net8297)
);

AOI22_X1 c7777(
.A1(net8289),
.A2(net8284),
.B1(net8294),
.B2(net7184),
.ZN(net8298)
);

INV_X4 c7778(
.A(net9847),
.ZN(net8299)
);

INV_X1 c7779(
.A(net11216),
.ZN(net8300)
);

OR2_X1 c7780(
.A1(net8276),
.A2(net6105),
.ZN(net8301)
);

NAND3_X4 c7781(
.A1(net8280),
.A2(net8287),
.A3(net7141),
.ZN(net8302)
);

XNOR2_X2 c7782(
.A(net8153),
.B(net11571),
.ZN(net8303)
);

OR3_X4 c7783(
.A1(net7228),
.A2(net8260),
.A3(net8180),
.ZN(net8304)
);

DFFRS_X1 c7784(
.D(net8266),
.RN(net8301),
.SN(net8289),
.CK(clk),
.Q(net8306),
.QN(net8305)
);

AND2_X4 c7785(
.A1(net8291),
.A2(net8304),
.ZN(net8307)
);

INV_X2 c7786(
.A(net10180),
.ZN(net8308)
);

AND2_X1 c7787(
.A1(net8262),
.A2(net10604),
.ZN(net8309)
);

AND3_X2 c7788(
.A1(net8237),
.A2(net8299),
.A3(net8305),
.ZN(net8310)
);

INV_X8 c7789(
.A(net9743),
.ZN(net8311)
);

NAND2_X1 c7790(
.A1(net8288),
.A2(net7141),
.ZN(net8312)
);

AND4_X4 c7791(
.A1(net8309),
.A2(net8287),
.A3(net8276),
.A4(net7288),
.ZN(net8313)
);

NOR3_X1 c7792(
.A1(net8300),
.A2(net8307),
.A3(net8309),
.ZN(net8314)
);

OR3_X2 c7793(
.A1(net8285),
.A2(net8299),
.A3(net8302),
.ZN(net8315)
);

NAND2_X2 c7794(
.A1(net8315),
.A2(net11028),
.ZN(net8316)
);

NAND4_X1 c7795(
.A1(net8312),
.A2(net8303),
.A3(net8315),
.A4(out13),
.ZN(net8317)
);

OAI21_X2 c7796(
.A(net8273),
.B1(net8276),
.B2(net11434),
.ZN(net8318)
);

OAI21_X1 c7797(
.A(net8314),
.B1(net8311),
.B2(net11434),
.ZN(net8319)
);

OAI222_X2 c7798(
.A1(net8277),
.A2(net8318),
.B1(net8315),
.B2(net8294),
.C1(net7213),
.C2(net8274),
.ZN(net8320)
);

DFFRS_X2 c7799(
.D(net8255),
.RN(net8217),
.SN(net8320),
.CK(clk),
.Q(net8322),
.QN(net8321)
);

OAI221_X1 c7800(
.A(net8240),
.B1(net8314),
.B2(net8321),
.C1(net8315),
.C2(net10603),
.ZN(net8323)
);

OR4_X1 c7801(
.A1(net8308),
.A2(net8318),
.A3(net8314),
.A4(net8321),
.ZN(net8324)
);

NAND2_X4 c7802(
.A1(net7348),
.A2(net7312),
.ZN(net8325)
);

AND2_X2 c7803(
.A1(net6413),
.A2(net7074),
.ZN(net8326)
);

INV_X16 c7804(
.A(net9689),
.ZN(net8327)
);

XOR2_X1 c7805(
.A(net7312),
.B(net8284),
.Z(net8328)
);

NOR2_X1 c7806(
.A1(net556),
.A2(net8264),
.ZN(net8329)
);

AOI21_X2 c7807(
.A(net8302),
.B1(net8294),
.B2(net7363),
.ZN(net8330)
);

AOI21_X1 c7808(
.A(net8260),
.B1(net7296),
.B2(net8128),
.ZN(net8331)
);

OR2_X2 c7809(
.A1(net6454),
.A2(net11261),
.ZN(net8332)
);

INV_X32 c7810(
.A(net10477),
.ZN(net8333)
);

INV_X4 c7811(
.A(net10405),
.ZN(net8334)
);

NOR2_X4 c7812(
.A1(net8334),
.A2(net7300),
.ZN(net8335)
);

NOR2_X2 c7813(
.A1(net7329),
.A2(net7126),
.ZN(net8336)
);

AOI21_X4 c7814(
.A(net8077),
.B1(net7405),
.B2(net6454),
.ZN(net8337)
);

XOR2_X2 c7815(
.A(net8294),
.B(net8024),
.Z(net8338)
);

AND3_X1 c7816(
.A1(net8219),
.A2(net7363),
.A3(net5234),
.ZN(net8339)
);

XNOR2_X1 c7817(
.A(net7393),
.B(net7342),
.ZN(net8340)
);

NAND3_X1 c7818(
.A1(net8290),
.A2(net8335),
.A3(net7329),
.ZN(net8341)
);

OR2_X4 c7819(
.A1(net7418),
.A2(net7405),
.ZN(net8342)
);

INV_X1 c7820(
.A(net10250),
.ZN(net8343)
);

INV_X2 c7821(
.A(net11404),
.ZN(net8344)
);

OR2_X1 c7822(
.A1(net8284),
.A2(net10883),
.ZN(net8345)
);

XNOR2_X2 c7823(
.A(net7409),
.B(net5431),
.ZN(net8346)
);

NOR3_X4 c7824(
.A1(net6165),
.A2(net8335),
.A3(net8012),
.ZN(net8347)
);

DFFR_X2 c7825(
.D(net8331),
.RN(net8330),
.CK(clk),
.Q(net8349),
.QN(net8348)
);

NOR3_X2 c7826(
.A1(net8155),
.A2(net7372),
.A3(net8329),
.ZN(net8350)
);

AND2_X4 c7827(
.A1(net6388),
.A2(net8339),
.ZN(net8351)
);

AND2_X1 c7828(
.A1(net8296),
.A2(net7372),
.ZN(net8352)
);

INV_X8 c7829(
.A(net11381),
.ZN(net8353)
);

INV_X16 c7830(
.A(net9969),
.ZN(net8354)
);

NAND2_X1 c7831(
.A1(net8344),
.A2(net8343),
.ZN(net8355)
);

INV_X32 c7832(
.A(net9876),
.ZN(net8356)
);

AND3_X4 c7833(
.A1(net8177),
.A2(net8356),
.A3(net8353),
.ZN(net8357)
);

NAND2_X2 c7834(
.A1(net5432),
.A2(net8316),
.ZN(net8358)
);

NAND3_X2 c7835(
.A1(net7379),
.A2(net7312),
.A3(net11431),
.ZN(net8359)
);

NAND2_X4 c7836(
.A1(net8002),
.A2(net8345),
.ZN(net8360)
);

INV_X4 c7837(
.A(net11314),
.ZN(net8361)
);

AND2_X2 c7838(
.A1(net8257),
.A2(net8352),
.ZN(net8362)
);

XOR2_X1 c7839(
.A(net7382),
.B(net8077),
.Z(net8363)
);

NOR2_X1 c7840(
.A1(net7296),
.A2(net8355),
.ZN(net8364)
);

OR3_X1 c7841(
.A1(net8157),
.A2(net8329),
.A3(net11166),
.ZN(net8365)
);

MUX2_X1 c7842(
.A(net8236),
.B(net7127),
.S(net8219),
.Z(net8366)
);

OAI21_X4 c7843(
.A(net8363),
.B1(net7356),
.B2(net8329),
.ZN(net8367)
);

OR2_X2 c7844(
.A1(net8250),
.A2(net6363),
.ZN(net8368)
);

NOR2_X4 c7845(
.A1(net7422),
.A2(net5100),
.ZN(net8369)
);

MUX2_X2 c7846(
.A(net6439),
.B(net7296),
.S(net3451),
.Z(net8370)
);

SDFFRS_X1 c7847(
.D(net8259),
.RN(net8330),
.SE(net8274),
.SI(net6437),
.SN(net6870),
.CK(clk),
.Q(net8372),
.QN(net8371)
);

NOR2_X2 c7848(
.A1(net6454),
.A2(net8337),
.ZN(net8373)
);

DFFS_X1 c7849(
.D(net8368),
.SN(net8373),
.CK(clk),
.Q(net8375),
.QN(net8374)
);

AOI222_X1 c7850(
.A1(net8354),
.A2(net8342),
.B1(net7372),
.B2(net8294),
.C1(net8284),
.C2(net7413),
.ZN(net8376)
);

NAND3_X4 c7851(
.A1(net8370),
.A2(net5432),
.A3(net7314),
.ZN(net8377)
);

OR3_X4 c7852(
.A1(net6240),
.A2(net8109),
.A3(net8348),
.ZN(net8378)
);

XOR2_X2 c7853(
.A(net3497),
.B(net10751),
.Z(net8379)
);

XNOR2_X1 c7854(
.A(net8264),
.B(net8217),
.ZN(net8380)
);

AND3_X2 c7855(
.A1(net5458),
.A2(net8337),
.A3(net7219),
.ZN(net8381)
);

NOR3_X1 c7856(
.A1(net8374),
.A2(net8378),
.A3(net11481),
.ZN(net8382)
);

OR2_X4 c7857(
.A1(net8301),
.A2(net11181),
.ZN(net8383)
);

OR2_X1 c7858(
.A1(net8281),
.A2(net11573),
.ZN(net8384)
);

INV_X1 c7859(
.A(net9982),
.ZN(net8385)
);

XNOR2_X2 c7860(
.A(net4187),
.B(net8373),
.ZN(net8386)
);

AOI222_X4 c7861(
.A1(net8349),
.A2(net8383),
.B1(net8352),
.B2(net8329),
.C1(net8294),
.C2(net8207),
.ZN(net8387)
);

AND2_X4 c7862(
.A1(net8340),
.A2(net8353),
.ZN(net8388)
);

OR3_X2 c7863(
.A1(net8157),
.A2(net7126),
.A3(net11574),
.ZN(net8389)
);

OAI21_X2 c7864(
.A(net8362),
.B1(net8335),
.B2(net8337),
.ZN(net8390)
);

INV_X2 c7865(
.A(net10163),
.ZN(net8391)
);

AND2_X1 c7866(
.A1(net8388),
.A2(net7314),
.ZN(net8392)
);

NAND2_X1 c7867(
.A1(net8384),
.A2(net8361),
.ZN(net8393)
);

OAI21_X1 c7868(
.A(net8365),
.B1(net7329),
.B2(net6240),
.ZN(net8394)
);

SDFF_X1 c7869(
.D(net8389),
.SE(net7397),
.SI(net8377),
.CK(clk),
.Q(net8396),
.QN(net8395)
);

AOI21_X2 c7870(
.A(net8369),
.B1(net8365),
.B2(net7299),
.ZN(net8397)
);

AOI21_X1 c7871(
.A(net7342),
.B1(net7329),
.B2(net10717),
.ZN(net8398)
);

AOI21_X4 c7872(
.A(net8393),
.B1(net8335),
.B2(net8395),
.ZN(net8399)
);

SDFF_X2 c7873(
.D(net8386),
.SE(net8392),
.SI(net11573),
.CK(clk),
.Q(net8401),
.QN(net8400)
);

AND3_X1 c7874(
.A1(net7372),
.A2(net8394),
.A3(net8399),
.ZN(net8402)
);

NAND3_X1 c7875(
.A1(net8241),
.A2(net8396),
.A3(net8393),
.ZN(net8403)
);

NOR3_X4 c7876(
.A1(net8130),
.A2(net5102),
.A3(net8155),
.ZN(net8404)
);

NOR3_X2 c7877(
.A1(net7342),
.A2(net8389),
.A3(net11572),
.ZN(net8405)
);

INV_X8 c7878(
.A(net9688),
.ZN(net8406)
);

OAI221_X4 c7879(
.A(net8402),
.B1(net8403),
.B2(net8405),
.C1(net8377),
.C2(net7252),
.ZN(net8407)
);

NAND2_X2 c7880(
.A1(net8406),
.A2(net11432),
.ZN(net8408)
);

NAND2_X4 c7881(
.A1(net8394),
.A2(net8399),
.ZN(net8409)
);

AND3_X4 c7882(
.A1(net7013),
.A2(net6425),
.A3(net8396),
.ZN(net8410)
);

NAND3_X2 c7883(
.A1(net8409),
.A2(net8410),
.A3(net11432),
.ZN(net8411)
);

DFFRS_X1 c7884(
.D(net8373),
.RN(net8410),
.SN(net8411),
.CK(clk),
.Q(net8413),
.QN(net8412)
);

INV_X16 c7885(
.A(net11388),
.ZN(net8414)
);

AND2_X2 c7886(
.A1(net5515),
.A2(net6528),
.ZN(net8415)
);

INV_X32 c7887(
.A(net7252),
.ZN(net8416)
);

INV_X4 c7888(
.A(net10439),
.ZN(net8417)
);

XOR2_X1 c7889(
.A(net5102),
.B(net11262),
.Z(net8418)
);

NOR2_X1 c7890(
.A1(net8356),
.A2(net8306),
.ZN(net8419)
);

INV_X1 c7891(
.A(net9931),
.ZN(net8420)
);

OR2_X2 c7892(
.A1(net5478),
.A2(net8385),
.ZN(net8421)
);

INV_X2 c7893(
.A(net11027),
.ZN(net8422)
);

INV_X8 c7894(
.A(net11334),
.ZN(net8423)
);

INV_X16 c7895(
.A(net7363),
.ZN(net8424)
);

INV_X32 c7896(
.A(net11561),
.ZN(net8425)
);

INV_X4 c7897(
.A(net9867),
.ZN(net8426)
);

NOR2_X4 c7898(
.A1(net6481),
.A2(net8419),
.ZN(net8427)
);

INV_X1 c7899(
.A(net10089),
.ZN(net8428)
);

INV_X2 c7900(
.A(net11487),
.ZN(net8429)
);

NOR2_X2 c7901(
.A1(net8424),
.A2(net7430),
.ZN(net8430)
);

XOR2_X2 c7902(
.A(net8422),
.B(net5515),
.Z(net8431)
);

INV_X8 c7903(
.A(net11487),
.ZN(net8432)
);

XNOR2_X1 c7904(
.A(net8306),
.B(net8426),
.ZN(net8433)
);

OR2_X4 c7905(
.A1(net8420),
.A2(net7314),
.ZN(net8434)
);

INV_X16 c7906(
.A(net10492),
.ZN(net8435)
);

OR2_X1 c7907(
.A1(net7458),
.A2(net8352),
.ZN(net8436)
);

OAI22_X1 c7908(
.A1(net8414),
.A2(net8415),
.B1(net8279),
.B2(net8321),
.ZN(net8437)
);

XNOR2_X2 c7909(
.A(net8336),
.B(net8332),
.ZN(net8438)
);

AND2_X4 c7910(
.A1(net8426),
.A2(net10891),
.ZN(net8439)
);

AND2_X1 c7911(
.A1(net7451),
.A2(net8425),
.ZN(net8440)
);

NAND2_X1 c7912(
.A1(net8408),
.A2(net11006),
.ZN(net8441)
);

NAND2_X2 c7913(
.A1(net6382),
.A2(net7363),
.ZN(net8442)
);

NAND2_X4 c7914(
.A1(net7430),
.A2(net7466),
.ZN(net8443)
);

AND2_X2 c7915(
.A1(net6298),
.A2(net7314),
.ZN(net8444)
);

XOR2_X1 c7916(
.A(net8432),
.B(net5496),
.Z(net8445)
);

INV_X32 c7917(
.A(net10293),
.ZN(net8446)
);

INV_X4 c7918(
.A(net9909),
.ZN(net8447)
);

NOR2_X1 c7919(
.A1(net7219),
.A2(net8440),
.ZN(net8448)
);

OR2_X2 c7920(
.A1(net8128),
.A2(net7441),
.ZN(net8449)
);

OR3_X1 c7921(
.A1(net8435),
.A2(net8445),
.A3(net8436),
.ZN(net8450)
);

NOR2_X4 c7922(
.A1(net8423),
.A2(net8426),
.ZN(net8451)
);

NOR2_X2 c7923(
.A1(net7356),
.A2(net8398),
.ZN(net8452)
);

MUX2_X1 c7924(
.A(net8426),
.B(net8425),
.S(net2606),
.Z(net8453)
);

XOR2_X2 c7925(
.A(net8445),
.B(net8024),
.Z(net8454)
);

XNOR2_X1 c7926(
.A(net8443),
.B(net10597),
.ZN(net8455)
);

OR2_X4 c7927(
.A1(net8417),
.A2(net8444),
.ZN(net8456)
);

AND4_X2 c7928(
.A1(net7494),
.A2(net8444),
.A3(net6476),
.A4(net11561),
.ZN(net8457)
);

OR2_X1 c7929(
.A1(net7444),
.A2(net7314),
.ZN(net8458)
);

INV_X1 c7930(
.A(net8450),
.ZN(net8459)
);

XNOR2_X2 c7931(
.A(net8437),
.B(net8456),
.ZN(net8460)
);

AND2_X4 c7932(
.A1(net8442),
.A2(net8415),
.ZN(net8461)
);

AND2_X1 c7933(
.A1(net7126),
.A2(net11262),
.ZN(net8462)
);

INV_X2 c7934(
.A(net8462),
.ZN(net8463)
);

NAND2_X1 c7935(
.A1(net7915),
.A2(out13),
.ZN(net8464)
);

INV_X8 c7936(
.A(net8461),
.ZN(net8465)
);

NAND2_X2 c7937(
.A1(net8024),
.A2(net8445),
.ZN(net8466)
);

AND4_X1 c7938(
.A1(net8333),
.A2(net8443),
.A3(net8466),
.A4(net7443),
.ZN(net8467)
);

OAI21_X4 c7939(
.A(net6451),
.B1(net8465),
.B2(net8448),
.ZN(net8468)
);

NAND2_X4 c7940(
.A1(net8458),
.A2(net7314),
.ZN(net8469)
);

INV_X16 c7941(
.A(net9977),
.ZN(net8470)
);

AND2_X2 c7942(
.A1(net8347),
.A2(net8311),
.ZN(net8471)
);

DFFRS_X2 c7943(
.D(net8438),
.RN(net8452),
.SN(net8378),
.CK(clk),
.Q(net8473),
.QN(net8472)
);

XOR2_X1 c7944(
.A(net5496),
.B(net8471),
.Z(net8474)
);

NOR2_X1 c7945(
.A1(net8429),
.A2(net8454),
.ZN(net8475)
);

MUX2_X2 c7946(
.A(net5351),
.B(net8456),
.S(net8452),
.Z(net8476)
);

OR2_X2 c7947(
.A1(net6407),
.A2(net7475),
.ZN(net8477)
);

NOR2_X4 c7948(
.A1(net8425),
.A2(net8465),
.ZN(net8478)
);

NAND3_X4 c7949(
.A1(net8466),
.A2(net8448),
.A3(net8441),
.ZN(net8479)
);

NOR2_X2 c7950(
.A1(net8449),
.A2(net8286),
.ZN(net8480)
);

XOR2_X2 c7951(
.A(net8454),
.B(net7444),
.Z(net8481)
);

SDFFS_X1 c7952(
.D(net8465),
.SE(net8478),
.SI(net8469),
.SN(net7451),
.CK(clk),
.Q(net8483),
.QN(net8482)
);

OR3_X4 c7953(
.A1(net8451),
.A2(net8464),
.A3(net8428),
.ZN(net8484)
);

AND3_X2 c7954(
.A1(net8479),
.A2(net8484),
.A3(net8482),
.ZN(net8485)
);

INV_X32 c7955(
.A(net11430),
.ZN(net8486)
);

NOR3_X1 c7956(
.A1(net8483),
.A2(net8446),
.A3(net8479),
.ZN(net8487)
);

AOI22_X4 c7957(
.A1(net8366),
.A2(net8480),
.B1(net8485),
.B2(net7445),
.ZN(net8488)
);

OR3_X2 c7958(
.A1(net7465),
.A2(net8464),
.A3(net8483),
.ZN(net8489)
);

SDFF_X1 c7959(
.D(net8459),
.SE(net6418),
.SI(net8484),
.CK(clk),
.Q(net8491),
.QN(net8490)
);

SDFF_X2 c7960(
.D(net2606),
.SE(net8491),
.SI(net8207),
.CK(clk),
.Q(net8493),
.QN(net8492)
);

OAI21_X2 c7961(
.A(net8474),
.B1(net8493),
.B2(net8490),
.ZN(net8494)
);

OAI21_X1 c7962(
.A(net7357),
.B1(net8486),
.B2(net8492),
.ZN(net8495)
);

OAI33_X1 c7963(
.A1(net8463),
.A2(net8482),
.A3(net8345),
.B1(net5545),
.B2(net6450),
.B3(net11065),
.ZN(net8496)
);

SDFFRS_X2 c7964(
.D(net8419),
.RN(net8487),
.SE(net8478),
.SI(net7356),
.SN(net11576),
.CK(clk),
.Q(net8498),
.QN(net8497)
);

OAI22_X4 c7965(
.A1(net8455),
.A2(net8449),
.B1(net8490),
.B2(net11576),
.ZN(net8499)
);

AOI22_X2 c7966(
.A1(net8485),
.A2(net8447),
.B1(net10716),
.B2(net11576),
.ZN(net8500)
);

AOI21_X2 c7967(
.A(net8484),
.B1(net10940),
.B2(net11240),
.ZN(net8501)
);

INV_X4 c7968(
.A(net11374),
.ZN(net8502)
);

NAND4_X4 c7969(
.A1(net6541),
.A2(net8345),
.A3(net7588),
.A4(net7559),
.ZN(net8503)
);

AOI21_X1 c7970(
.A(net6333),
.B1(net7535),
.B2(net8415),
.ZN(net8504)
);

INV_X1 c7971(
.A(net11428),
.ZN(net8505)
);

XNOR2_X1 c7972(
.A(net8352),
.B(net6423),
.ZN(net8506)
);

OR2_X4 c7973(
.A1(net7606),
.A2(net7563),
.ZN(net8507)
);

OR2_X1 c7974(
.A1(net8364),
.A2(net8506),
.ZN(net8508)
);

XNOR2_X2 c7975(
.A(net7589),
.B(net11577),
.ZN(net8509)
);

AOI21_X4 c7976(
.A(net8481),
.B1(net8508),
.B2(net7441),
.ZN(net8510)
);

AND2_X4 c7977(
.A1(net8505),
.A2(net8430),
.ZN(net8511)
);

AND3_X1 c7978(
.A1(net5616),
.A2(net6558),
.A3(net7455),
.ZN(net8512)
);

AND2_X1 c7979(
.A1(net7466),
.A2(net8412),
.ZN(net8513)
);

NAND2_X1 c7980(
.A1(net8447),
.A2(net8471),
.ZN(net8514)
);

NAND3_X1 c7981(
.A1(net8441),
.A2(net8408),
.A3(net7597),
.ZN(net8515)
);

NOR3_X4 c7982(
.A1(net7600),
.A2(net8508),
.A3(net7414),
.ZN(net8516)
);

INV_X2 c7983(
.A(net10032),
.ZN(net8517)
);

INV_X8 c7984(
.A(net10046),
.ZN(net8518)
);

DFFRS_X1 c7985(
.D(net7590),
.RN(net8507),
.SN(net8506),
.CK(clk),
.Q(net8520),
.QN(net8519)
);

NAND2_X2 c7986(
.A1(net7530),
.A2(net8508),
.ZN(net8521)
);

NAND2_X4 c7987(
.A1(net8516),
.A2(net10571),
.ZN(net8522)
);

NOR3_X2 c7988(
.A1(net8513),
.A2(net8472),
.A3(net7561),
.ZN(net8523)
);

AND3_X4 c7989(
.A1(net1732),
.A2(net8521),
.A3(net11573),
.ZN(net8524)
);

NAND3_X2 c7990(
.A1(net8501),
.A2(net5623),
.A3(net11575),
.ZN(net8525)
);

INV_X16 c7991(
.A(net9932),
.ZN(net8526)
);

INV_X32 c7992(
.A(net9868),
.ZN(net8527)
);

AND2_X2 c7993(
.A1(net8439),
.A2(net8506),
.ZN(net8528)
);

OR3_X1 c7994(
.A1(net6423),
.A2(net8510),
.A3(net8519),
.ZN(net8529)
);

INV_X4 c7995(
.A(net10030),
.ZN(net8530)
);

DFFRS_X2 c7996(
.D(net7571),
.RN(net8529),
.SN(net8522),
.CK(clk),
.Q(net8532),
.QN(net8531)
);

XOR2_X1 c7997(
.A(net6553),
.B(net8322),
.Z(net8533)
);

NOR2_X1 c7998(
.A1(net7455),
.A2(net8528),
.ZN(net8534)
);

SDFF_X1 c7999(
.D(net8526),
.SE(net8523),
.SI(net8528),
.CK(clk),
.Q(net8536),
.QN(net8535)
);

INV_X1 c8000(
.A(net9808),
.ZN(net8537)
);

MUX2_X1 c8001(
.A(net7543),
.B(net8533),
.S(net7517),
.Z(net8538)
);

OR2_X2 c8002(
.A1(net6397),
.A2(net8518),
.ZN(net8539)
);

NOR2_X4 c8003(
.A1(net7514),
.A2(net8517),
.ZN(net8540)
);

OAI21_X4 c8004(
.A(net8530),
.B1(net6423),
.B2(net7546),
.ZN(net8541)
);

MUX2_X2 c8005(
.A(net7521),
.B(net6600),
.S(net8415),
.Z(net8542)
);

NOR2_X2 c8006(
.A1(net7127),
.A2(net7535),
.ZN(net8543)
);

SDFF_X2 c8007(
.D(net7517),
.SE(net8533),
.SI(net8478),
.CK(clk),
.Q(net8545),
.QN(net8544)
);

NAND3_X4 c8008(
.A1(net4392),
.A2(net8518),
.A3(net7414),
.ZN(net8546)
);

XOR2_X2 c8009(
.A(net8512),
.B(net7541),
.Z(net8547)
);

OR3_X4 c8010(
.A1(net8541),
.A2(net8415),
.A3(net8542),
.ZN(net8548)
);

OAI211_X2 c8011(
.A(net8537),
.B(net4604),
.C1(net8535),
.C2(net11572),
.ZN(net8549)
);

INV_X2 c8012(
.A(net11464),
.ZN(net8550)
);

XNOR2_X1 c8013(
.A(net8543),
.B(net8545),
.ZN(net8551)
);

OR2_X4 c8014(
.A1(net8551),
.A2(net8441),
.ZN(net8552)
);

AND3_X2 c8015(
.A1(net8539),
.A2(net8528),
.A3(net8542),
.ZN(net8553)
);

OR4_X2 c8016(
.A1(net8501),
.A2(net8552),
.A3(net8542),
.A4(net8517),
.ZN(net8554)
);

NOR3_X1 c8017(
.A1(net4604),
.A2(net8531),
.A3(net2713),
.ZN(net8555)
);

SDFFRS_X1 c8018(
.D(net8428),
.RN(net7915),
.SE(net8553),
.SI(net8528),
.SN(net8377),
.CK(clk),
.Q(net8557),
.QN(net8556)
);

OR3_X2 c8019(
.A1(net8375),
.A2(net8555),
.A3(net8544),
.ZN(net8558)
);

AOI211_X1 c8020(
.A(net8520),
.B(net6423),
.C1(net5545),
.C2(net10598),
.ZN(net8559)
);

OAI21_X2 c8021(
.A(net8380),
.B1(net8550),
.B2(net8553),
.ZN(net8560)
);

OAI21_X1 c8022(
.A(net8286),
.B1(net8557),
.B2(net7449),
.ZN(net8561)
);

DFFRS_X1 c8023(
.D(net8478),
.RN(net8552),
.SN(net7588),
.CK(clk),
.Q(net8563),
.QN(net8562)
);

OAI221_X2 c8024(
.A(net8548),
.B1(net8478),
.B2(net8492),
.C1(net11186),
.C2(net11562),
.ZN(net8564)
);

AOI21_X2 c8025(
.A(net6550),
.B1(net7441),
.B2(net11154),
.ZN(net8565)
);

DFFRS_X2 c8026(
.D(net8540),
.RN(net8555),
.SN(net7812),
.CK(clk),
.Q(net8567),
.QN(net8566)
);

AOI21_X1 c8027(
.A(net7442),
.B1(net6550),
.B2(net8562),
.ZN(net8568)
);

AOI21_X4 c8028(
.A(net8567),
.B1(net8528),
.B2(net8549),
.ZN(net8569)
);

AOI221_X4 c8029(
.A(net5621),
.B1(net8377),
.B2(net8556),
.C1(net8012),
.C2(net8353),
.ZN(net8570)
);

AND3_X1 c8030(
.A1(net7441),
.A2(net8563),
.A3(net11253),
.ZN(net8571)
);

OR2_X1 c8031(
.A1(net8550),
.A2(net8364),
.ZN(net8572)
);

NAND3_X1 c8032(
.A1(net8563),
.A2(net4598),
.A3(net10721),
.ZN(net8573)
);

NOR3_X4 c8033(
.A1(net6600),
.A2(net8522),
.A3(net5383),
.ZN(net8574)
);

NOR3_X2 c8034(
.A1(net8571),
.A2(net8377),
.A3(net8569),
.ZN(net8575)
);

SDFF_X1 c8035(
.D(net8436),
.SE(net7580),
.SI(net8207),
.CK(clk),
.Q(net8577),
.QN(net8576)
);

AND3_X4 c8036(
.A1(net8560),
.A2(net8514),
.A3(net8528),
.ZN(net8578)
);

NAND4_X2 c8037(
.A1(net8532),
.A2(net8546),
.A3(net3615),
.A4(net8556),
.ZN(net8579)
);

INV_X8 c8038(
.A(net11428),
.ZN(net8580)
);

NAND3_X2 c8039(
.A1(net8536),
.A2(net8412),
.A3(net10557),
.ZN(net8581)
);

XNOR2_X2 c8040(
.A(net11091),
.B(net11187),
.ZN(net8582)
);

SDFF_X2 c8041(
.D(net8502),
.SE(net8579),
.SI(net8477),
.CK(clk),
.Q(net8584),
.QN(net8583)
);

AND2_X4 c8042(
.A1(net8527),
.A2(net10556),
.ZN(net8585)
);

OR3_X1 c8043(
.A1(net8572),
.A2(net8580),
.A3(net8581),
.ZN(net8586)
);

MUX2_X1 c8044(
.A(net8586),
.B(net8581),
.S(net8540),
.Z(net8587)
);

OAI21_X4 c8045(
.A(net8582),
.B1(net8517),
.B2(net10939),
.ZN(net8588)
);

MUX2_X2 c8046(
.A(net8565),
.B(net8582),
.S(net11202),
.Z(net8589)
);

NAND3_X4 c8047(
.A1(net7449),
.A2(net8588),
.A3(net8587),
.ZN(net8590)
);

OR3_X4 c8048(
.A1(net8583),
.A2(net10772),
.A3(net11147),
.ZN(net8591)
);

DFFRS_X1 c8049(
.D(net7587),
.RN(net8585),
.SN(net8566),
.CK(clk),
.Q(net8593),
.QN(net8592)
);

AOI222_X2 c8050(
.A1(net8584),
.A2(net8591),
.B1(net8593),
.B2(net8556),
.C1(net8353),
.C2(net8519),
.ZN(net8594)
);

AND2_X1 c8051(
.A1(net8398),
.A2(net8553),
.ZN(net8595)
);

NAND2_X1 c8052(
.A1(net8495),
.A2(net2751),
.ZN(net8596)
);

NAND2_X2 c8053(
.A1(net3627),
.A2(out25),
.ZN(net8597)
);

AND3_X2 c8054(
.A1(net840),
.A2(net8491),
.A3(net7359),
.ZN(net8598)
);

DFFRS_X2 c8055(
.D(net8378),
.RN(net8329),
.SN(net5383),
.CK(clk),
.Q(net8600),
.QN(net8599)
);

NAND2_X4 c8056(
.A1(net5685),
.A2(net7627),
.ZN(net8601)
);

NOR3_X1 c8057(
.A1(net8345),
.A2(net4753),
.A3(net6689),
.ZN(net8602)
);

SDFF_X1 c8058(
.D(net8521),
.SE(net7674),
.SI(net5482),
.CK(clk),
.Q(net8604),
.QN(net8603)
);

OR3_X2 c8059(
.A1(net7627),
.A2(net6682),
.A3(net7673),
.ZN(net8605)
);

OAI21_X2 c8060(
.A(net8605),
.B1(net8557),
.B2(net2606),
.ZN(net8606)
);

AOI221_X2 c8061(
.A(net7559),
.B1(net8603),
.B2(net7627),
.C1(net6507),
.C2(net7577),
.ZN(net8607)
);

SDFF_X2 c8062(
.D(net8311),
.SE(net7359),
.SI(net8493),
.CK(clk),
.Q(net8609),
.QN(net8608)
);

AND2_X2 c8063(
.A1(net5449),
.A2(net1730),
.ZN(net8610)
);

OAI21_X1 c8064(
.A(net7664),
.B1(net7559),
.B2(net7640),
.ZN(net8611)
);

AOI21_X2 c8065(
.A(net3742),
.B1(out25),
.B2(net3452),
.ZN(net8612)
);

XOR2_X1 c8066(
.A(net8473),
.B(net8549),
.Z(net8613)
);

AOI21_X1 c8067(
.A(net8607),
.B1(net5704),
.B2(net11577),
.ZN(net8614)
);

INV_X16 c8068(
.A(net11374),
.ZN(net8615)
);

DFFRS_X1 c8069(
.D(net7688),
.RN(net8599),
.SN(net8610),
.CK(clk),
.Q(net8617),
.QN(net8616)
);

DFFRS_X2 c8070(
.D(net7560),
.RN(net7690),
.SN(net7693),
.CK(clk),
.Q(net8619),
.QN(net8618)
);

AOI21_X4 c8071(
.A(net6689),
.B1(net8590),
.B2(net7673),
.ZN(net8620)
);

AOI221_X1 c8072(
.A(net7695),
.B1(net8521),
.B2(net8573),
.C1(net8329),
.C2(net8608),
.ZN(net8621)
);

SDFF_X1 c8073(
.D(net7541),
.SE(net8517),
.SI(net8514),
.CK(clk),
.Q(net8623),
.QN(net8622)
);

OR4_X4 c8074(
.A1(net6679),
.A2(net4539),
.A3(net7359),
.A4(net8608),
.ZN(net8624)
);

AND3_X1 c8075(
.A1(net3750),
.A2(net8616),
.A3(net8619),
.ZN(net8625)
);

NAND3_X1 c8076(
.A1(net8605),
.A2(net5449),
.A3(net11236),
.ZN(net8626)
);

SDFF_X2 c8077(
.D(net5482),
.SE(net5704),
.SI(net3742),
.CK(clk),
.Q(net8628),
.QN(net8627)
);

NOR3_X4 c8078(
.A1(net8470),
.A2(net8521),
.A3(net3750),
.ZN(net8629)
);

NOR2_X1 c8079(
.A1(net7692),
.A2(net8279),
.ZN(net8630)
);

NOR3_X2 c8080(
.A1(net7448),
.A2(net8604),
.A3(net8628),
.ZN(net8631)
);

AND3_X4 c8081(
.A1(net8484),
.A2(net7211),
.A3(net10856),
.ZN(net8632)
);

NAND3_X2 c8082(
.A1(net7640),
.A2(net8610),
.A3(net8573),
.ZN(net8633)
);

OR3_X1 c8083(
.A1(net7673),
.A2(net8568),
.A3(net8484),
.ZN(net8634)
);

MUX2_X1 c8084(
.A(net8517),
.B(net8619),
.S(net8623),
.Z(net8635)
);

OR2_X2 c8085(
.A1(net7661),
.A2(net11443),
.ZN(net8636)
);

OAI21_X4 c8086(
.A(net6558),
.B1(net8493),
.B2(net6559),
.ZN(net8637)
);

MUX2_X2 c8087(
.A(net6507),
.B(net8636),
.S(net8619),
.Z(net8638)
);

INV_X32 c8088(
.A(net9727),
.ZN(net8639)
);

NAND3_X4 c8089(
.A1(net8638),
.A2(net8636),
.A3(net8569),
.ZN(net8640)
);

OR3_X4 c8090(
.A1(net8596),
.A2(net7540),
.A3(net8635),
.ZN(net8641)
);

INV_X4 c8091(
.A(net9835),
.ZN(net8642)
);

OAI222_X1 c8092(
.A1(net5685),
.A2(net7577),
.B1(net8610),
.B2(net8618),
.C1(net11082),
.C2(net11266),
.ZN(net8643)
);

AND3_X2 c8093(
.A1(net6716),
.A2(net8617),
.A3(net2777),
.ZN(net8644)
);

NOR3_X1 c8094(
.A1(net8332),
.A2(net8609),
.A3(net8596),
.ZN(net8645)
);

OR3_X2 c8095(
.A1(net8497),
.A2(net8596),
.A3(net10712),
.ZN(net8646)
);

OAI21_X2 c8096(
.A(net4592),
.B1(net3750),
.B2(net8608),
.ZN(net8647)
);

DFFRS_X1 c8097(
.D(net8639),
.RN(net7693),
.SN(net10963),
.CK(clk),
.Q(net8649),
.QN(net8648)
);

OAI21_X1 c8098(
.A(net8609),
.B1(net6679),
.B2(net8618),
.ZN(net8650)
);

AOI21_X2 c8099(
.A(net4753),
.B1(net8613),
.B2(net8635),
.ZN(net8651)
);

AOI21_X1 c8100(
.A(net6668),
.B1(net6715),
.B2(net10809),
.ZN(net8652)
);

AOI21_X4 c8101(
.A(net8555),
.B1(net8632),
.B2(net8647),
.ZN(net8653)
);

AND3_X1 c8102(
.A1(net7628),
.A2(net8642),
.A3(net8623),
.ZN(net8654)
);

OAI221_X1 c8103(
.A(net6682),
.B1(net8642),
.B2(net8596),
.C1(net7674),
.C2(net6548),
.ZN(net8655)
);

NAND3_X1 c8104(
.A1(net6548),
.A2(net8649),
.A3(net8596),
.ZN(net8656)
);

NOR3_X4 c8105(
.A1(net6559),
.A2(net8630),
.A3(net8647),
.ZN(net8657)
);

OAI22_X2 c8106(
.A1(net8608),
.A2(net8627),
.B1(net11204),
.B2(net11211),
.ZN(net8658)
);

NOR3_X2 c8107(
.A1(net8658),
.A2(net8651),
.A3(net8647),
.ZN(net8659)
);

NOR2_X4 c8108(
.A1(net8652),
.A2(net8659),
.ZN(net8660)
);

AND3_X4 c8109(
.A1(net8329),
.A2(net8619),
.A3(net6715),
.ZN(net8661)
);

NAND3_X2 c8110(
.A1(net8647),
.A2(net8635),
.A3(net8612),
.ZN(net8662)
);

OR3_X1 c8111(
.A1(net7674),
.A2(net8655),
.A3(net8661),
.ZN(net8663)
);

OAI211_X4 c8112(
.A(net6682),
.B(net8609),
.C1(net10808),
.C2(net11443),
.ZN(net8664)
);

MUX2_X1 c8113(
.A(net8569),
.B(net8663),
.S(net8609),
.Z(net8665)
);

OAI21_X4 c8114(
.A(net8553),
.B1(net8662),
.B2(net8660),
.ZN(net8666)
);

NOR2_X2 c8115(
.A1(net8661),
.A2(net10914),
.ZN(net8667)
);

MUX2_X2 c8116(
.A(net8408),
.B(net8636),
.S(net8647),
.Z(net8668)
);

XOR2_X2 c8117(
.A(net8668),
.B(net8640),
.Z(net8669)
);

NAND3_X4 c8118(
.A1(net8346),
.A2(net8669),
.A3(net8491),
.ZN(net8670)
);

OR3_X4 c8119(
.A1(net8656),
.A2(net8547),
.A3(net8648),
.ZN(net8671)
);

DFFRS_X2 c8120(
.D(net7475),
.RN(net8557),
.SN(net8666),
.CK(clk),
.Q(net8673),
.QN(net8672)
);

AND3_X2 c8121(
.A1(net8650),
.A2(net8577),
.A3(net10941),
.ZN(net8674)
);

NOR3_X1 c8122(
.A1(net8660),
.A2(net8596),
.A3(net10713),
.ZN(net8675)
);

OR3_X2 c8123(
.A1(net8514),
.A2(net8645),
.A3(net8644),
.ZN(net8676)
);

SDFF_X1 c8124(
.D(net7667),
.SE(net7693),
.SI(net11448),
.CK(clk),
.Q(net8678),
.QN(net8677)
);

OAI21_X2 c8125(
.A(net8654),
.B1(net8674),
.B2(net8650),
.ZN(net8679)
);

OAI21_X1 c8126(
.A(net8679),
.B1(net6715),
.B2(net3742),
.ZN(net8680)
);

INV_X1 c8127(
.A(net9726),
.ZN(net8681)
);

AOI21_X2 c8128(
.A(net7673),
.B1(net10723),
.B2(net10855),
.ZN(net8682)
);

AOI21_X1 c8129(
.A(net7512),
.B1(net8644),
.B2(net8682),
.ZN(net8683)
);

AOI21_X4 c8130(
.A(net8664),
.B1(net7693),
.B2(net8671),
.ZN(net8684)
);

AND3_X1 c8131(
.A1(net8631),
.A2(net8680),
.A3(net8647),
.ZN(net8685)
);

NAND3_X1 c8132(
.A1(net8549),
.A2(net8628),
.A3(net11259),
.ZN(net8686)
);

NOR3_X4 c8133(
.A1(net8685),
.A2(net8610),
.A3(net11141),
.ZN(net8687)
);

OAI211_X1 c8160(
.A(net6772),
.B(net4792),
.C1(out3),
.C2(net5791),
.ZN(net8688)
);

SDFF_X2 c8161(
.D(net8610),
.SE(net8413),
.SI(net8728),
.CK(clk),
.Q(net8690),
.QN(net8689)
);

NOR4_X4 c8162(
.A1(net7778),
.A2(net8678),
.A3(net6779),
.A4(net8733),
.ZN(net8691)
);

NOR3_X2 c8163(
.A1(net7546),
.A2(net8690),
.A3(net8730),
.ZN(net8692)
);

INV_X2 c8164(
.A(net11589),
.ZN(out6)
);

NOR4_X2 c8165(
.A1(net6607),
.A2(net6801),
.A3(net5795),
.A4(net8610),
.ZN(net8693)
);

AOI211_X4 c8166(
.A(net7720),
.B(net7787),
.C1(net8721),
.C2(net11282),
.ZN(net8694)
);

NOR4_X1 c8167(
.A1(net7754),
.A2(net7633),
.A3(net8730),
.A4(net10514),
.ZN(net8695)
);

AND3_X4 c8168(
.A1(net8690),
.A2(net8721),
.A3(net11294),
.ZN(net8696)
);

NAND3_X2 c8169(
.A1(net8694),
.A2(net8696),
.A3(net8641),
.ZN(net8697)
);

OR3_X1 c8170(
.A1(net5795),
.A2(net7770),
.A3(net8721),
.ZN(net8698)
);

MUX2_X1 c8171(
.A(net8568),
.B(net8696),
.S(net8734),
.Z(net8699)
);

SDFFS_X2 c8172(
.D(net8729),
.SE(net8727),
.SI(net6800),
.SN(net8736),
.CK(clk),
.Q(net8701),
.QN(net8700)
);

OAI21_X4 c8173(
.A(net8577),
.B1(net8678),
.B2(net7787),
.ZN(net8702)
);

MUX2_X2 c8174(
.A(net5742),
.B(net7582),
.S(net8736),
.Z(net8703)
);

NAND3_X4 c8175(
.A1(net5580),
.A2(net7582),
.A3(net8723),
.ZN(out20)
);

OAI221_X4 c8176(
.A(net8698),
.B1(net8734),
.B2(net8689),
.C1(net8721),
.C2(net8610),
.ZN(net8704)
);

OR3_X4 c8177(
.A1(net6643),
.A2(net8736),
.A3(net5815),
.ZN(net8705)
);

AND3_X2 c8178(
.A1(net8573),
.A2(net8741),
.A3(net8688),
.ZN(net8706)
);

NOR3_X1 c8179(
.A1(net8720),
.A2(net8700),
.A3(net11281),
.ZN(out21)
);

OR3_X2 c8180(
.A1(net8737),
.A2(net7727),
.A3(net8738),
.ZN(net8707)
);

OAI21_X2 c8181(
.A(net8721),
.B1(net8692),
.B2(net8690),
.ZN(net8708)
);

OAI21_X1 c8182(
.A(net8688),
.B1(net8701),
.B2(net7546),
.ZN(out11)
);

AOI21_X2 c8183(
.A(net2894),
.B1(net7766),
.B2(net10998),
.ZN(net8709)
);

DFFRS_X1 c8184(
.D(net8590),
.RN(net8706),
.SN(net11293),
.CK(clk),
.Q(out17),
.QN(net8710)
);

OAI221_X2 c8185(
.A(net8726),
.B1(net7739),
.B2(net8576),
.C1(net6803),
.ZN(net11304)
);

OAI222_X4 c8186(
.A1(net8728),
.A2(net8691),
.B1(net8689),
.B2(net8710),
.C1(out25),
.C2(net7633),
.ZN(net8712)
);

AOI211_X2 c8187(
.A(net8702),
.B(out17),
.C1(out1),
.C2(net11273),
.ZN(net8713)
);

AOI221_X4 c8188(
.A(net4791),
.B1(net8710),
.B2(net8736),
.C1(net11083),
.C2(net11156),
.ZN(net8714)
);

OAI222_X2 c8189(
.A1(net6779),
.A2(net8707),
.B1(net8736),
.B2(out17),
.C1(net5704),
.C2(net8673),
.ZN(net8715)
);

AOI222_X1 c8190(
.A1(net7686),
.A2(net8695),
.B1(net8733),
.B2(net7770),
.C1(net8721),
.C2(net11319),
.ZN(net8716)
);

AOI21_X1 c8191(
.A(net8730),
.B1(net5792),
.B2(net10513),
.ZN(out18)
);

AOI21_X4 c8192(
.A(out18),
.B1(net11161),
.B2(net11387),
.ZN(net8717)
);

AND3_X1 c8193(
.A1(net6732),
.A2(net7782),
.A3(net5704),
.ZN(net8718)
);

DFFRS_X2 c8194(
.D(net7732),
.RN(net7787),
.SN(out16),
.CK(clk),
.Q(net8720),
.QN(net8719)
);

NAND3_X1 c8195(
.A1(net4792),
.A2(net7754),
.A3(net8587),
.ZN(out24)
);

NOR3_X4 c8196(
.A1(net7676),
.A2(net7713),
.A3(net8719),
.ZN(net8721)
);

NOR3_X2 c8197(
.A1(net7633),
.A2(net8641),
.A3(net5792),
.ZN(net8722)
);

SDFF_X1 c8198(
.D(net7700),
.SE(net5704),
.SI(net2894),
.CK(clk),
.Q(net8724),
.QN(net8723)
);

AND3_X4 c8199(
.A1(net6728),
.A2(out9),
.A3(net6643),
.ZN(net8725)
);

NAND3_X2 c8200(
.A1(net8725),
.A2(net4853),
.A3(net8576),
.ZN(net8726)
);

AOI22_X1 c8201(
.A1(net7755),
.A2(net8724),
.B1(net8641),
.B2(out9),
.ZN(net8727)
);

OR3_X1 c8202(
.A1(net7727),
.A2(net8722),
.A3(net8721),
.ZN(net8728)
);

MUX2_X1 c8203(
.A(net7670),
.B(net7720),
.S(net5704),
.Z(net8729)
);

OAI21_X4 c8204(
.A(net5815),
.B1(net6772),
.B2(net7633),
.ZN(net8730)
);

AND4_X4 c8205(
.A1(net6766),
.A2(net6643),
.A3(net8730),
.A4(net11001),
.ZN(out22)
);

MUX2_X2 c8206(
.A(net2892),
.B(net6803),
.S(net7787),
.Z(net8731)
);

NAND4_X1 c8207(
.A1(net8597),
.A2(net7766),
.A3(net7770),
.A4(net6643),
.ZN(net8732)
);

SDFF_X2 c8208(
.D(net7784),
.SE(net7641),
.SI(net7781),
.CK(clk),
.Q(net8734),
.QN(net8733)
);

NAND3_X4 c8209(
.A1(net6734),
.A2(net6607),
.A3(net8677),
.ZN(out14)
);

OR3_X4 c8210(
.A1(net8587),
.A2(net8610),
.A3(net4791),
.ZN(net8735)
);

AND3_X2 c8211(
.A1(net7779),
.A2(net8730),
.A3(net7720),
.ZN(net8736)
);

NOR3_X1 c8212(
.A1(net5792),
.A2(net4853),
.A3(net10936),
.ZN(net8737)
);

DFFRS_X1 c8213(
.D(net8732),
.RN(net8734),
.SN(net7582),
.CK(clk),
.Q(net8739),
.QN(net8738)
);

OR3_X2 c8214(
.A1(net7739),
.A2(net8739),
.A3(net8736),
.ZN(net8740)
);

OAI21_X2 c8215(
.A(net8413),
.B1(net7676),
.B2(net11230),
.ZN(out12)
);

INV_X8 c8216(
.A(net11588),
.ZN(net8741)
);

INV_X16 c8217(
.A(net7875),
.ZN(net8742)
);

INV_X32 c8218(
.A(net9775),
.ZN(net8743)
);

XNOR2_X1 c8219(
.A(net4862),
.B(net7836),
.ZN(net8744)
);

INV_X4 c8220(
.A(net8742),
.ZN(net8745)
);

INV_X1 c8221(
.A(net7851),
.ZN(net8746)
);

INV_X2 c8222(
.A(net8743),
.ZN(net8747)
);

INV_X8 c8223(
.A(net6899),
.ZN(net8748)
);

INV_X16 c8224(
.A(net7875),
.ZN(net8749)
);

OR2_X4 c8225(
.A1(net5894),
.A2(net6873),
.ZN(net8750)
);

INV_X32 c8226(
.A(net6838),
.ZN(net8751)
);

INV_X4 c8227(
.A(net7847),
.ZN(net8752)
);

INV_X1 c8228(
.A(net8743),
.ZN(net8753)
);

OAI21_X1 c8229(
.A(net4929),
.B1(net8749),
.B2(net7800),
.ZN(net8754)
);

OR2_X1 c8230(
.A1(net6883),
.A2(net7875),
.ZN(net8755)
);

INV_X2 c8231(
.A(net5913),
.ZN(net8756)
);

INV_X8 c8232(
.A(net8756),
.ZN(net8757)
);

INV_X16 c8233(
.A(net8749),
.ZN(net8758)
);

INV_X32 c8234(
.A(net9774),
.ZN(net8759)
);

INV_X4 c8235(
.A(net7829),
.ZN(net8760)
);

INV_X1 c8236(
.A(net8749),
.ZN(net8761)
);

INV_X2 c8237(
.A(net8747),
.ZN(net8762)
);

INV_X8 c8238(
.A(net7836),
.ZN(net8763)
);

INV_X16 c8239(
.A(net7885),
.ZN(net8764)
);

XNOR2_X2 c8240(
.A(net8751),
.B(net7820),
.ZN(net8765)
);

AND2_X4 c8241(
.A1(net8756),
.A2(net8765),
.ZN(net8766)
);

INV_X32 c8242(
.A(net8766),
.ZN(net8767)
);

INV_X4 c8243(
.A(net8765),
.ZN(net8768)
);

INV_X1 c8244(
.A(net8746),
.ZN(net8769)
);

INV_X2 c8245(
.A(net7853),
.ZN(net8770)
);

DFFS_X2 c8246(
.D(net5883),
.SN(net8754),
.CK(clk),
.Q(net8772),
.QN(net8771)
);

INV_X8 c8247(
.A(net5839),
.ZN(net8773)
);

INV_X16 c8248(
.A(net8758),
.ZN(net8774)
);

INV_X32 c8249(
.A(net6893),
.ZN(net8775)
);

INV_X4 c8250(
.A(net8745),
.ZN(net8776)
);

INV_X1 c8251(
.A(net7828),
.ZN(net8777)
);

INV_X2 c8252(
.A(net9840),
.ZN(net8778)
);

INV_X8 c8253(
.A(net8771),
.ZN(net8779)
);

INV_X16 c8254(
.A(net8768),
.ZN(net8780)
);

INV_X32 c8255(
.A(net8778),
.ZN(net8781)
);

AND2_X1 c8256(
.A1(net8777),
.A2(net8764),
.ZN(net8782)
);

NAND2_X1 c8257(
.A1(net8776),
.A2(net8765),
.ZN(net8783)
);

NAND2_X2 c8258(
.A1(net8770),
.A2(net8750),
.ZN(net8784)
);

NAND2_X4 c8259(
.A1(net8758),
.A2(net8781),
.ZN(net8785)
);

AND2_X2 c8260(
.A1(net8783),
.A2(net8752),
.ZN(net8786)
);

INV_X4 c8261(
.A(net8782),
.ZN(net8787)
);

XOR2_X1 c8262(
.A(net7845),
.B(net8770),
.Z(net8788)
);

INV_X1 c8263(
.A(net7877),
.ZN(net8789)
);

NOR2_X1 c8264(
.A1(net8774),
.A2(net7875),
.ZN(net8790)
);

INV_X2 c8265(
.A(net8781),
.ZN(net8791)
);

OR2_X2 c8266(
.A1(net8759),
.A2(net8788),
.ZN(net8792)
);

INV_X8 c8267(
.A(net8791),
.ZN(net8793)
);

NOR2_X4 c8268(
.A1(net8774),
.A2(net8753),
.ZN(net8794)
);

NOR2_X2 c8269(
.A1(net8794),
.A2(net8781),
.ZN(net8795)
);

INV_X16 c8270(
.A(net8762),
.ZN(net8796)
);

XOR2_X2 c8271(
.A(net8786),
.B(net8782),
.Z(net8797)
);

XNOR2_X1 c8272(
.A(net8767),
.B(net8797),
.ZN(net8798)
);

OR2_X4 c8273(
.A1(net6873),
.A2(net8787),
.ZN(net8799)
);

AOI21_X2 c8274(
.A(net8760),
.B1(net8778),
.B2(net8787),
.ZN(net8800)
);

OR2_X1 c8275(
.A1(net8744),
.A2(net8797),
.ZN(net8801)
);

XNOR2_X2 c8276(
.A(net8764),
.B(net8750),
.ZN(net8802)
);

AND2_X4 c8277(
.A1(net8788),
.A2(net8778),
.ZN(net8803)
);

AND2_X1 c8278(
.A1(net8803),
.A2(net8792),
.ZN(net8804)
);

NAND2_X1 c8279(
.A1(net8779),
.A2(net6873),
.ZN(net8805)
);

NAND2_X2 c8280(
.A1(net8783),
.A2(net8791),
.ZN(net8806)
);

NAND2_X4 c8281(
.A1(net8804),
.A2(net8805),
.ZN(net8807)
);

OR4_X1 c8282(
.A1(net8795),
.A2(net8803),
.A3(net8805),
.A4(net8769),
.ZN(net8808)
);

AND2_X2 c8283(
.A1(net8755),
.A2(net8807),
.ZN(net8809)
);

OAI22_X1 c8284(
.A1(net8809),
.A2(net8807),
.B1(net7877),
.B2(net8805),
.ZN(net8810)
);

SDFFR_X1 c8285(
.D(net8798),
.RN(net7853),
.SE(net7816),
.SI(net8787),
.CK(clk),
.Q(net8812),
.QN(net8811)
);

AOI21_X1 c8286(
.A(net8775),
.B1(net8811),
.B2(net5898),
.ZN(net8813)
);

AOI21_X4 c8287(
.A(net8806),
.B1(net8800),
.B2(net8792),
.ZN(net8814)
);

DFFRS_X2 c8288(
.D(net8772),
.RN(net8807),
.SN(net8808),
.CK(clk),
.Q(net8816),
.QN(net8815)
);

SDFF_X1 c8289(
.D(net8799),
.SE(net8798),
.SI(net8807),
.CK(clk),
.Q(net8818),
.QN(net8817)
);

XOR2_X1 c8290(
.A(net7847),
.B(net8809),
.Z(net8819)
);

NOR2_X1 c8291(
.A1(net7829),
.A2(net8803),
.ZN(net8820)
);

AND4_X2 c8292(
.A1(net8796),
.A2(net8815),
.A3(net8801),
.A4(net8814),
.ZN(net8821)
);

AND4_X1 c8293(
.A1(net8790),
.A2(net8779),
.A3(net8744),
.A4(net8787),
.ZN(net8822)
);

OR2_X2 c8294(
.A1(net8822),
.A2(net8820),
.ZN(net8823)
);

AND3_X1 c8295(
.A1(net8761),
.A2(net8753),
.A3(net8814),
.ZN(net8824)
);

AOI22_X4 c8296(
.A1(net8824),
.A2(net8778),
.B1(net8807),
.ZN(net8825)
);

SDFF_X2 c8297(
.D(net8800),
.SE(net8799),
.SI(net8824),
.CK(clk),
.Q(net8827),
.QN(net8826)
);

OAI22_X4 c8298(
.A1(net8824),
.A2(net8806),
.B1(net8765),
.B2(net10550),
.ZN(net8828)
);

AOI222_X4 c8299(
.A1(net8824),
.A2(net8826),
.B1(net8769),
.B2(net8765),
.C1(net7819),
.C2(net10814),
.ZN(net8829)
);

NOR2_X4 c8300(
.A1(net7919),
.A2(net8789),
.ZN(net8830)
);

NOR2_X2 c8301(
.A1(net7825),
.A2(net6910),
.ZN(net8831)
);

XOR2_X2 c8302(
.A(net8814),
.B(net8763),
.Z(net8832)
);

INV_X32 c8303(
.A(net9794),
.ZN(net8833)
);

XNOR2_X1 c8304(
.A(net8819),
.B(net7948),
.ZN(net8834)
);

OR2_X4 c8305(
.A1(net8792),
.A2(net8814),
.ZN(net8835)
);

OR2_X1 c8306(
.A1(net8812),
.A2(net6927),
.ZN(net8836)
);

INV_X4 c8307(
.A(net3976),
.ZN(net8837)
);

XNOR2_X2 c8308(
.A(net7817),
.B(net5945),
.ZN(net8838)
);

AND2_X4 c8309(
.A1(net8807),
.A2(net8770),
.ZN(net8839)
);

AND2_X1 c8310(
.A1(net5885),
.A2(net8746),
.ZN(net8840)
);

INV_X1 c8311(
.A(net8751),
.ZN(net8841)
);

NAND2_X1 c8312(
.A1(net8836),
.A2(net6980),
.ZN(net8842)
);

INV_X2 c8313(
.A(net7869),
.ZN(net8843)
);

NAND2_X2 c8314(
.A1(net8813),
.A2(net6908),
.ZN(net8844)
);

INV_X8 c8315(
.A(net8763),
.ZN(net8845)
);

NAND2_X4 c8316(
.A1(net6838),
.A2(net3976),
.ZN(net8846)
);

AND2_X2 c8317(
.A1(net8810),
.A2(net11578),
.ZN(net8847)
);

INV_X16 c8318(
.A(net7972),
.ZN(net8848)
);

XOR2_X1 c8319(
.A(net7800),
.B(net8769),
.Z(net8849)
);

NOR2_X1 c8320(
.A1(net8823),
.A2(net6883),
.ZN(net8850)
);

OR2_X2 c8321(
.A1(net8827),
.A2(net11579),
.ZN(net8851)
);

NOR2_X4 c8322(
.A1(net8816),
.A2(net8831),
.ZN(net8852)
);

INV_X32 c8323(
.A(net8847),
.ZN(net8853)
);

NOR2_X2 c8324(
.A1(net8843),
.A2(net7868),
.ZN(net8854)
);

INV_X4 c8325(
.A(net8842),
.ZN(net8855)
);

NAND3_X1 c8326(
.A1(net8853),
.A2(net5898),
.A3(net8852),
.ZN(net8856)
);

XOR2_X2 c8327(
.A(net7948),
.B(net7825),
.Z(net8857)
);

INV_X1 c8328(
.A(net8780),
.ZN(net8858)
);

XNOR2_X1 c8329(
.A(net6911),
.B(net7894),
.ZN(net8859)
);

INV_X2 c8330(
.A(net8789),
.ZN(net8860)
);

INV_X8 c8331(
.A(net9793),
.ZN(net8861)
);

OR2_X4 c8332(
.A1(net8753),
.A2(net8838),
.ZN(net8862)
);

OR2_X1 c8333(
.A1(net8850),
.A2(net8773),
.ZN(net8863)
);

DFFRS_X1 c8334(
.D(net8801),
.RN(net8860),
.SN(net8814),
.CK(clk),
.Q(net8865),
.QN(net8864)
);

NOR3_X4 c8335(
.A1(net8848),
.A2(net6984),
.A3(net7948),
.ZN(net8866)
);

XNOR2_X2 c8336(
.A(net8855),
.B(net8860),
.ZN(net8867)
);

AND2_X4 c8337(
.A1(net7962),
.A2(net10681),
.ZN(net8868)
);

AND2_X1 c8338(
.A1(net8746),
.A2(net8784),
.ZN(net8869)
);

NOR3_X2 c8339(
.A1(net7843),
.A2(net8859),
.A3(net8841),
.ZN(net8870)
);

INV_X16 c8340(
.A(net10054),
.ZN(net8871)
);

NAND2_X1 c8341(
.A1(net8834),
.A2(net8861),
.ZN(net8872)
);

INV_X32 c8342(
.A(net8857),
.ZN(net8873)
);

DFFR_X1 c8343(
.D(net8872),
.RN(net8857),
.CK(clk),
.Q(net8875),
.QN(net8874)
);

NAND2_X2 c8344(
.A1(net8859),
.A2(net8851),
.ZN(net8876)
);

INV_X4 c8345(
.A(net8845),
.ZN(net8877)
);

AND3_X4 c8346(
.A1(net8797),
.A2(net8846),
.A3(net8763),
.ZN(net8878)
);

NAND2_X4 c8347(
.A1(net8770),
.A2(net8763),
.ZN(net8879)
);

AND2_X2 c8348(
.A1(net8876),
.A2(net8859),
.ZN(net8880)
);

INV_X1 c8349(
.A(net10461),
.ZN(net8881)
);

DFFR_X2 c8350(
.D(net8773),
.RN(net8801),
.CK(clk),
.Q(net8883),
.QN(net8882)
);

XOR2_X1 c8351(
.A(net8866),
.B(net8877),
.Z(net8884)
);

NOR2_X1 c8352(
.A1(net7805),
.A2(net8855),
.ZN(net8885)
);

NAND3_X2 c8353(
.A1(net8791),
.A2(net8857),
.A3(net8846),
.ZN(net8886)
);

OR2_X2 c8354(
.A1(net8875),
.A2(net8870),
.ZN(net8887)
);

OR3_X1 c8355(
.A1(net8752),
.A2(net8884),
.A3(net6927),
.ZN(net8888)
);

AOI221_X2 c8356(
.A(net8839),
.B1(net8861),
.B2(net8882),
.C1(net8860),
.C2(net8871),
.ZN(net8889)
);

MUX2_X1 c8357(
.A(net8793),
.B(net8873),
.S(net7900),
.Z(net8890)
);

OAI21_X4 c8358(
.A(net8867),
.B1(net8883),
.B2(net8884),
.ZN(net8891)
);

DFFRS_X2 c8359(
.D(net8886),
.RN(net8810),
.SN(net7800),
.CK(clk),
.Q(net8893),
.QN(net8892)
);

MUX2_X2 c8360(
.A(net8827),
.B(net8875),
.S(net8882),
.Z(net8894)
);

NOR2_X4 c8361(
.A1(net7949),
.A2(net8787),
.ZN(net8895)
);

NAND3_X4 c8362(
.A1(net8870),
.A2(net8893),
.A3(net8861),
.ZN(net8896)
);

OR3_X4 c8363(
.A1(net8895),
.A2(net8894),
.A3(net8892),
.ZN(net8897)
);

AND3_X2 c8364(
.A1(net6885),
.A2(net8896),
.A3(net7972),
.ZN(net8898)
);

NOR3_X1 c8365(
.A1(net6921),
.A2(net6012),
.A3(net8851),
.ZN(net8899)
);

NOR2_X2 c8366(
.A1(net8898),
.A2(net8893),
.ZN(net8900)
);

OR3_X2 c8367(
.A1(net8802),
.A2(net8884),
.A3(net8814),
.ZN(net8901)
);

OAI21_X2 c8368(
.A(net8900),
.B1(net8884),
.B2(net11050),
.ZN(net8902)
);

XOR2_X2 c8369(
.A(net8883),
.B(net8897),
.Z(net8903)
);

OAI21_X1 c8370(
.A(net5839),
.B1(net8808),
.B2(net8900),
.ZN(net8904)
);

XNOR2_X1 c8371(
.A(net8863),
.B(net8830),
.ZN(net8905)
);

AOI21_X2 c8372(
.A(net8903),
.B1(net8885),
.B2(net8797),
.ZN(net8906)
);

SDFF_X1 c8373(
.D(net8873),
.SE(net8905),
.SI(net11096),
.CK(clk),
.Q(net8908),
.QN(net8907)
);

AOI21_X1 c8374(
.A(net8906),
.B1(net8905),
.B2(net8879),
.ZN(net8909)
);

AOI21_X4 c8375(
.A(net8880),
.B1(net8901),
.B2(net7843),
.ZN(net8910)
);

SDFFRS_X2 c8376(
.D(net8899),
.RN(net7961),
.SE(net8897),
.SI(net7889),
.SN(net8748),
.CK(clk),
.Q(net8912),
.QN(net8911)
);

OR2_X4 c8377(
.A1(net8885),
.A2(net8874),
.ZN(net8913)
);

OAI33_X1 c8378(
.A1(net8852),
.A2(net8913),
.A3(net8912),
.B1(net8894),
.B2(net8871),
.B3(net7903),
.ZN(net8914)
);

AND3_X1 c8379(
.A1(net8878),
.A2(net4904),
.A3(net10835),
.ZN(net8915)
);

NAND3_X1 c8380(
.A1(net8900),
.A2(net7934),
.A3(net8908),
.ZN(net8916)
);

SDFFR_X2 c8381(
.D(net8835),
.RN(net8906),
.SE(net7889),
.SI(net10813),
.CK(clk),
.Q(net8918),
.QN(net8917)
);

AOI22_X2 c8382(
.A1(net8917),
.A2(net8911),
.B1(net10680),
.B2(net10786),
.ZN(net8919)
);

OR2_X1 c8383(
.A1(net7052),
.A2(net6984),
.ZN(net8920)
);

XNOR2_X2 c8384(
.A(net7894),
.B(net8784),
.ZN(net8921)
);

AND2_X4 c8385(
.A1(net6961),
.A2(net8897),
.ZN(net8922)
);

AND2_X1 c8386(
.A1(net8871),
.A2(net10769),
.ZN(net8923)
);

NOR3_X4 c8387(
.A1(net7933),
.A2(net8908),
.A3(net8769),
.ZN(net8924)
);

NAND2_X1 c8388(
.A1(net8921),
.A2(net8023),
.ZN(net8925)
);

INV_X2 c8389(
.A(net11375),
.ZN(net8926)
);

INV_X8 c8390(
.A(net8818),
.ZN(net8927)
);

INV_X16 c8391(
.A(net10127),
.ZN(net8928)
);

NAND2_X2 c8392(
.A1(net8835),
.A2(net8008),
.ZN(net8929)
);

NAND2_X4 c8393(
.A1(net8926),
.A2(net7061),
.ZN(net8930)
);

AND2_X2 c8394(
.A1(net7835),
.A2(net5102),
.ZN(net8931)
);

AOI221_X1 c8395(
.A(net8846),
.B1(net8905),
.B2(net8055),
.C1(net8012),
.C2(net8871),
.ZN(net8932)
);

XOR2_X1 c8396(
.A(net8837),
.B(net6097),
.Z(net8933)
);

NOR2_X1 c8397(
.A1(net8840),
.A2(net8912),
.ZN(net8934)
);

OR2_X2 c8398(
.A1(net8008),
.A2(net8927),
.ZN(net8935)
);

NOR2_X4 c8399(
.A1(net8879),
.A2(net8924),
.ZN(net8936)
);

NOR2_X2 c8400(
.A1(net8918),
.A2(net8931),
.ZN(net8937)
);

XOR2_X2 c8401(
.A(net7053),
.B(net8784),
.Z(net8938)
);

XNOR2_X1 c8402(
.A(net8861),
.B(net8769),
.ZN(net8939)
);

INV_X32 c8403(
.A(net10344),
.ZN(net8940)
);

OR2_X4 c8404(
.A1(net7792),
.A2(net8887),
.ZN(net8941)
);

SDFF_X2 c8405(
.D(net8939),
.SE(net7911),
.SI(net8846),
.CK(clk),
.Q(net8943),
.QN(net8942)
);

OR2_X1 c8406(
.A1(net6892),
.A2(net8940),
.ZN(net8944)
);

NOR3_X2 c8407(
.A1(net7962),
.A2(net8931),
.A3(net8935),
.ZN(net8945)
);

XNOR2_X2 c8408(
.A(net8897),
.B(net10630),
.ZN(net8946)
);

INV_X4 c8409(
.A(net10275),
.ZN(net8947)
);

INV_X1 c8410(
.A(net10287),
.ZN(net8948)
);

AND2_X4 c8411(
.A1(net5120),
.A2(net8946),
.ZN(net8949)
);

AND2_X1 c8412(
.A1(net7061),
.A2(net8861),
.ZN(net8950)
);

NAND2_X1 c8413(
.A1(net8754),
.A2(net8881),
.ZN(net8951)
);

AND3_X4 c8414(
.A1(net8833),
.A2(net8057),
.A3(net6908),
.ZN(net8952)
);

NAND2_X2 c8415(
.A1(net8881),
.A2(net8943),
.ZN(net8953)
);

NAND3_X2 c8416(
.A1(net8950),
.A2(net8817),
.A3(net7792),
.ZN(net8954)
);

OR3_X1 c8417(
.A1(net7928),
.A2(net7980),
.A3(net8953),
.ZN(net8955)
);

NAND2_X4 c8418(
.A1(net8787),
.A2(net8951),
.ZN(net8956)
);

AND2_X2 c8419(
.A1(net8907),
.A2(net11244),
.ZN(net8957)
);

INV_X2 c8420(
.A(net10126),
.ZN(net8958)
);

XOR2_X1 c8421(
.A(net8784),
.B(net8889),
.Z(net8959)
);

INV_X8 c8422(
.A(net9694),
.ZN(net8960)
);

NOR2_X1 c8423(
.A1(net6999),
.A2(net7019),
.ZN(net8961)
);

OAI221_X1 c8424(
.A(net8854),
.B1(net3976),
.B2(net8920),
.C1(net8911),
.C2(net11244),
.ZN(net8962)
);

SDFFS_X1 c8425(
.D(net7942),
.SE(net8933),
.SI(net8935),
.SN(net8931),
.CK(clk),
.Q(net8964),
.QN(net8963)
);

DFFRS_X1 c8426(
.D(net8957),
.RN(net8925),
.SN(net8961),
.CK(clk),
.Q(net8966),
.QN(net8965)
);

SDFFS_X2 c8427(
.D(net8891),
.SE(net8961),
.SI(net8894),
.SN(net8911),
.CK(clk),
.Q(net8968),
.QN(net8967)
);

OR2_X2 c8428(
.A1(net8935),
.A2(net8057),
.ZN(net8969)
);

OAI221_X4 c8429(
.A(net8890),
.B1(net8955),
.B2(net8919),
.C1(net7903),
.C2(net8860),
.ZN(net8970)
);

NOR2_X4 c8430(
.A1(net8933),
.A2(net11310),
.ZN(net8971)
);

NOR2_X2 c8431(
.A1(net8894),
.A2(net8967),
.ZN(net8972)
);

MUX2_X1 c8432(
.A(net6908),
.B(net8748),
.S(net8831),
.Z(net8973)
);

NAND4_X4 c8433(
.A1(net8808),
.A2(net7982),
.A3(net8925),
.A4(net8785),
.ZN(net8974)
);

OAI221_X2 c8434(
.A(net8947),
.B1(net8945),
.B2(net8963),
.C1(net6098),
.C2(net8750),
.ZN(net8975)
);

OAI21_X4 c8435(
.A(net8964),
.B1(net8931),
.B2(net8933),
.ZN(net8976)
);

DFFS_X1 c8436(
.D(net8769),
.SN(net8004),
.CK(clk),
.Q(net8978),
.QN(net8977)
);

XOR2_X2 c8437(
.A(net8805),
.B(net11162),
.Z(net8979)
);

XNOR2_X1 c8438(
.A(net8930),
.B(net8946),
.ZN(net8980)
);

INV_X16 c8439(
.A(net11375),
.ZN(net8981)
);

OR2_X4 c8440(
.A1(net8868),
.A2(net8055),
.ZN(net8982)
);

OR2_X1 c8441(
.A1(net8944),
.A2(net7982),
.ZN(net8983)
);

INV_X32 c8442(
.A(net10444),
.ZN(net8984)
);

XNOR2_X2 c8443(
.A(net8958),
.B(net8966),
.ZN(net8985)
);

AND2_X4 c8444(
.A1(net8985),
.A2(net6050),
.ZN(net8986)
);

AND2_X1 c8445(
.A1(net7982),
.A2(net8945),
.ZN(net8987)
);

NAND2_X1 c8446(
.A1(net8951),
.A2(net8897),
.ZN(net8988)
);

NAND2_X2 c8447(
.A1(net8988),
.A2(net11077),
.ZN(net8989)
);

NAND2_X4 c8448(
.A1(net8948),
.A2(net8908),
.ZN(net8990)
);

MUX2_X2 c8449(
.A(net8956),
.B(net8964),
.S(net8988),
.Z(net8991)
);

AND2_X2 c8450(
.A1(net8988),
.A2(net8918),
.ZN(net8992)
);

XOR2_X1 c8451(
.A(net8055),
.B(net11310),
.Z(net8993)
);

INV_X4 c8452(
.A(net9693),
.ZN(net8994)
);

NAND3_X4 c8453(
.A1(net8844),
.A2(net8968),
.A3(net8933),
.ZN(net8995)
);

OR3_X4 c8454(
.A1(net8994),
.A2(net8952),
.A3(net8985),
.ZN(net8996)
);

INV_X1 c8455(
.A(net10191),
.ZN(net8997)
);

NOR2_X1 c8456(
.A1(net8962),
.A2(net8985),
.ZN(net8998)
);

AND3_X2 c8457(
.A1(net7019),
.A2(net7928),
.A3(net11391),
.ZN(net8999)
);

OR2_X2 c8458(
.A1(net8979),
.A2(net8981),
.ZN(net9000)
);

NOR3_X1 c8459(
.A1(net7066),
.A2(net8963),
.A3(net10629),
.ZN(net9001)
);

NOR2_X4 c8460(
.A1(net9001),
.A2(net8992),
.ZN(net9002)
);

NOR2_X2 c8461(
.A1(net8869),
.A2(net7013),
.ZN(net9003)
);

OR3_X2 c8462(
.A1(net8987),
.A2(net8998),
.A3(net8965),
.ZN(net9004)
);

SDFFR_X1 c8463(
.D(net8057),
.RN(net8993),
.SE(net8869),
.SI(net8983),
.CK(clk),
.Q(net9006),
.QN(net9005)
);

SDFFRS_X1 c8464(
.D(net9002),
.RN(net9000),
.SE(net9003),
.SI(net8985),
.SN(net7812),
.CK(clk),
.Q(net9008),
.QN(net9007)
);

XOR2_X2 c8465(
.A(net8969),
.B(net9007),
.Z(net9009)
);

INV_X2 c8466(
.A(net11331),
.ZN(net9010)
);

XNOR2_X1 c8467(
.A(net6980),
.B(net8997),
.ZN(net9011)
);

INV_X8 c8468(
.A(net11249),
.ZN(net9012)
);

OR2_X4 c8469(
.A1(net7078),
.A2(net8098),
.ZN(net9013)
);

OAI21_X2 c8470(
.A(net7988),
.B1(net8757),
.B2(net7820),
.ZN(net9014)
);

OAI21_X1 c8471(
.A(net8118),
.B1(net8961),
.B2(net11247),
.ZN(net9015)
);

INV_X16 c8472(
.A(net11388),
.ZN(net9016)
);

OR2_X1 c8473(
.A1(net9015),
.A2(net11478),
.ZN(net9017)
);

INV_X32 c8474(
.A(net10368),
.ZN(net9018)
);

AOI21_X2 c8475(
.A(net8887),
.B1(net8984),
.B2(net8943),
.ZN(net9019)
);

XNOR2_X2 c8476(
.A(net7934),
.B(net8087),
.ZN(net9020)
);

AOI21_X1 c8477(
.A(net8143),
.B1(net8997),
.B2(net8931),
.ZN(net9021)
);

AND2_X4 c8478(
.A1(net7979),
.A2(net7078),
.ZN(net9022)
);

AND2_X1 c8479(
.A1(net8093),
.A2(net8076),
.ZN(net9023)
);

AOI21_X4 c8480(
.A(net4140),
.B1(net9023),
.B2(net8945),
.ZN(net9024)
);

NAND2_X1 c8481(
.A1(net5945),
.A2(net8851),
.ZN(net9025)
);

NAND2_X2 c8482(
.A1(net6170),
.A2(net9019),
.ZN(net9026)
);

AND3_X1 c8483(
.A1(net7160),
.A2(net6927),
.A3(net8750),
.ZN(net9027)
);

NAND2_X4 c8484(
.A1(net7907),
.A2(net11489),
.ZN(net9028)
);

AND2_X2 c8485(
.A1(net7159),
.A2(net8045),
.ZN(net9029)
);

NAND3_X1 c8486(
.A1(net7985),
.A2(net8748),
.A3(net11025),
.ZN(net9030)
);

DFFRS_X2 c8487(
.D(net7122),
.RN(net8945),
.SN(net8851),
.CK(clk),
.Q(net9032),
.QN(net9031)
);

DFFS_X2 c8488(
.D(net6098),
.SN(net8999),
.CK(clk),
.Q(net9034),
.QN(net9033)
);

NOR3_X4 c8489(
.A1(net8858),
.A2(net8838),
.A3(net7886),
.ZN(net9035)
);

NOR3_X2 c8490(
.A1(net8080),
.A2(net8946),
.A3(net8805),
.ZN(net9036)
);

XOR2_X1 c8491(
.A(net7037),
.B(net11173),
.Z(net9037)
);

SDFF_X1 c8492(
.D(net9014),
.SE(net8113),
.SI(net8919),
.CK(clk),
.Q(net9039),
.QN(net9038)
);

AND3_X4 c8493(
.A1(net9027),
.A2(net8012),
.A3(net7934),
.ZN(net9040)
);

NAND3_X2 c8494(
.A1(net8923),
.A2(net9028),
.A3(net8871),
.ZN(net9041)
);

NOR2_X1 c8495(
.A1(net8978),
.A2(net9005),
.ZN(net9042)
);

DFFR_X1 c8496(
.D(net8113),
.RN(net9012),
.CK(clk),
.Q(net9044),
.QN(net9043)
);

SDFF_X2 c8497(
.D(net8888),
.SE(net8098),
.SI(net9027),
.CK(clk),
.Q(net9046),
.QN(net9045)
);

OR2_X2 c8498(
.A1(net7137),
.A2(net5945),
.ZN(net9047)
);

OR3_X1 c8499(
.A1(net8050),
.A2(net8977),
.A3(net8938),
.ZN(net9048)
);

NOR2_X4 c8500(
.A1(net8076),
.A2(net8757),
.ZN(net9049)
);

NOR2_X2 c8501(
.A1(net9040),
.A2(net7980),
.ZN(net9050)
);

INV_X4 c8502(
.A(net10369),
.ZN(net9051)
);

XOR2_X2 c8503(
.A(net8978),
.B(net11042),
.Z(net9052)
);

XNOR2_X1 c8504(
.A(net9052),
.B(net9008),
.ZN(net9053)
);

OR2_X4 c8505(
.A1(net8968),
.A2(net9003),
.ZN(net9054)
);

OR2_X1 c8506(
.A1(net8750),
.A2(net8966),
.ZN(net9055)
);

XNOR2_X2 c8507(
.A(net7037),
.B(net9050),
.ZN(net9056)
);

AND2_X4 c8508(
.A1(net9009),
.A2(net9015),
.ZN(net9057)
);

DFFRS_X1 c8509(
.D(net7820),
.RN(net9045),
.SN(net9026),
.CK(clk),
.Q(net9059),
.QN(net9058)
);

MUX2_X1 c8510(
.A(net9022),
.B(net7078),
.S(net8865),
.Z(net9060)
);

AND2_X1 c8511(
.A1(net8111),
.A2(net11127),
.ZN(net9061)
);

INV_X1 c8512(
.A(net10410),
.ZN(net9062)
);

DFFR_X2 c8513(
.D(net9048),
.RN(net8757),
.CK(clk),
.Q(net9064),
.QN(net9063)
);

NAND2_X1 c8514(
.A1(net9059),
.A2(net8960),
.ZN(net9065)
);

OAI21_X4 c8515(
.A(net9020),
.B1(net8830),
.B2(net7137),
.ZN(net9066)
);

MUX2_X2 c8516(
.A(net9044),
.B(net8997),
.S(net8940),
.Z(net9067)
);

NAND2_X2 c8517(
.A1(net7019),
.A2(net9064),
.ZN(net9068)
);

NAND2_X4 c8518(
.A1(net9068),
.A2(net8940),
.ZN(net9069)
);

AND2_X2 c8519(
.A1(net8990),
.A2(net8858),
.ZN(net9070)
);

XOR2_X1 c8520(
.A(net9066),
.B(net9069),
.Z(net9071)
);

NOR2_X1 c8521(
.A1(net9067),
.A2(net8785),
.ZN(net9072)
);

NAND3_X4 c8522(
.A1(net7985),
.A2(net8118),
.A3(net8888),
.ZN(net9073)
);

OR3_X4 c8523(
.A1(net9017),
.A2(net8865),
.A3(net9015),
.ZN(net9074)
);

INV_X2 c8524(
.A(net11249),
.ZN(net9075)
);

OR2_X2 c8525(
.A1(net8931),
.A2(net11026),
.ZN(net9076)
);

OAI211_X2 c8526(
.A(net9068),
.B(net9043),
.C1(net8133),
.C2(net11435),
.ZN(net9077)
);

NOR2_X4 c8527(
.A1(net9065),
.A2(net7084),
.ZN(net9078)
);

NOR2_X2 c8528(
.A1(net9062),
.A2(net11009),
.ZN(net9079)
);

DFFRS_X2 c8529(
.D(net9079),
.RN(net9026),
.SN(net9075),
.CK(clk),
.Q(net9081),
.QN(net9080)
);

AND3_X2 c8530(
.A1(net8750),
.A2(net9014),
.A3(net10897),
.ZN(net9082)
);

NOR3_X1 c8531(
.A1(net7979),
.A2(net9065),
.A3(net11414),
.ZN(net9083)
);

OR3_X2 c8532(
.A1(net9050),
.A2(net9061),
.A3(net9077),
.ZN(net9084)
);

XOR2_X2 c8533(
.A(net9046),
.B(net9076),
.Z(net9085)
);

SDFF_X1 c8534(
.D(net8838),
.SE(net9058),
.SI(net8983),
.CK(clk),
.Q(net9087),
.QN(net9086)
);

SDFF_X2 c8535(
.D(net8830),
.SE(net9070),
.SI(net9087),
.CK(clk),
.Q(net9089),
.QN(net9088)
);

OAI21_X2 c8536(
.A(net9075),
.B1(net9059),
.B2(net9086),
.ZN(net9090)
);

OAI21_X1 c8537(
.A(net9025),
.B1(net9085),
.B2(net9087),
.ZN(net9091)
);

AOI21_X2 c8538(
.A(net7109),
.B1(net9087),
.B2(net8079),
.ZN(net9092)
);

AOI21_X1 c8539(
.A(net9076),
.B1(net10890),
.B2(net10927),
.ZN(net9093)
);

AOI21_X4 c8540(
.A(net9083),
.B1(net9068),
.B2(net9019),
.ZN(net9094)
);

AND3_X1 c8541(
.A1(net8945),
.A2(net9042),
.A3(net11247),
.ZN(net9095)
);

NAND3_X1 c8542(
.A1(net9078),
.A2(net9089),
.A3(net10975),
.ZN(net9096)
);

DFFRS_X1 c8543(
.D(net9095),
.RN(net11097),
.SN(net11488),
.CK(clk),
.Q(net9098),
.QN(net9097)
);

NOR3_X4 c8544(
.A1(net9035),
.A2(net9094),
.A3(net9097),
.ZN(net9099)
);

OR4_X2 c8545(
.A1(net9060),
.A2(net9072),
.A3(net9020),
.A4(net8911),
.ZN(net9100)
);

XNOR2_X1 c8546(
.A(net8105),
.B(net10762),
.ZN(net9101)
);

AOI221_X4 c8547(
.A(net9101),
.B1(net9096),
.B2(net9090),
.C1(net9086),
.C2(net8091),
.ZN(net9102)
);

NOR3_X2 c8548(
.A1(net9086),
.A2(net10627),
.A3(net10742),
.ZN(net9103)
);

AND3_X4 c8549(
.A1(net8045),
.A2(net9081),
.A3(net9038),
.ZN(net9104)
);

NAND3_X2 c8550(
.A1(net8231),
.A2(net9026),
.A3(net9077),
.ZN(net9105)
);

INV_X8 c8551(
.A(net11329),
.ZN(net9106)
);

OR2_X4 c8552(
.A1(net6927),
.A2(net9008),
.ZN(net9107)
);

OR2_X1 c8553(
.A1(net8149),
.A2(net8993),
.ZN(net9108)
);

XNOR2_X2 c8554(
.A(net8166),
.B(net9063),
.ZN(net9109)
);

OR3_X1 c8555(
.A1(net8928),
.A2(net9108),
.A3(net9088),
.ZN(net9110)
);

AND2_X4 c8556(
.A1(net9034),
.A2(net8959),
.ZN(net9111)
);

MUX2_X1 c8557(
.A(net9041),
.B(net9089),
.S(net8991),
.Z(net9112)
);

OAI21_X4 c8558(
.A(net7907),
.B1(net8989),
.B2(net9108),
.ZN(net9113)
);

AOI222_X2 c8559(
.A1(net8938),
.A2(net5234),
.B1(net9107),
.B2(net9026),
.C1(net9051),
.C2(net9080),
.ZN(net9114)
);

MUX2_X2 c8560(
.A(net8035),
.B(net9012),
.S(net8126),
.Z(net9115)
);

NAND3_X4 c8561(
.A1(net8993),
.A2(net9110),
.A3(net9055),
.ZN(net9116)
);

AND2_X1 c8562(
.A1(net8785),
.A2(net9116),
.ZN(net9117)
);

DFFS_X1 c8563(
.D(net8884),
.SN(net9026),
.CK(clk),
.Q(net9119),
.QN(net9118)
);

OR3_X4 c8564(
.A1(net7886),
.A2(net9119),
.A3(net8965),
.ZN(net9120)
);

INV_X16 c8565(
.A(net10441),
.ZN(net9121)
);

AND3_X2 c8566(
.A1(net9029),
.A2(net8035),
.A3(net8222),
.ZN(net9122)
);

NAND2_X1 c8567(
.A1(net9051),
.A2(net9011),
.ZN(net9123)
);

NOR3_X1 c8568(
.A1(net8991),
.A2(net8785),
.A3(net8232),
.ZN(net9124)
);

INV_X32 c8569(
.A(net10499),
.ZN(net9125)
);

NAND2_X2 c8570(
.A1(net8058),
.A2(net8946),
.ZN(net9126)
);

OR3_X2 c8571(
.A1(net9053),
.A2(net9097),
.A3(net11076),
.ZN(net9127)
);

NAND2_X4 c8572(
.A1(net9055),
.A2(net8919),
.ZN(net9128)
);

AND2_X2 c8573(
.A1(net8982),
.A2(net9082),
.ZN(net9129)
);

OAI21_X2 c8574(
.A(net9126),
.B1(net8233),
.B2(net8133),
.ZN(net9130)
);

OAI21_X1 c8575(
.A(net8229),
.B1(net8884),
.B2(net11568),
.ZN(net9131)
);

AOI21_X2 c8576(
.A(net8233),
.B1(net8805),
.B2(net6011),
.ZN(net9132)
);

AOI21_X1 c8577(
.A(net6175),
.B1(net9094),
.B2(net7184),
.ZN(net9133)
);

XOR2_X1 c8578(
.A(net8087),
.B(net8112),
.Z(net9134)
);

AOI21_X4 c8579(
.A(net9006),
.B1(net9102),
.B2(net11033),
.ZN(net9135)
);

DFFRS_X2 c8580(
.D(net8966),
.RN(net9103),
.SN(net7176),
.CK(clk),
.Q(net9137),
.QN(net9136)
);

NOR2_X1 c8581(
.A1(net11041),
.A2(net11569),
.ZN(net9138)
);

AND3_X1 c8582(
.A1(net8152),
.A2(net9106),
.A3(net9021),
.ZN(net9139)
);

OAI222_X1 c8583(
.A1(net8079),
.A2(net9021),
.B1(net9107),
.B2(net9138),
.C1(net9122),
.C2(net8213),
.ZN(net9140)
);

NAND3_X1 c8584(
.A1(net8169),
.A2(net8748),
.A3(net9021),
.ZN(net9141)
);

OR2_X2 c8585(
.A1(net8060),
.A2(net9032),
.ZN(net9142)
);

NOR3_X4 c8586(
.A1(net9003),
.A2(net9132),
.A3(net8841),
.ZN(net9143)
);

NOR3_X2 c8587(
.A1(net8174),
.A2(net7889),
.A3(net8192),
.ZN(net9144)
);

AND3_X4 c8588(
.A1(net9128),
.A2(net9106),
.A3(net8222),
.ZN(net9145)
);

SDFF_X1 c8589(
.D(net9119),
.SE(net9116),
.SI(net8222),
.CK(clk),
.Q(net9147),
.QN(net9146)
);

SDFF_X2 c8590(
.D(net7903),
.SE(net9129),
.SI(net7176),
.CK(clk),
.Q(net9149),
.QN(net9148)
);

DFFRS_X1 c8591(
.D(net9070),
.RN(net9148),
.SN(net10974),
.CK(clk),
.Q(net9151),
.QN(net9150)
);

NAND3_X2 c8592(
.A1(net9144),
.A2(net9129),
.A3(net8058),
.ZN(net9152)
);

OR3_X1 c8593(
.A1(net7176),
.A2(net9130),
.A3(net8785),
.ZN(net9153)
);

MUX2_X1 c8594(
.A(net9016),
.B(net9132),
.S(net8109),
.Z(net9154)
);

OAI21_X4 c8595(
.A(net8953),
.B1(net9134),
.B2(net6175),
.ZN(net9155)
);

MUX2_X2 c8596(
.A(net8748),
.B(net8831),
.S(net9124),
.Z(net9156)
);

NAND3_X4 c8597(
.A1(net8937),
.A2(net8235),
.A3(net9013),
.ZN(net9157)
);

DFFRS_X2 c8598(
.D(net9006),
.RN(net9124),
.SN(net11559),
.CK(clk),
.Q(net9159),
.QN(net9158)
);

OR3_X4 c8599(
.A1(net9155),
.A2(net8952),
.A3(net9136),
.ZN(net9160)
);

AND3_X2 c8600(
.A1(net8222),
.A2(net9154),
.A3(net9136),
.ZN(net9161)
);

NOR3_X1 c8601(
.A1(net8126),
.A2(net8952),
.A3(net9150),
.ZN(net9162)
);

SDFF_X1 c8602(
.D(net8946),
.SE(net9112),
.SI(net9039),
.CK(clk),
.Q(net9164),
.QN(net9163)
);

OR3_X2 c8603(
.A1(net9115),
.A2(net9110),
.A3(net11172),
.ZN(net9165)
);

SDFF_X2 c8604(
.D(net9124),
.SE(net9134),
.SI(net9033),
.CK(clk),
.Q(net9167),
.QN(net9166)
);

INV_X4 c8605(
.A(net11329),
.ZN(net9168)
);

INV_X1 c8606(
.A(net10143),
.ZN(net9169)
);

OAI21_X2 c8607(
.A(net8919),
.B1(net9121),
.B2(net11559),
.ZN(net9170)
);

AOI221_X2 c8608(
.A(net8213),
.B1(net8166),
.B2(net9138),
.C1(net9146),
.C2(net9032),
.ZN(net9171)
);

OAI222_X4 c8609(
.A1(net8112),
.A2(net9164),
.B1(net9162),
.B2(net9077),
.C1(net9090),
.C2(net9122),
.ZN(net9172)
);

DFFRS_X1 c8610(
.D(net9057),
.RN(net7980),
.SN(net9162),
.CK(clk),
.Q(net9174),
.QN(net9173)
);

INV_X2 c8611(
.A(net9846),
.ZN(net9175)
);

OAI21_X1 c8612(
.A(net8757),
.B1(net9095),
.B2(net11376),
.ZN(net9176)
);

AOI21_X2 c8613(
.A(net9161),
.B1(net9165),
.B2(net9163),
.ZN(net9177)
);

DFFRS_X2 c8614(
.D(net9070),
.RN(net9174),
.SN(net8200),
.CK(clk),
.Q(net9179),
.QN(net9178)
);

OAI222_X2 c8615(
.A1(net9104),
.A2(net9179),
.B1(net9166),
.B2(net9088),
.C1(net9122),
.C2(net8207),
.ZN(net9180)
);

INV_X8 c8616(
.A(net9981),
.ZN(net9181)
);

AOI21_X1 c8617(
.A(net9010),
.B1(net8785),
.B2(net10909),
.ZN(net9182)
);

AOI21_X4 c8618(
.A(net9162),
.B1(net9181),
.B2(net9168),
.ZN(net9183)
);

AND3_X1 c8619(
.A1(net9169),
.A2(net9088),
.A3(net10926),
.ZN(net9184)
);

NAND3_X1 c8620(
.A1(net9124),
.A2(net9175),
.A3(net10554),
.ZN(net9185)
);

NOR3_X4 c8621(
.A1(net9164),
.A2(net8919),
.A3(net11330),
.ZN(net9186)
);

NOR3_X2 c8622(
.A1(net9182),
.A2(net9016),
.A3(net11433),
.ZN(net9187)
);

AND3_X4 c8623(
.A1(net9175),
.A2(net9181),
.A3(net11163),
.ZN(net9188)
);

SDFF_X1 c8624(
.D(net9131),
.SE(net9127),
.SI(net9173),
.CK(clk),
.Q(net9190),
.QN(net9189)
);

NAND3_X2 c8625(
.A1(net9103),
.A2(net9190),
.A3(net11330),
.ZN(net9191)
);

SDFF_X2 c8626(
.D(net9187),
.SE(net9154),
.SI(net9131),
.CK(clk),
.Q(net9193),
.QN(net9192)
);

OR3_X1 c8627(
.A1(net9191),
.A2(net9178),
.A3(net9170),
.ZN(net9194)
);

MUX2_X1 c8628(
.A(net9145),
.B(net9093),
.S(net11032),
.Z(net9195)
);

OAI21_X4 c8629(
.A(net9188),
.B1(net9122),
.B2(net11261),
.ZN(net9196)
);

DFFS_X2 c8630(
.D(net9095),
.SN(net9194),
.CK(clk),
.Q(net9198),
.QN(net9197)
);

DFFRS_X1 c8631(
.D(net9113),
.RN(net9170),
.SN(net10555),
.CK(clk),
.Q(net9200),
.QN(net9199)
);

MUX2_X2 c8632(
.A(net9135),
.B(net8983),
.S(net9036),
.Z(net9201)
);

NOR2_X4 c8633(
.A1(net8153),
.A2(net9098),
.ZN(net9202)
);

NAND3_X4 c8634(
.A1(net9186),
.A2(net9135),
.A3(net8292),
.ZN(net9203)
);

INV_X16 c8635(
.A(net11453),
.ZN(net9204)
);

INV_X32 c8636(
.A(net11453),
.ZN(net9205)
);

NOR2_X2 c8637(
.A1(net9110),
.A2(net8920),
.ZN(net9206)
);

OR3_X4 c8638(
.A1(net9109),
.A2(net8961),
.A3(net8299),
.ZN(net9207)
);

AND3_X2 c8639(
.A1(net9192),
.A2(net9166),
.A3(net11409),
.ZN(net9208)
);

NOR3_X1 c8640(
.A1(net8193),
.A2(net9012),
.A3(net11454),
.ZN(net9209)
);

XOR2_X2 c8641(
.A(net9081),
.B(net7309),
.Z(net9210)
);

DFFRS_X2 c8642(
.D(net8201),
.RN(net9150),
.SN(net9202),
.CK(clk),
.Q(net9212),
.QN(net9211)
);

XNOR2_X1 c8643(
.A(net9200),
.B(net6851),
.ZN(net9213)
);

INV_X4 c8644(
.A(net10360),
.ZN(net9214)
);

OR2_X4 c8645(
.A1(net9013),
.A2(net9151),
.ZN(net9215)
);

OR2_X1 c8646(
.A1(net9108),
.A2(net9102),
.ZN(net9216)
);

XNOR2_X2 c8647(
.A(net7287),
.B(net9204),
.ZN(net9217)
);

SDFF_X1 c8648(
.D(net7184),
.SE(net8201),
.SI(net9216),
.CK(clk),
.Q(net9219),
.QN(net9218)
);

AND2_X4 c8649(
.A1(net8961),
.A2(net9208),
.ZN(net9220)
);

OR3_X2 c8650(
.A1(net9149),
.A2(net8912),
.A3(net8091),
.ZN(net9221)
);

AND2_X1 c8651(
.A1(net8299),
.A2(net7211),
.ZN(net9222)
);

NAND2_X1 c8652(
.A1(net8278),
.A2(net9207),
.ZN(net9223)
);

NAND2_X2 c8653(
.A1(net8193),
.A2(net7184),
.ZN(net9224)
);

NAND2_X4 c8654(
.A1(net8295),
.A2(net9190),
.ZN(net9225)
);

AND2_X2 c8655(
.A1(net8249),
.A2(net8310),
.ZN(net9226)
);

SDFFR_X2 c8656(
.D(net8292),
.RN(net9167),
.SE(net9211),
.SI(net9012),
.CK(clk),
.Q(net9228),
.QN(net9227)
);

XOR2_X1 c8657(
.A(net8256),
.B(net9227),
.Z(net9229)
);

OAI21_X2 c8658(
.A(net9082),
.B1(net9121),
.B2(net9229),
.ZN(net9230)
);

NOR2_X1 c8659(
.A1(net9228),
.A2(net9120),
.ZN(net9231)
);

OAI21_X1 c8660(
.A(net9168),
.B1(net9219),
.B2(net9199),
.ZN(net9232)
);

AOI21_X2 c8661(
.A(net9100),
.B1(net8091),
.B2(net10628),
.ZN(net9233)
);

AOI21_X1 c8662(
.A(net9224),
.B1(net8059),
.B2(net11438),
.ZN(net9234)
);

OR2_X2 c8663(
.A1(net9107),
.A2(net11196),
.ZN(net9235)
);

AOI21_X4 c8664(
.A(net8841),
.B1(net8059),
.B2(net9170),
.ZN(net9236)
);

AND3_X1 c8665(
.A1(net9222),
.A2(net8283),
.A3(net8249),
.ZN(net9237)
);

NAND3_X1 c8666(
.A1(net9221),
.A2(net9193),
.A3(net9138),
.ZN(net9238)
);

NOR3_X4 c8667(
.A1(net9206),
.A2(net9236),
.A3(net9202),
.ZN(net9239)
);

NOR3_X2 c8668(
.A1(net9232),
.A2(net9235),
.A3(net8192),
.ZN(net9240)
);

NOR2_X4 c8669(
.A1(net8098),
.A2(net8212),
.ZN(net9241)
);

AND3_X4 c8670(
.A1(net8851),
.A2(net9013),
.A3(net9018),
.ZN(net9242)
);

NAND3_X2 c8671(
.A1(net9229),
.A2(net9137),
.A3(net5383),
.ZN(net9243)
);

SDFF_X2 c8672(
.D(net9159),
.SE(net9236),
.SI(net8059),
.CK(clk),
.Q(net9245),
.QN(net9244)
);

OR3_X1 c8673(
.A1(net9039),
.A2(net9224),
.A3(net8248),
.ZN(net9246)
);

MUX2_X1 c8674(
.A(net8091),
.B(net8860),
.S(net9218),
.Z(net9247)
);

OAI21_X4 c8675(
.A(net9120),
.B1(net9209),
.B2(net9224),
.ZN(net9248)
);

MUX2_X2 c8676(
.A(net9241),
.B(net8201),
.S(net6354),
.Z(net9249)
);

NAND3_X4 c8677(
.A1(net8912),
.A2(net9225),
.A3(net8841),
.ZN(net9250)
);

AOI222_X1 c8678(
.A1(net9210),
.A2(net8059),
.B1(net8295),
.B2(net9224),
.C1(net9202),
.C2(net9189),
.ZN(net9251)
);

OR3_X4 c8679(
.A1(net9234),
.A2(net9246),
.A3(net8292),
.ZN(net9252)
);

NOR2_X2 c8680(
.A1(net8133),
.A2(net8278),
.ZN(net9253)
);

AND3_X2 c8681(
.A1(net7309),
.A2(net9248),
.A3(net9158),
.ZN(net9254)
);

NOR3_X1 c8682(
.A1(net9147),
.A2(net9250),
.A3(net9202),
.ZN(net9255)
);

DFFRS_X1 c8683(
.D(net9142),
.RN(net5383),
.SN(net9244),
.CK(clk),
.Q(net9257),
.QN(net9256)
);

XOR2_X2 c8684(
.A(net9012),
.B(net8984),
.Z(net9258)
);

OR3_X2 c8685(
.A1(net8212),
.A2(net9256),
.A3(net11454),
.ZN(net9259)
);

OAI21_X2 c8686(
.A(net9121),
.B1(net9109),
.B2(net10869),
.ZN(net9260)
);

OAI21_X1 c8687(
.A(net9259),
.B1(net9250),
.B2(net9241),
.ZN(net9261)
);

XNOR2_X1 c8688(
.A(net11128),
.B(net11197),
.ZN(net9262)
);

OR2_X4 c8689(
.A1(net7889),
.A2(net9247),
.ZN(net9263)
);

AOI21_X2 c8690(
.A(net8283),
.B1(net7331),
.B2(net8274),
.ZN(net9264)
);

AOI21_X1 c8691(
.A(net9263),
.B1(net9261),
.B2(net9246),
.ZN(net9265)
);

AOI21_X4 c8692(
.A(net6966),
.B1(net8998),
.B2(net9181),
.ZN(net9266)
);

AND3_X1 c8693(
.A1(net8315),
.A2(net9205),
.A3(net9122),
.ZN(net9267)
);

OR2_X1 c8694(
.A1(net9265),
.A2(net9018),
.ZN(net9268)
);

AOI211_X1 c8695(
.A(net9260),
.B(net9214),
.C1(out13),
.C2(net11409),
.ZN(net9269)
);

NAND3_X1 c8696(
.A1(net9213),
.A2(net9262),
.A3(net9244),
.ZN(net9270)
);

NOR3_X4 c8697(
.A1(net8984),
.A2(net9254),
.A3(net9263),
.ZN(net9271)
);

NOR3_X2 c8698(
.A1(net9242),
.A2(net9270),
.A3(net8283),
.ZN(net9272)
);

AND3_X4 c8699(
.A1(net9270),
.A2(net8960),
.A3(net8315),
.ZN(net9273)
);

NAND3_X2 c8700(
.A1(net8998),
.A2(net9273),
.A3(net9147),
.ZN(net9274)
);

OR3_X1 c8701(
.A1(net9272),
.A2(net9229),
.A3(net11094),
.ZN(net9275)
);

XNOR2_X2 c8702(
.A(net9260),
.B(net9247),
.ZN(net9276)
);

NAND4_X2 c8703(
.A1(net7331),
.A2(net9276),
.A3(net9270),
.A4(net9122),
.ZN(net9277)
);

MUX2_X1 c8704(
.A(net9093),
.B(net9261),
.S(net9216),
.Z(net9278)
);

OAI21_X4 c8705(
.A(net9250),
.B1(net9270),
.B2(net10868),
.ZN(net9279)
);

MUX2_X2 c8706(
.A(net9151),
.B(net8960),
.S(net8212),
.Z(net9280)
);

SDFFRS_X2 c8707(
.D(net9231),
.RN(net9271),
.SE(net9264),
.SI(net9100),
.SN(net8279),
.CK(clk),
.Q(net9282),
.QN(net9281)
);

NAND3_X4 c8708(
.A1(net8251),
.A2(net9262),
.A3(net9257),
.ZN(net9283)
);

OR4_X4 c8709(
.A1(net9258),
.A2(net9273),
.A3(net9281),
.A4(net11194),
.ZN(net9284)
);

OR3_X4 c8710(
.A1(net9125),
.A2(net9246),
.A3(net9276),
.ZN(net9285)
);

AND3_X2 c8711(
.A1(net9284),
.A2(net9280),
.A3(net10980),
.ZN(net9286)
);

OAI22_X2 c8712(
.A1(net9286),
.A2(net9276),
.B1(net9102),
.B2(net11095),
.ZN(net9287)
);

NOR3_X1 c8713(
.A1(net9254),
.A2(net9257),
.A3(net8091),
.ZN(net9288)
);

AOI222_X4 c8714(
.A1(net9269),
.A2(net9288),
.B1(net9287),
.B2(net9216),
.C1(net9189),
.C2(net9202),
.ZN(net9289)
);

AND2_X4 c8715(
.A1(net9226),
.A2(net10921),
.ZN(net9290)
);

OAI211_X4 c8716(
.A(net8337),
.B(net9138),
.C1(net8983),
.C2(net9224),
.ZN(net9291)
);

AND2_X1 c8717(
.A1(net8275),
.A2(net9290),
.ZN(net9292)
);

DFFRS_X2 c8718(
.D(net9089),
.RN(net9122),
.SN(net8831),
.CK(clk),
.Q(net9294),
.QN(net9293)
);

INV_X1 c8719(
.A(net11354),
.ZN(net9295)
);

OR3_X2 c8720(
.A1(net9047),
.A2(net7812),
.A3(net9122),
.ZN(net9296)
);

SDFF_X1 c8721(
.D(net8405),
.SE(net9287),
.SI(net9100),
.CK(clk),
.Q(net9298),
.QN(net9297)
);

NAND2_X1 c8722(
.A1(net8391),
.A2(net8920),
.ZN(net9299)
);

OAI21_X2 c8723(
.A(net9102),
.B1(net9198),
.B2(net11148),
.ZN(net9300)
);

INV_X2 c8724(
.A(net10288),
.ZN(net9301)
);

SDFF_X2 c8725(
.D(net8338),
.SE(net7287),
.SI(net9285),
.CK(clk),
.Q(net9303),
.QN(net9302)
);

NAND2_X2 c8726(
.A1(net9217),
.A2(net9214),
.ZN(net9304)
);

OAI21_X1 c8727(
.A(net9214),
.B1(net7915),
.B2(net10542),
.ZN(net9305)
);

NAND2_X4 c8728(
.A1(net8358),
.A2(net8411),
.ZN(net9306)
);

INV_X8 c8729(
.A(net9877),
.ZN(net9307)
);

AOI21_X2 c8730(
.A(net8327),
.B1(net8284),
.B2(net9307),
.ZN(net9308)
);

INV_X16 c8731(
.A(net9949),
.ZN(net9309)
);

AND2_X2 c8732(
.A1(net9290),
.A2(net9036),
.ZN(net9310)
);

XOR2_X1 c8733(
.A(net9238),
.B(net8358),
.Z(net9311)
);

AOI21_X1 c8734(
.A(net6363),
.B1(net9197),
.B2(net8871),
.ZN(net9312)
);

INV_X32 c8735(
.A(net9783),
.ZN(net9313)
);

NOR2_X1 c8736(
.A1(net6354),
.A2(net9220),
.ZN(net9314)
);

OAI33_X1 c8737(
.A1(net7405),
.A2(net8272),
.A3(net9276),
.B1(net8805),
.B2(net9224),
.B3(net9202),
.ZN(net9315)
);

AOI21_X4 c8738(
.A(net9295),
.B1(net3452),
.B2(net9290),
.ZN(net9316)
);

AND3_X1 c8739(
.A1(net9273),
.A2(net8337),
.A3(net11581),
.ZN(net9317)
);

NAND3_X1 c8740(
.A1(net9137),
.A2(net9301),
.A3(net9316),
.ZN(net9318)
);

OR2_X2 c8741(
.A1(net9292),
.A2(net9309),
.ZN(net9319)
);

NOR3_X4 c8742(
.A1(net7300),
.A2(net9226),
.A3(net9307),
.ZN(net9320)
);

NOR3_X2 c8743(
.A1(net9305),
.A2(net9138),
.A3(net8275),
.ZN(net9321)
);

AND3_X4 c8744(
.A1(net8217),
.A2(net7300),
.A3(net9264),
.ZN(net9322)
);

NAND3_X2 c8745(
.A1(net6437),
.A2(net9307),
.A3(net8927),
.ZN(net9323)
);

DFFRS_X1 c8746(
.D(net8831),
.RN(net8207),
.SN(net8217),
.CK(clk),
.Q(net9325),
.QN(net9324)
);

NOR2_X4 c8747(
.A1(net9285),
.A2(net8371),
.ZN(net9326)
);

DFFRS_X2 c8748(
.D(net9268),
.RN(net9320),
.SN(net6437),
.CK(clk),
.Q(net9328),
.QN(net9327)
);

OR3_X1 c8749(
.A1(net9264),
.A2(net9100),
.A3(net8411),
.ZN(net9329)
);

SDFF_X1 c8750(
.D(net3452),
.SE(net9313),
.SI(net9100),
.CK(clk),
.Q(net9331),
.QN(net9330)
);

MUX2_X1 c8751(
.A(net7175),
.B(net9190),
.S(net9309),
.Z(net9332)
);

OAI21_X4 c8752(
.A(net9320),
.B1(net9299),
.B2(net10957),
.ZN(net9333)
);

MUX2_X2 c8753(
.A(net9121),
.B(net9302),
.S(net9202),
.Z(net9334)
);

INV_X4 c8754(
.A(net9968),
.ZN(net9335)
);

NOR2_X2 c8755(
.A1(net9215),
.A2(net9311),
.ZN(net9336)
);

NAND3_X4 c8756(
.A1(net9325),
.A2(net9273),
.A3(net9301),
.ZN(net9337)
);

OR3_X4 c8757(
.A1(net8272),
.A2(net9294),
.A3(net9320),
.ZN(net9338)
);

SDFFS_X1 c8758(
.D(net9335),
.SE(net9336),
.SI(net7287),
.SN(net11582),
.CK(clk),
.Q(net9340),
.QN(net9339)
);

AND3_X2 c8759(
.A1(net9326),
.A2(net9188),
.A3(net11064),
.ZN(net9341)
);

INV_X1 c8760(
.A(net9782),
.ZN(net9342)
);

NOR3_X1 c8761(
.A1(net9313),
.A2(net9332),
.A3(net9319),
.ZN(net9343)
);

OAI211_X1 c8762(
.A(net9247),
.B(net9342),
.C1(net9324),
.C2(net7399),
.ZN(net9344)
);

SDFF_X2 c8763(
.D(net8284),
.SE(net9047),
.SI(net9338),
.CK(clk),
.Q(net9346),
.QN(net9345)
);

DFFRS_X1 c8764(
.D(net9011),
.RN(net9220),
.SN(net9122),
.CK(clk),
.Q(net9348),
.QN(net9347)
);

XOR2_X2 c8765(
.A(net9319),
.B(net9089),
.Z(net9349)
);

OR3_X2 c8766(
.A1(net9336),
.A2(net9343),
.A3(net7175),
.ZN(net9350)
);

OAI21_X2 c8767(
.A(net9098),
.B1(net9343),
.B2(net10981),
.ZN(net9351)
);

AOI221_X1 c8768(
.A(net9202),
.B1(net9340),
.B2(net9318),
.C1(net8983),
.C2(net8284),
.ZN(net9352)
);

OAI21_X1 c8769(
.A(net9102),
.B1(net9338),
.B2(net9340),
.ZN(net9353)
);

XNOR2_X1 c8770(
.A(net9345),
.B(net11426),
.ZN(net9354)
);

AOI21_X2 c8771(
.A(net9338),
.B1(net9330),
.B2(net8012),
.ZN(net9355)
);

OR2_X4 c8772(
.A1(net9316),
.A2(net11123),
.ZN(net9356)
);

NOR4_X4 c8773(
.A1(net7900),
.A2(net9331),
.A3(net8275),
.A4(net9339),
.ZN(net9357)
);

NOR4_X2 c8774(
.A1(net9245),
.A2(net9357),
.A3(net9339),
.A4(net10910),
.ZN(net9358)
);

OR2_X1 c8775(
.A1(net9272),
.A2(net9064),
.ZN(net9359)
);

DFFRS_X2 c8776(
.D(net9353),
.RN(net9358),
.SN(net9338),
.CK(clk),
.Q(net9361),
.QN(net9360)
);

XNOR2_X2 c8777(
.A(net9355),
.B(net9356),
.ZN(net9362)
);

AOI211_X4 c8778(
.A(net9354),
.B(net9346),
.C1(net4187),
.C2(net9356),
.ZN(net9363)
);

OAI221_X1 c8779(
.A(net9279),
.B1(net9212),
.B2(net9283),
.C1(net8109),
.C2(net9356),
.ZN(net9364)
);

AND2_X4 c8780(
.A1(net9188),
.A2(net9011),
.ZN(net9365)
);

OAI221_X4 c8781(
.A(net9337),
.B1(net9358),
.B2(net9309),
.C1(net9202),
.C2(net9339),
.ZN(net9366)
);

AOI21_X1 c8782(
.A(net9351),
.B1(net9100),
.B2(net9138),
.ZN(net9367)
);

AOI21_X4 c8783(
.A(net9346),
.B1(net9362),
.B2(net7012),
.ZN(net9368)
);

AND3_X1 c8784(
.A1(net9279),
.A2(net9340),
.A3(net11125),
.ZN(net9369)
);

NAND3_X1 c8785(
.A1(net8392),
.A2(net9363),
.A3(net6437),
.ZN(net9370)
);

NOR4_X1 c8786(
.A1(net9333),
.A2(net9369),
.A3(net9330),
.A4(net9339),
.ZN(net9371)
);

NOR3_X4 c8787(
.A1(net9331),
.A2(net9272),
.A3(net11122),
.ZN(net9372)
);

SDFF_X1 c8788(
.D(net9230),
.SE(net8927),
.SI(net9371),
.CK(clk),
.Q(net9374),
.QN(net9373)
);

AND2_X1 c8789(
.A1(net9317),
.A2(net9364),
.ZN(net9375)
);

SDFFRS_X1 c8790(
.D(net9375),
.RN(net9212),
.SE(net9342),
.SI(net9102),
.SN(net9202),
.CK(clk),
.Q(net9377),
.QN(net9376)
);

SDFF_X2 c8791(
.D(net9372),
.SE(net9358),
.SI(net11140),
.CK(clk),
.Q(net9379),
.QN(net9378)
);

NOR3_X2 c8792(
.A1(net9371),
.A2(net9369),
.A3(net11209),
.ZN(net9380)
);

AND3_X4 c8793(
.A1(net9036),
.A2(net9368),
.A3(net9369),
.ZN(net9381)
);

NAND3_X2 c8794(
.A1(net9362),
.A2(net9374),
.A3(net9356),
.ZN(net9382)
);

OR3_X1 c8795(
.A1(net9382),
.A2(net9373),
.A3(net10818),
.ZN(net9383)
);

DFFRS_X1 c8796(
.D(net9216),
.RN(net9378),
.SN(net10765),
.CK(clk),
.Q(net9385),
.QN(net9384)
);

DFFRS_X2 c8797(
.D(net9379),
.RN(net9372),
.SN(net11007),
.CK(clk),
.Q(net9387),
.QN(net9386)
);

NAND2_X1 c8798(
.A1(net8434),
.A2(net8475),
.ZN(net9388)
);

MUX2_X1 c8799(
.A(net9361),
.B(net9282),
.S(net6883),
.Z(net9389)
);

NAND2_X2 c8800(
.A1(net9098),
.A2(net11583),
.ZN(net9390)
);

NAND2_X4 c8801(
.A1(net4539),
.A2(net9184),
.ZN(net9391)
);

OAI21_X4 c8802(
.A(net9308),
.B1(net9340),
.B2(net10541),
.ZN(net9392)
);

INV_X2 c8803(
.A(net10105),
.ZN(net9393)
);

AND2_X2 c8804(
.A1(net9304),
.A2(net9344),
.ZN(net9394)
);

XOR2_X1 c8805(
.A(net9340),
.B(net11447),
.Z(net9395)
);

INV_X8 c8806(
.A(net9682),
.ZN(net9396)
);

OAI221_X2 c8807(
.A(net9391),
.B1(net8415),
.B2(net8475),
.C1(net9344),
.C2(net9189),
.ZN(net9397)
);

NOR2_X1 c8808(
.A1(net8279),
.A2(net9090),
.ZN(net9398)
);

MUX2_X2 c8809(
.A(net8238),
.B(net8871),
.S(net9360),
.Z(net9399)
);

NAND3_X4 c8810(
.A1(net9388),
.A2(net9184),
.A3(net9297),
.ZN(net9400)
);

OR3_X4 c8811(
.A1(net9392),
.A2(net9090),
.A3(net8377),
.ZN(net9401)
);

OR2_X2 c8812(
.A1(net5234),
.A2(net9389),
.ZN(net9402)
);

DFFR_X1 c8813(
.D(net9077),
.RN(net8469),
.CK(clk),
.Q(net9404),
.QN(net9403)
);

INV_X16 c8814(
.A(net11334),
.ZN(net9405)
);

AOI211_X2 c8815(
.A(net7435),
.B(net7509),
.C1(net8411),
.C2(net9400),
.ZN(net9406)
);

AOI22_X1 c8816(
.A1(net6306),
.A2(net8401),
.B1(net9327),
.B2(net8927),
.ZN(net9407)
);

SDFF_X1 c8817(
.D(net8207),
.SE(net7013),
.SI(net9400),
.CK(clk),
.Q(net9409),
.QN(net9408)
);

AND3_X2 c8818(
.A1(net7911),
.A2(net9282),
.A3(net9400),
.ZN(net9410)
);

NOR3_X1 c8819(
.A1(net8446),
.A2(out13),
.A3(net9356),
.ZN(net9411)
);

OR3_X2 c8820(
.A1(net9280),
.A2(net9198),
.A3(net9392),
.ZN(net9412)
);

OAI21_X2 c8821(
.A(net9411),
.B1(net9245),
.B2(net9322),
.ZN(net9413)
);

OAI21_X1 c8822(
.A(net9312),
.B1(net9376),
.B2(net11426),
.ZN(net9414)
);

AOI21_X2 c8823(
.A(net8469),
.B1(net9392),
.B2(net9318),
.ZN(net9415)
);

NOR2_X4 c8824(
.A1(net9407),
.A2(net9405),
.ZN(net9416)
);

AOI21_X1 c8825(
.A(net9299),
.B1(net7235),
.B2(net11577),
.ZN(net9417)
);

AOI21_X4 c8826(
.A(net9405),
.B1(net9167),
.B2(net9357),
.ZN(net9418)
);

AND3_X1 c8827(
.A1(net9321),
.A2(net9393),
.A3(net7509),
.ZN(net9419)
);

NOR2_X2 c8828(
.A1(net9184),
.A2(net9418),
.ZN(net9420)
);

XOR2_X2 c8829(
.A(net9416),
.B(net9413),
.Z(net9421)
);

XNOR2_X1 c8830(
.A(net9415),
.B(net9280),
.ZN(net9422)
);

SDFFRS_X2 c8831(
.D(net9021),
.RN(net9409),
.SE(net9090),
.SI(net8207),
.SN(net7445),
.CK(clk),
.Q(net9424),
.QN(net9423)
);

DFFR_X2 c8832(
.D(net9359),
.RN(net9398),
.CK(clk),
.Q(net9426),
.QN(net9425)
);

NAND3_X1 c8833(
.A1(net9356),
.A2(net7460),
.A3(net9166),
.ZN(net9427)
);

OR2_X4 c8834(
.A1(net9276),
.A2(net9415),
.ZN(net9428)
);

NOR3_X4 c8835(
.A1(net7509),
.A2(net10766),
.A3(net10976),
.ZN(net9429)
);

INV_X32 c8836(
.A(net10104),
.ZN(net9430)
);

SDFF_X2 c8837(
.D(net7483),
.SE(net9321),
.SI(net9021),
.CK(clk),
.Q(net9432),
.QN(net9431)
);

NOR3_X2 c8838(
.A1(net9426),
.A2(net9392),
.A3(net8468),
.ZN(net9433)
);

DFFS_X1 c8839(
.D(net7509),
.SN(net9422),
.CK(clk),
.Q(net9435),
.QN(net9434)
);

OR2_X1 c8840(
.A1(net8871),
.A2(net9420),
.ZN(net9436)
);

AND3_X4 c8841(
.A1(net8468),
.A2(net8983),
.A3(net8400),
.ZN(net9437)
);

NAND3_X2 c8842(
.A1(net9427),
.A2(net7399),
.A3(net11576),
.ZN(net9438)
);

XNOR2_X2 c8843(
.A(net8431),
.B(net9430),
.ZN(net9439)
);

INV_X4 c8844(
.A(net10172),
.ZN(net9440)
);

OR3_X1 c8845(
.A1(net7399),
.A2(out13),
.A3(net11203),
.ZN(net9441)
);

MUX2_X1 c8846(
.A(net9390),
.B(net9432),
.S(net11258),
.Z(net9442)
);

INV_X1 c8847(
.A(net9821),
.ZN(net9443)
);

OAI21_X4 c8848(
.A(net9303),
.B1(net9412),
.B2(net9423),
.ZN(net9444)
);

MUX2_X2 c8849(
.A(net8464),
.B(net9441),
.S(net9344),
.Z(net9445)
);

NAND3_X4 c8850(
.A1(net9394),
.A2(net7482),
.A3(net10722),
.ZN(net9446)
);

OR3_X4 c8851(
.A1(net8475),
.A2(net9408),
.A3(net9311),
.ZN(net9447)
);

AND3_X2 c8852(
.A1(net9322),
.A2(net9280),
.A3(net9423),
.ZN(net9448)
);

AND2_X4 c8853(
.A1(net9410),
.A2(net9090),
.ZN(net9449)
);

NOR3_X1 c8854(
.A1(net9438),
.A2(net7452),
.A3(net8871),
.ZN(net9450)
);

OR3_X2 c8855(
.A1(net9240),
.A2(net9318),
.A3(net9312),
.ZN(net9451)
);

OAI21_X2 c8856(
.A(net9415),
.B1(net8238),
.B2(net10516),
.ZN(net9452)
);

OAI21_X1 c8857(
.A(net9413),
.B1(net9431),
.B2(net10958),
.ZN(net9453)
);

AND2_X1 c8858(
.A1(net8411),
.A2(net9320),
.ZN(net9454)
);

AOI21_X2 c8859(
.A(net8109),
.B1(net9448),
.B2(net9389),
.ZN(net9455)
);

DFFRS_X1 c8860(
.D(net9443),
.RN(net9428),
.SN(net9412),
.CK(clk),
.Q(net9457),
.QN(net9456)
);

NAND2_X1 c8861(
.A1(net9436),
.A2(net9457),
.ZN(net9458)
);

AOI21_X1 c8862(
.A(net9449),
.B1(net9448),
.B2(net11583),
.ZN(net9459)
);

INV_X2 c8863(
.A(net9681),
.ZN(net9460)
);

AOI21_X4 c8864(
.A(net9442),
.B1(net9458),
.B2(net9403),
.ZN(net9461)
);

AND3_X1 c8865(
.A1(net9461),
.A2(net9458),
.A3(net9425),
.ZN(net9462)
);

NAND3_X1 c8866(
.A1(net9431),
.A2(net10720),
.A3(net11180),
.ZN(net9463)
);

AOI222_X2 c8867(
.A1(net9417),
.A2(net9413),
.B1(net9189),
.B2(net9444),
.C1(net8415),
.C2(net9456),
.ZN(net9464)
);

NOR3_X4 c8868(
.A1(net8421),
.A2(net9462),
.A3(net9460),
.ZN(net9465)
);

NOR3_X2 c8869(
.A1(net9465),
.A2(net9460),
.A3(net11066),
.ZN(net9466)
);

AND3_X4 c8870(
.A1(net9447),
.A2(net9441),
.A3(net8468),
.ZN(net9467)
);

NAND3_X2 c8871(
.A1(net8372),
.A2(net9430),
.A3(net9465),
.ZN(net9468)
);

NAND2_X2 c8872(
.A1(net9460),
.A2(net11242),
.ZN(net9469)
);

OR3_X1 c8873(
.A1(net7414),
.A2(net9395),
.A3(net9307),
.ZN(net9470)
);

NAND2_X4 c8874(
.A1(net9377),
.A2(net9307),
.ZN(net9471)
);

OAI222_X1 c8875(
.A1(net9470),
.A2(net9471),
.B1(net9181),
.B2(net9444),
.C1(net9465),
.C2(net11582),
.ZN(net9472)
);

MUX2_X1 c8876(
.A(net9434),
.B(net10955),
.S(net11153),
.Z(net9473)
);

OAI21_X4 c8877(
.A(net9473),
.B1(net9281),
.B2(net11257),
.ZN(net9474)
);

MUX2_X2 c8878(
.A(net9469),
.B(net11195),
.S(net11584),
.Z(net9475)
);

NAND3_X4 c8879(
.A1(net9474),
.A2(net9475),
.A3(net9224),
.ZN(net9476)
);

AOI221_X4 c8880(
.A(net9445),
.B1(net9438),
.B2(net9476),
.C1(net6472),
.C2(net11585),
.ZN(net9477)
);

AND2_X2 c8881(
.A1(net8805),
.A2(net9435),
.ZN(net9478)
);

OR3_X4 c8882(
.A1(net9460),
.A2(net9287),
.A3(net9440),
.ZN(net9479)
);

AND4_X4 c8883(
.A1(net8498),
.A2(net8328),
.A3(net8594),
.A4(net9123),
.ZN(net9480)
);

AND3_X2 c8884(
.A1(net9452),
.A2(net9312),
.A3(net9123),
.ZN(net9481)
);

AOI221_X2 c8885(
.A(net9298),
.B1(net9428),
.B2(net6472),
.C1(net9400),
.C2(net9460),
.ZN(net9482)
);

NOR3_X1 c8886(
.A1(net7460),
.A2(net7414),
.A3(net7519),
.ZN(net9483)
);

XOR2_X1 c8887(
.A(net9429),
.B(net11396),
.Z(net9484)
);

NOR2_X1 c8888(
.A1(net9446),
.A2(net7561),
.ZN(net9485)
);

DFFRS_X2 c8889(
.D(net9249),
.RN(net10817),
.SN(net11254),
.CK(clk),
.Q(net9487),
.QN(net9486)
);

OR2_X2 c8890(
.A1(net7211),
.A2(net9484),
.ZN(net9488)
);

OR3_X2 c8891(
.A1(net7235),
.A2(net9400),
.A3(net9310),
.ZN(net9489)
);

INV_X8 c8892(
.A(net9684),
.ZN(net9490)
);

SDFF_X1 c8893(
.D(net9349),
.SE(net9465),
.SI(net11135),
.CK(clk),
.Q(net9492),
.QN(net9491)
);

SDFF_X2 c8894(
.D(net8983),
.SE(net9344),
.SI(net11395),
.CK(clk),
.Q(net9494),
.QN(net9493)
);

OAI21_X2 c8895(
.A(net9328),
.B1(net9494),
.B2(net11425),
.ZN(net9495)
);

NOR2_X4 c8896(
.A1(net6469),
.A2(net9460),
.ZN(net9496)
);

OAI21_X1 c8897(
.A(net7445),
.B1(net9387),
.B2(net9281),
.ZN(net9497)
);

NOR2_X2 c8898(
.A1(net9484),
.A2(net11448),
.ZN(net9498)
);

AOI21_X2 c8899(
.A(net5601),
.B1(net9484),
.B2(net9344),
.ZN(net9499)
);

INV_X16 c8900(
.A(net9962),
.ZN(net9500)
);

XOR2_X2 c8901(
.A(net9480),
.B(net9484),
.Z(net9501)
);

AOI21_X1 c8902(
.A(net9312),
.B1(net8353),
.B2(net9500),
.ZN(net9502)
);

XNOR2_X1 c8903(
.A(net9123),
.B(net8418),
.ZN(net9503)
);

OR2_X4 c8904(
.A1(net7452),
.A2(net7460),
.ZN(net9504)
);

AOI21_X4 c8905(
.A(net7544),
.B1(net9490),
.B2(net9460),
.ZN(net9505)
);

INV_X32 c8906(
.A(net9683),
.ZN(net9506)
);

NAND4_X1 c8907(
.A1(net9505),
.A2(net9190),
.A3(net8511),
.A4(net9491),
.ZN(net9507)
);

AND3_X1 c8908(
.A1(net9424),
.A2(net9446),
.A3(net9297),
.ZN(net9508)
);

OR4_X1 c8909(
.A1(net9369),
.A2(net9487),
.A3(net8592),
.A4(net8927),
.ZN(net9509)
);

NAND3_X1 c8910(
.A1(net4598),
.A2(net8235),
.A3(net8511),
.ZN(net9510)
);

NOR3_X4 c8911(
.A1(net9440),
.A2(net9484),
.A3(net9486),
.ZN(net9511)
);

NOR3_X2 c8912(
.A1(net8511),
.A2(net9509),
.A3(net9505),
.ZN(net9512)
);

AND3_X4 c8913(
.A1(net9506),
.A2(net1730),
.A3(net10913),
.ZN(net9513)
);

OAI22_X1 c8914(
.A1(net5584),
.A2(net9404),
.B1(net8805),
.B2(net11142),
.ZN(net9514)
);

NAND3_X2 c8915(
.A1(net9432),
.A2(net9500),
.A3(net9123),
.ZN(net9515)
);

OR3_X1 c8916(
.A1(net9506),
.A2(net9181),
.A3(net9485),
.ZN(net9516)
);

MUX2_X1 c8917(
.A(net9298),
.B(net7445),
.S(net11395),
.Z(net9517)
);

OR2_X1 c8918(
.A1(net9515),
.A2(net10600),
.ZN(net9518)
);

OAI21_X4 c8919(
.A(net9500),
.B1(net7445),
.B2(net11463),
.ZN(net9519)
);

MUX2_X2 c8920(
.A(net9397),
.B(net9503),
.S(net8920),
.Z(net9520)
);

NAND3_X4 c8921(
.A1(net7607),
.A2(net9344),
.A3(net3615),
.ZN(net9521)
);

OR3_X4 c8922(
.A1(net9516),
.A2(net9517),
.A3(net9431),
.ZN(net9522)
);

AND3_X2 c8923(
.A1(net9521),
.A2(net9167),
.A3(net9357),
.ZN(net9523)
);

NOR3_X1 c8924(
.A1(net9435),
.A2(net8589),
.A3(net9492),
.ZN(net9524)
);

OR3_X2 c8925(
.A1(net9485),
.A2(net8519),
.A3(net11581),
.ZN(net9525)
);

OAI21_X2 c8926(
.A(net9181),
.B1(net9522),
.B2(net9347),
.ZN(net9526)
);

OAI21_X1 c8927(
.A(net8353),
.B1(net8511),
.B2(net10988),
.ZN(net9527)
);

AOI21_X2 c8928(
.A(net8538),
.B1(net8012),
.B2(net9514),
.ZN(net9528)
);

AOI21_X1 c8929(
.A(net7558),
.B1(net9476),
.B2(net9397),
.ZN(net9529)
);

SDFFS_X2 c8930(
.D(net9501),
.SE(net9498),
.SI(net9282),
.SN(net9529),
.CK(clk),
.Q(net9531),
.QN(net9530)
);

DFFRS_X1 c8931(
.D(net9508),
.RN(net9507),
.SN(net9514),
.CK(clk),
.Q(net9533),
.QN(net9532)
);

AOI21_X4 c8932(
.A(net9511),
.B1(net9527),
.B2(net9369),
.ZN(net9534)
);

AND3_X1 c8933(
.A1(net9528),
.A2(net9499),
.A3(net9444),
.ZN(net9535)
);

NAND3_X1 c8934(
.A1(net9463),
.A2(net9530),
.A3(net11463),
.ZN(net9536)
);

NOR3_X4 c8935(
.A1(net8418),
.A2(net9432),
.A3(net11342),
.ZN(net9537)
);

NOR3_X2 c8936(
.A1(net9429),
.A2(net9500),
.A3(net9369),
.ZN(net9538)
);

AND3_X4 c8937(
.A1(net7562),
.A2(net9533),
.A3(net9531),
.ZN(net9539)
);

XNOR2_X2 c8938(
.A(net8448),
.B(net9519),
.ZN(net9540)
);

NAND3_X2 c8939(
.A1(net9527),
.A2(net9496),
.A3(net9529),
.ZN(net9541)
);

AND2_X4 c8940(
.A1(net9504),
.A2(net9282),
.ZN(net9542)
);

OR3_X1 c8941(
.A1(net9520),
.A2(net9518),
.A3(net9446),
.ZN(net9543)
);

MUX2_X1 c8942(
.A(net9540),
.B(net9531),
.S(net9529),
.Z(net9544)
);

OAI21_X4 c8943(
.A(net6472),
.B1(net7544),
.B2(net9434),
.ZN(net9545)
);

MUX2_X2 c8944(
.A(net3615),
.B(net5584),
.S(net9522),
.Z(net9546)
);

NAND3_X4 c8945(
.A1(net9542),
.A2(net9524),
.A3(net8509),
.ZN(net9547)
);

OR3_X4 c8946(
.A1(net9523),
.A2(net7563),
.A3(net3626),
.ZN(net9548)
);

INV_X4 c8947(
.A(net9820),
.ZN(net9549)
);

AND3_X2 c8948(
.A1(net9539),
.A2(net9465),
.A3(net11396),
.ZN(net9550)
);

NOR3_X1 c8949(
.A1(net9245),
.A2(net9349),
.A3(net8520),
.ZN(net9551)
);

OR3_X2 c8950(
.A1(net9545),
.A2(net9513),
.A3(net9514),
.ZN(net9552)
);

OAI21_X2 c8951(
.A(net9522),
.B1(net9493),
.B2(net11427),
.ZN(net9553)
);

OAI21_X1 c8952(
.A(net9553),
.B1(net9485),
.B2(net11210),
.ZN(net9554)
);

OAI222_X4 c8953(
.A1(net9497),
.A2(net9546),
.B1(net9522),
.B2(net8519),
.C1(net7445),
.C2(net9396),
.ZN(net9555)
);

AOI21_X2 c8954(
.A(net9404),
.B1(net9526),
.B2(net9522),
.ZN(net9556)
);

AOI221_X1 c8955(
.A(net9525),
.B1(net8520),
.B2(net9529),
.C1(net7445),
.C2(net11587),
.ZN(net9557)
);

AOI21_X1 c8956(
.A(net9548),
.B1(net7445),
.B2(net11229),
.ZN(net9558)
);

AOI21_X4 c8957(
.A(net9536),
.B1(net9552),
.B2(net9424),
.ZN(net9559)
);

AND3_X1 c8958(
.A1(net8415),
.A2(net9551),
.A3(net11586),
.ZN(net9560)
);

NAND3_X1 c8959(
.A1(net9523),
.A2(net11260),
.A3(net11580),
.ZN(net9561)
);

OAI222_X2 c8960(
.A1(net9548),
.A2(net9540),
.B1(net9561),
.B2(net9514),
.C1(net9506),
.C2(net11235),
.ZN(net9562)
);

NOR3_X4 c8961(
.A1(net8534),
.A2(net9559),
.A3(net9532),
.ZN(net9563)
);

NOR3_X2 c8962(
.A1(net9538),
.A2(net9561),
.A3(net10962),
.ZN(net9564)
);

OAI221_X1 c8963(
.A(net9485),
.B1(net9561),
.B2(net9529),
.C1(net11218),
.C2(net11427),
.ZN(net9565)
);

AND3_X4 c8964(
.A1(net9465),
.A2(net7211),
.A3(net9493),
.ZN(net9566)
);

NAND3_X2 c8965(
.A1(net8328),
.A2(net8634),
.A3(net8927),
.ZN(net9567)
);

AND2_X1 c8966(
.A1(net7577),
.A2(net8322),
.ZN(net9568)
);

OR3_X1 c8967(
.A1(net7359),
.A2(net9494),
.A3(net9529),
.ZN(net9569)
);

NAND2_X1 c8968(
.A1(net9402),
.A2(net8600),
.ZN(net9570)
);

INV_X1 c8969(
.A(net9686),
.ZN(net9571)
);

MUX2_X1 c8970(
.A(net9568),
.B(net6559),
.S(net9514),
.Z(net9572)
);

DFFRS_X2 c8971(
.D(net8927),
.RN(net8634),
.SN(net10599),
.CK(clk),
.Q(net9574),
.QN(net9573)
);

OAI21_X4 c8972(
.A(net9384),
.B1(net9495),
.B2(net10989),
.ZN(net9575)
);

NAND2_X2 c8973(
.A1(net2777),
.A2(net11136),
.ZN(net9576)
);

MUX2_X2 c8974(
.A(net9348),
.B(net7519),
.S(net8322),
.Z(net9577)
);

NAND3_X4 c8975(
.A1(net9570),
.A2(net7649),
.A3(net9492),
.ZN(net9578)
);

NAND2_X4 c8976(
.A1(net8594),
.A2(net11577),
.ZN(net9579)
);

AND2_X2 c8977(
.A1(net8646),
.A2(net11143),
.ZN(net9580)
);

OR3_X4 c8978(
.A1(net9444),
.A2(net11126),
.A3(net11563),
.ZN(net9581)
);

AND3_X2 c8979(
.A1(net8518),
.A2(net9429),
.A3(net9444),
.ZN(net9582)
);

INV_X2 c8980(
.A(net9685),
.ZN(net9583)
);

NOR3_X1 c8981(
.A1(net8600),
.A2(net8686),
.A3(net9574),
.ZN(net9584)
);

OR3_X2 c8982(
.A1(net8440),
.A2(net9357),
.A3(net9529),
.ZN(net9585)
);

OAI21_X2 c8983(
.A(net9357),
.B1(net8279),
.B2(net9491),
.ZN(net9586)
);

OAI21_X1 c8984(
.A(net8667),
.B1(net9478),
.B2(net9439),
.ZN(net9587)
);

AOI21_X2 c8985(
.A(net8675),
.B1(net9498),
.B2(net11000),
.ZN(net9588)
);

XOR2_X1 c8986(
.A(net9444),
.B(net9588),
.Z(net9589)
);

AND4_X2 c8987(
.A1(net9307),
.A2(net9465),
.A3(net9478),
.A4(net8627),
.ZN(net9590)
);

NOR2_X1 c8988(
.A1(net8594),
.A2(net11263),
.ZN(net9591)
);

AOI21_X1 c8989(
.A(net7684),
.B1(net8682),
.B2(net10999),
.ZN(net9592)
);

AOI21_X4 c8990(
.A(net8615),
.B1(net9574),
.B2(net9583),
.ZN(net9593)
);

SDFF_X1 c8991(
.D(net3626),
.SE(net8634),
.SI(net9583),
.CK(clk),
.Q(net9595),
.QN(net9594)
);

AND3_X1 c8992(
.A1(net6495),
.A2(net9478),
.A3(net11219),
.ZN(net9596)
);

NAND3_X1 c8993(
.A1(net6636),
.A2(net9592),
.A3(net9594),
.ZN(net9597)
);

NOR3_X4 c8994(
.A1(net8920),
.A2(net9586),
.A3(net8628),
.ZN(net9598)
);

NOR3_X2 c8995(
.A1(net9578),
.A2(net9573),
.A3(net11291),
.ZN(net9599)
);

AND3_X4 c8996(
.A1(net9310),
.A2(net9444),
.A3(net11387),
.ZN(net9600)
);

AND4_X1 c8997(
.A1(net9529),
.A2(net8681),
.A3(net9573),
.A4(net7519),
.ZN(net9601)
);

NAND3_X2 c8998(
.A1(net8509),
.A2(net9579),
.A3(net8628),
.ZN(net9602)
);

OR3_X1 c8999(
.A1(net9476),
.A2(net8440),
.A3(net10690),
.ZN(net9603)
);

MUX2_X1 c9000(
.A(net9598),
.B(net9492),
.S(net9439),
.Z(net9604)
);

OAI21_X4 c9001(
.A(net9275),
.B1(net9580),
.B2(net9357),
.ZN(net9605)
);

MUX2_X2 c9002(
.A(net8593),
.B(net9498),
.S(net10994),
.Z(net9606)
);

NAND3_X4 c9003(
.A1(net9400),
.A2(net9596),
.A3(net6559),
.ZN(net9607)
);

INV_X8 c9004(
.A(net9886),
.ZN(net9608)
);

INV_X16 c9005(
.A(net9887),
.ZN(net9609)
);

OR2_X2 c9006(
.A1(net9591),
.A2(net10871),
.ZN(net9610)
);

OR3_X4 c9007(
.A1(net9602),
.A2(net9575),
.A3(net8440),
.ZN(net9611)
);

AND3_X2 c9008(
.A1(net9595),
.A2(net9583),
.A3(net11425),
.ZN(net9612)
);

NOR3_X1 c9009(
.A1(net8430),
.A2(net9609),
.A3(net9611),
.ZN(net9613)
);

OR3_X2 c9010(
.A1(net9584),
.A2(net9613),
.A3(net9610),
.ZN(net9614)
);

OAI21_X2 c9011(
.A(net9478),
.B1(net9608),
.B2(net11316),
.ZN(net9615)
);

OAI21_X1 c9012(
.A(net9604),
.B1(net9615),
.B2(net11144),
.ZN(net9616)
);

AOI21_X2 c9013(
.A(net6675),
.B1(net8682),
.B2(net9492),
.ZN(net9617)
);

AOI21_X1 c9014(
.A(net8520),
.B1(net9385),
.B2(net9595),
.ZN(net9618)
);

AOI21_X4 c9015(
.A(net9595),
.B1(net10602),
.B2(net11292),
.ZN(net9619)
);

AOI222_X1 c9016(
.A1(net9593),
.A2(net9610),
.B1(net9608),
.B2(net9618),
.C1(net9594),
.C2(net9491),
.ZN(net9620)
);

AND3_X1 c9017(
.A1(net9571),
.A2(net9576),
.A3(net8509),
.ZN(net9621)
);

NAND3_X1 c9018(
.A1(net9581),
.A2(net9616),
.A3(net9606),
.ZN(net9622)
);

NOR3_X4 c9019(
.A1(net9412),
.A2(net9615),
.A3(net9602),
.ZN(net9623)
);

NOR3_X2 c9020(
.A1(net9618),
.A2(net9587),
.A3(net9610),
.ZN(net9624)
);

AOI222_X4 c9021(
.A1(net5623),
.A2(net9623),
.B1(net9610),
.B2(net9618),
.C1(net8279),
.C2(net9594),
.ZN(net9625)
);

AND3_X4 c9022(
.A1(net8612),
.A2(net9396),
.A3(net9606),
.ZN(net9626)
);

NAND3_X2 c9023(
.A1(net7672),
.A2(net9439),
.A3(net9618),
.ZN(net9627)
);

AOI22_X4 c9024(
.A1(net9620),
.A2(net9514),
.B1(net9616),
.B2(net9618),
.ZN(net9628)
);

OR3_X1 c9025(
.A1(net9419),
.A2(net9612),
.A3(net9618),
.ZN(net9629)
);

MUX2_X1 c9026(
.A(net7649),
.B(net9621),
.S(net9625),
.Z(net9630)
);

OAI21_X4 c9027(
.A(net9583),
.B1(net9622),
.B2(net9606),
.ZN(net9631)
);

MUX2_X2 c9028(
.A(net9627),
.B(net9597),
.S(net9603),
.Z(net9632)
);

NAND3_X4 c9029(
.A1(net9589),
.A2(net9631),
.A3(net9629),
.ZN(net9633)
);

OR3_X4 c9030(
.A1(net9614),
.A2(net9595),
.A3(net10718),
.ZN(net9634)
);

AND3_X2 c9031(
.A1(net9619),
.A2(net9629),
.A3(net11324),
.ZN(net9635)
);

OAI33_X1 c9032(
.A1(net9624),
.A2(net9549),
.A3(net9629),
.B1(net9491),
.B2(net8627),
.B3(net9618),
.ZN(net9636)
);

NOR3_X1 c9033(
.A1(net9495),
.A2(net9636),
.A3(net11325),
.ZN(net9637)
);

OR3_X2 c9034(
.A1(net9561),
.A2(net9629),
.A3(net9626),
.ZN(net9638)
);

OAI21_X2 c9035(
.A(net9628),
.B1(net9494),
.B2(net9637),
.ZN(net9639)
);

OAI21_X1 c9036(
.A(net9498),
.B1(net10689),
.B2(net11315),
.ZN(net9640)
);

AOI21_X2 c9037(
.A(net9630),
.B1(net9618),
.B2(net11098),
.ZN(net9641)
);

AOI21_X1 c9038(
.A(net9637),
.B1(net9641),
.B2(net9640),
.ZN(net9642)
);

OAI22_X4 c9039(
.A1(net8322),
.A2(net9635),
.B1(net10601),
.B2(net11328)
);

SDFFR_X1 merge9040(
.D(net5156),
.RN(net6199),
.SE(net6201),
.SI(net6030),
.CK(clk),
.Q(net9644),
.QN(net9643)
);

INV_X32 merge9041(
.A(net10078),
.ZN(net9645)
);

SDFF_X2 merge9042(
.D(net1806),
.SE(net1681),
.SI(net1782),
.CK(clk),
.Q(net9647),
.QN(net9646)
);

DFFRS_X1 merge9043(
.D(net4907),
.RN(net3904),
.SN(net3936),
.CK(clk),
.Q(net9649),
.QN(net9648)
);

DFFS_X2 merge9044(
.D(net888),
.SN(net864),
.CK(clk),
.Q(net9651),
.QN(net9650)
);

DFFR_X1 merge9045(
.D(net421),
.RN(net153),
.CK(clk),
.Q(net9653),
.QN(net9652)
);

DFFR_X2 merge9046(
.D(net6939),
.RN(net7870),
.CK(clk),
.Q(net9655),
.QN(net9654)
);

NOR2_X4 merge9047(
.A1(net1535),
.A2(net1542),
.ZN(net9656)
);

SDFFR_X2 merge9048(
.D(net2876),
.RN(net3418),
.SE(net3832),
.SI(net3821),
.CK(clk),
.Q(net9658),
.QN(net9657)
);

SDFFS_X1 merge9049(
.D(net7447),
.SE(net5383),
.SI(net7602),
.SN(net11562),
.CK(clk),
.Q(net9660),
.QN(net9659)
);

DFFRS_X2 merge9050(
.D(net2923),
.RN(net2929),
.SN(net1968),
.CK(clk),
.Q(net9662),
.QN(net9661)
);

DFFS_X1 merge9051(
.D(net3246),
.SN(net3172),
.CK(clk),
.Q(net9664),
.QN(net9663)
);

INV_X4 merge9052(
.A(net10019),
.ZN(net9665)
);

AOI22_X2 merge9053(
.A1(net6616),
.A2(net8378),
.B1(net8542),
.B2(net8561),
.ZN(net9666)
);

DFFS_X2 merge9054(
.D(net88),
.SN(net527),
.CK(clk),
.Q(net9668),
.QN(net9667)
);

SDFFS_X2 merge9055(
.D(net5383),
.SE(net6548),
.SI(net5676),
.SN(net5694),
.CK(clk),
.Q(net9670),
.QN(net9669)
);

NAND4_X4 merge9056(
.A1(net5525),
.A2(net5567),
.A3(net5610),
.A4(net5637),
.ZN(net9671)
);

INV_X1 merge9057(
.A(net9917),
.ZN(net9672)
);

INV_X2 merge9058(
.A(net10381),
.ZN(net9673)
);

INV_X8 merge9059(
.A(net11175),
.ZN(net9674)
);

DFFR_X1 merge9060(
.D(net1094),
.RN(net1065),
.CK(clk),
.Q(net9676),
.QN(net9675)
);

SDFFR_X1 merge9061(
.D(net8151),
.RN(net8156),
.SE(net8172),
.SI(net8215),
.CK(clk),
.Q(net9678),
.QN(net9677)
);

DFFR_X2 merge9062(
.D(net1944),
.RN(net3005),
.CK(clk),
.Q(net9680),
.QN(net9679)
);

SDFFR_X2 merge9063(
.D(net9311),
.RN(net9223),
.SE(net9448),
.SI(net10863),
.CK(clk),
.Q(net9682),
.QN(net9681)
);

SDFFS_X1 merge9064(
.D(net7597),
.SE(net9485),
.SI(net9386),
.SN(net9488),
.CK(clk),
.Q(net9684),
.QN(net9683)
);

SDFFS_X2 merge9065(
.D(net8627),
.SE(net9529),
.SI(net9582),
.SN(net9249),
.CK(clk),
.Q(net9686),
.QN(net9685)
);

NOR2_X2 merge9066(
.A1(net8416),
.A2(net7812),
.ZN(net9687)
);

SDFFR_X1 merge9067(
.D(net8313),
.RN(net8260),
.SE(net8339),
.SI(net8405),
.CK(clk),
.Q(net9689),
.QN(net9688)
);

INV_X16 merge9068(
.A(net10136),
.ZN(net9690)
);

DFFS_X1 merge9069(
.D(net6891),
.SN(net5028),
.CK(clk),
.Q(net9692),
.QN(net9691)
);

SDFFR_X2 merge9070(
.D(net8907),
.RN(net8955),
.SE(net8975),
.SI(net8889),
.CK(clk),
.Q(net9694),
.QN(net9693)
);

AOI21_X4 merge9071(
.A(net3189),
.B1(net2987),
.B2(net3167),
.ZN(net9695)
);

INV_X32 merge9072(
.A(net10289),
.ZN(net9696)
);

AND3_X1 merge9073(
.A1(net560),
.A2(net1545),
.A3(net2241),
.ZN(net9697)
);

NAND3_X1 merge9074(
.A1(net4506),
.A2(net4500),
.A3(net10744),
.ZN(net9698)
);

INV_X4 merge9075(
.A(net10110),
.ZN(net9699)
);

DFFS_X2 merge9076(
.D(net215),
.SN(net192),
.CK(clk),
.Q(net9701),
.QN(net9700)
);

INV_X1 merge9077(
.A(net10036),
.ZN(net9702)
);

XOR2_X2 merge9078(
.A(net3503),
.B(net3612),
.Z(net9703)
);

NOR3_X4 merge9079(
.A1(net3352),
.A2(net4210),
.A3(net10885),
.ZN(net9704)
);

DFFR_X1 merge9080(
.D(net855),
.RN(net772),
.CK(clk),
.Q(net9706),
.QN(net9705)
);

OAI211_X2 merge9081(
.A(net9031),
.B(net9021),
.C1(net8016),
.C2(net9152),
.ZN(net9707)
);

SDFFRS_X1 merge9082(
.D(net6765),
.RN(net6782),
.SE(net7269),
.SI(net7742),
.SN(net6533),
.CK(clk),
.Q(net9709),
.QN(net9708)
);

SDFFS_X1 merge9083(
.D(net3836),
.SE(net2848),
.SI(net3816),
.SN(net1868),
.CK(clk),
.Q(net9711),
.QN(net9710)
);

OR4_X2 merge9084(
.A1(net8986),
.A2(net8991),
.A3(net8925),
.A4(net8830),
.ZN(net9712)
);

INV_X2 merge9085(
.A(net9990),
.ZN(net9713)
);

INV_X8 merge9086(
.A(net11302),
.ZN(net9714)
);

SDFF_X1 merge9087(
.D(net6808),
.SE(net4404),
.SI(net6364),
.CK(clk),
.Q(net9716),
.QN(net9715)
);

DFFR_X2 merge9088(
.D(net1024),
.RN(net1119),
.CK(clk),
.Q(net9718),
.QN(net9717)
);

INV_X16 merge9089(
.A(net10013),
.ZN(net9719)
);

XNOR2_X1 merge9090(
.A(net220),
.B(net1140),
.ZN(net9720)
);

DFFS_X1 merge9091(
.D(net3371),
.SN(net4361),
.CK(clk),
.Q(net9722),
.QN(net9721)
);

INV_X32 merge9092(
.A(net11471),
.ZN(net9723)
);

OR2_X4 merge9093(
.A1(net1306),
.A2(net1455),
.ZN(net9724)
);

AOI222_X2 merge9094(
.A1(net8672),
.A2(net8622),
.B1(net8732),
.B2(net7641),
.C1(net8718),
.C2(net6732),
.ZN(net9725)
);

SDFFS_X2 merge9095(
.D(net8601),
.SE(net5545),
.SI(net8625),
.SN(net11389),
.CK(clk),
.Q(net9727),
.QN(net9726)
);

AOI211_X1 merge9096(
.A(net4520),
.B(net4736),
.C1(net4737),
.C2(net11439),
.ZN(net9728)
);

DFFS_X2 merge9097(
.D(net3974),
.SN(net3988),
.CK(clk),
.Q(net9730),
.QN(net9729)
);

INV_X4 merge9098(
.A(net9809),
.ZN(net9731)
);

DFFR_X1 merge9099(
.D(net1393),
.RN(net465),
.CK(clk),
.Q(net9733),
.QN(net9732)
);

INV_X1 merge9100(
.A(net10354),
.ZN(net9734)
);

OR2_X1 merge9101(
.A1(net514),
.A2(net680),
.ZN(net9735)
);

DFFR_X2 merge9102(
.D(net5900),
.RN(net5914),
.CK(clk),
.Q(net9737),
.QN(net9736)
);

DFFS_X1 merge9103(
.D(net7795),
.SN(net7814),
.CK(clk),
.Q(net9739),
.QN(net9738)
);

INV_X2 merge9104(
.A(net11106),
.ZN(net9740)
);

INV_X8 merge9105(
.A(net10177),
.ZN(net9741)
);

INV_X16 merge9106(
.A(net10200),
.ZN(net9742)
);

SDFF_X2 merge9107(
.D(net8215),
.SE(net6104),
.SI(net8303),
.CK(clk),
.Q(net9744),
.QN(net9743)
);

INV_X32 merge9108(
.A(net10117),
.ZN(net9745)
);

NAND4_X2 merge9109(
.A1(net5583),
.A2(net4755),
.A3(net5738),
.A4(net5736),
.ZN(net9746)
);

INV_X4 merge9110(
.A(net10396),
.ZN(net9747)
);

XNOR2_X2 merge9111(
.A(net220),
.B(net354),
.ZN(net9748)
);

DFFRS_X1 merge9112(
.D(net6365),
.RN(net6277),
.SN(net6476),
.CK(clk),
.Q(net9750),
.QN(net9749)
);

DFFRS_X2 merge9113(
.D(net3426),
.RN(net3413),
.SN(net11370),
.CK(clk),
.Q(net9752),
.QN(net9751)
);

OR4_X4 merge9114(
.A1(net7103),
.A2(net7796),
.A3(net8123),
.A4(net8135),
.ZN(net9753)
);

INV_X1 merge9115(
.A(net10193),
.ZN(net9754)
);

SDFFR_X1 merge9116(
.D(net1768),
.RN(net1880),
.SE(net1904),
.SI(net2866),
.CK(clk),
.Q(net9756),
.QN(net9755)
);

DFFS_X2 merge9117(
.D(net5836),
.SN(net5940),
.CK(clk),
.Q(net9758),
.QN(net9757)
);

SDFFR_X2 merge9118(
.D(net3846),
.RN(net5744),
.SE(net5789),
.SI(net5658),
.CK(clk),
.Q(net9760),
.QN(net9759)
);

DFFR_X1 merge9119(
.D(net2990),
.RN(net1944),
.CK(clk),
.Q(net9762),
.QN(net9761)
);

SDFFS_X1 merge9120(
.D(net4067),
.SE(net5170),
.SI(net5168),
.SN(net5126),
.CK(clk),
.Q(net9764),
.QN(net9763)
);

OAI22_X2 merge9121(
.A1(net1658),
.A2(net1525),
.B1(net1663),
.B2(net1667),
.ZN(net9765)
);

SDFF_X1 merge9122(
.D(net6640),
.SE(net5652),
.SI(net3775),
.CK(clk),
.Q(net9767),
.QN(net9766)
);

AND2_X4 merge9123(
.A1(net1959),
.A2(net1036),
.ZN(net9768)
);

INV_X2 merge9124(
.A(net10318),
.ZN(net9769)
);

INV_X8 merge9125(
.A(net10059),
.ZN(net9770)
);

INV_X16 merge9126(
.A(net9811),
.ZN(net9771)
);

DFFR_X2 merge9127(
.D(net490),
.RN(net491),
.CK(clk),
.Q(net9773),
.QN(net9772)
);

DFFS_X1 merge9128(
.D(net7804),
.SN(net6870),
.CK(clk),
.Q(net9775),
.QN(net9774)
);

INV_X32 merge9129(
.A(net10380),
.ZN(net9776)
);

OAI211_X4 merge9130(
.A(net8243),
.B(net9188),
.C1(net9094),
.C2(net8012),
.ZN(net9777)
);

INV_X4 merge9131(
.A(net10239),
.ZN(net9778)
);

INV_X1 merge9132(
.A(net10192),
.ZN(net9779)
);

SDFFS_X2 merge9133(
.D(net7339),
.SE(net7345),
.SI(net6453),
.SN(net7135),
.CK(clk),
.Q(net9781),
.QN(net9780)
);

SDFFR_X1 merge9134(
.D(net8377),
.RN(net9264),
.SE(net9314),
.SI(net8391),
.CK(clk),
.Q(net9783),
.QN(net9782)
);

NOR3_X2 merge9135(
.A1(net4130),
.A2(net4227),
.A3(net4065),
.ZN(net9784)
);

INV_X2 merge9136(
.A(net9812),
.ZN(net9785)
);

OAI211_X1 merge9137(
.A(net489),
.B(net4367),
.C1(net4473),
.C2(net3518),
.ZN(net9786)
);

AND3_X4 merge9138(
.A1(net5975),
.A2(net6115),
.A3(net7078),
.ZN(net9787)
);

DFFS_X2 merge9139(
.D(net5835),
.SN(net5854),
.CK(clk),
.Q(net9789),
.QN(net9788)
);

INV_X8 merge9140(
.A(net10185),
.ZN(net9790)
);

DFFR_X1 merge9141(
.D(net6053),
.RN(net6103),
.CK(clk),
.Q(net9792),
.QN(net9791)
);

SDFF_X2 merge9142(
.D(net5883),
.SE(net8832),
.SI(net8835),
.CK(clk),
.Q(net9794),
.QN(net9793)
);

DFFR_X2 merge9143(
.D(net6229),
.RN(net5364),
.CK(clk),
.Q(net9796),
.QN(net9795)
);

INV_X16 merge9144(
.A(net9927),
.ZN(net9797)
);

DFFS_X1 merge9145(
.D(net1023),
.SN(net1019),
.CK(clk),
.Q(net9799),
.QN(net9798)
);

INV_X32 merge9146(
.A(net11087),
.ZN(net9800)
);

SDFFR_X2 merge9147(
.D(net3810),
.RN(net3878),
.SE(net5820),
.SI(net5764),
.CK(clk),
.Q(net9802),
.QN(net9801)
);

INV_X4 merge9148(
.A(net10316),
.ZN(net9803)
);

SDFFS_X1 merge9149(
.D(net5332),
.SE(net4755),
.SI(net1635),
.SN(net3736),
.CK(clk),
.Q(net9805),
.QN(net9804)
);

INV_X1 merge9150(
.A(net10242),
.ZN(net9806)
);

SDFFS_X2 merge9151(
.D(net8522),
.SE(net8207),
.SI(net6645),
.SN(net4664),
.CK(clk),
.Q(net9808),
.QN(net9807)
);

INV_X2 merge9152(
.A(net10696),
.ZN(net9809)
);

NOR4_X4 merge9153(
.A1(net6608),
.A2(net6632),
.A3(net2849),
.A4(net5776),
.ZN(net9810)
);

DFFRS_X1 merge9154(
.D(net41),
.RN(net37),
.SN(net108),
.CK(clk),
.Q(net9812),
.QN(net9811)
);

DFFS_X2 merge9155(
.D(net235),
.SN(net1108),
.CK(clk),
.Q(net9814),
.QN(net9813)
);

INV_X8 merge9156(
.A(net10159),
.ZN(net9815)
);

INV_X16 merge9157(
.A(net10363),
.ZN(net9816)
);

DFFR_X1 merge9158(
.D(net5848),
.RN(net5854),
.CK(clk),
.Q(net9818),
.QN(net9817)
);

INV_X32 merge9159(
.A(net11460),
.ZN(net9819)
);

SDFFR_X1 merge9160(
.D(net4512),
.RN(net9077),
.SE(net9546),
.SI(net9537),
.CK(clk),
.Q(net9821),
.QN(net9820)
);

NOR4_X2 merge9161(
.A1(net8433),
.A2(net4588),
.A3(net7689),
.A4(net7674),
.ZN(net9822)
);

DFFR_X2 merge9162(
.D(net6850),
.RN(net6989),
.CK(clk),
.Q(net9824),
.QN(net9823)
);

DFFS_X1 merge9163(
.D(net4365),
.SN(net5329),
.CK(clk),
.Q(net9826),
.QN(net9825)
);

AND2_X1 merge9164(
.A1(net1190),
.A2(net342),
.ZN(net9827)
);

INV_X4 merge9165(
.A(net10029),
.ZN(net9828)
);

DFFS_X2 merge9166(
.D(net6821),
.SN(net6867),
.CK(clk),
.Q(net9830),
.QN(net9829)
);

INV_X1 merge9167(
.A(net10119),
.ZN(net9831)
);

INV_X2 merge9168(
.A(net10304),
.ZN(net9832)
);

SDFFR_X2 merge9169(
.D(net2772),
.RN(net5375),
.SE(net6625),
.SI(net6629),
.CK(clk),
.Q(net9834),
.QN(net9833)
);

SDFFS_X1 merge9170(
.D(net6657),
.SE(net7495),
.SI(net8595),
.SN(net8618),
.CK(clk),
.Q(net9836),
.QN(net9835)
);

DFFR_X1 merge9171(
.D(net7798),
.RN(net5086),
.CK(clk),
.Q(net9838),
.QN(net9837)
);

DFFR_X2 merge9172(
.D(net8748),
.RN(net5838),
.CK(clk),
.Q(net9840),
.QN(net9839)
);

DFFS_X1 merge9173(
.D(net4028),
.SN(net4163),
.CK(clk),
.Q(net9842),
.QN(net9841)
);

INV_X8 merge9174(
.A(net10147),
.ZN(net9843)
);

NAND2_X1 merge9175(
.A1(net192),
.A2(net284),
.ZN(net9844)
);

INV_X16 merge9176(
.A(net11473),
.ZN(net9845)
);

SDFFS_X2 merge9177(
.D(net8297),
.SE(net7312),
.SI(net9165),
.SN(net8953),
.CK(clk),
.Q(net9847),
.QN(net9846)
);

INV_X32 merge9178(
.A(net11465),
.ZN(net9848)
);

INV_X4 merge9179(
.A(net11441),
.ZN(net9849)
);

INV_X1 merge9180(
.A(net10414),
.ZN(net9850)
);

DFFS_X2 merge9181(
.D(net6833),
.SN(net6848),
.CK(clk),
.Q(net9852),
.QN(net9851)
);

INV_X2 merge9182(
.A(net10201),
.ZN(net9853)
);

DFFR_X1 merge9183(
.D(net527),
.RN(net640),
.CK(clk),
.Q(net9855),
.QN(net9854)
);

INV_X8 merge9184(
.A(net10249),
.ZN(net9856)
);

DFFR_X2 merge9185(
.D(net3445),
.RN(net4500),
.CK(clk),
.Q(net9858),
.QN(net9857)
);

INV_X16 merge9186(
.A(net10393),
.ZN(net9859)
);

DFFS_X1 merge9187(
.D(net1970),
.SN(net166),
.CK(clk),
.Q(net9861),
.QN(net9860)
);

DFFS_X2 merge9188(
.D(net5947),
.SN(net5882),
.CK(clk),
.Q(net9863),
.QN(net9862)
);

NAND2_X2 merge9189(
.A1(net259),
.A2(net218),
.ZN(net9864)
);

INV_X32 merge9190(
.A(net10044),
.ZN(net9865)
);

NAND2_X4 merge9191(
.A1(net5933),
.A2(net6942),
.ZN(net9866)
);

SDFFR_X1 merge9192(
.D(net7551),
.RN(net7359),
.SE(net5351),
.SI(net11429),
.CK(clk),
.Q(net9868),
.QN(net9867)
);

INV_X4 merge9193(
.A(net10349),
.ZN(net9869)
);

INV_X1 merge9194(
.A(net10695),
.ZN(net9870)
);

NAND3_X2 merge9195(
.A1(net4558),
.A2(net6478),
.A3(net5556),
.ZN(net9871)
);

DFFRS_X2 merge9196(
.D(net6308),
.RN(net7167),
.SN(net7255),
.CK(clk),
.Q(net9873),
.QN(net9872)
);

DFFR_X1 merge9197(
.D(net5042),
.RN(net5076),
.CK(clk),
.Q(net9875),
.QN(net9874)
);

SDFFR_X2 merge9198(
.D(net9300),
.RN(net7900),
.SE(net8343),
.SI(net8330),
.CK(clk),
.Q(net9877),
.QN(net9876)
);

DFFR_X2 merge9199(
.D(net1019),
.RN(net1029),
.CK(clk),
.Q(net9879),
.QN(net9878)
);

SDFFS_X1 merge9200(
.D(net6212),
.SE(net5595),
.SI(net4682),
.SN(net4588),
.CK(clk),
.Q(net9881),
.QN(net9880)
);

INV_X2 merge9201(
.A(net10432),
.ZN(net9882)
);

DFFS_X1 merge9202(
.D(net5886),
.SN(net5938),
.CK(clk),
.Q(net9884),
.QN(net9883)
);

INV_X8 merge9203(
.A(net11193),
.ZN(net9885)
);

SDFFS_X2 merge9204(
.D(net7634),
.SE(net8666),
.SI(net7519),
.SN(net9606),
.CK(clk),
.Q(net9887),
.QN(net9886)
);

INV_X16 merge9205(
.A(net10243),
.ZN(net9888)
);

INV_X32 merge9206(
.A(net10321),
.ZN(net9889)
);

INV_X4 merge9207(
.A(net10196),
.ZN(net9890)
);

INV_X1 merge9208(
.A(net10129),
.ZN(net9891)
);

OR3_X1 merge9209(
.A1(net6982),
.A2(net8942),
.A3(net7109),
.ZN(net9892)
);

AOI211_X4 merge9210(
.A(net3610),
.B(net1806),
.C1(net4684),
.C2(net3780),
.ZN(net9893)
);

SDFFR_X1 merge9211(
.D(net7186),
.RN(net5181),
.SE(net8186),
.SI(net8166),
.CK(clk),
.Q(net9895),
.QN(net9894)
);

INV_X2 merge9212(
.A(net11084),
.ZN(net9896)
);

DFFS_X2 merge9213(
.D(net2983),
.SN(net3899),
.CK(clk),
.Q(net9898),
.QN(net9897)
);

SDFFR_X2 merge9214(
.D(net8099),
.RN(net8089),
.SE(net8150),
.SI(net8214),
.CK(clk),
.Q(net9900),
.QN(net9899)
);

NOR4_X1 merge9215(
.A1(net5664),
.A2(net5684),
.A3(net5634),
.A4(net5669),
.ZN(net9901)
);

INV_X8 merge9216(
.A(net10109),
.ZN(net9902)
);

AOI211_X2 merge9217(
.A(net1382),
.B(net4028),
.C1(net4212),
.C2(net3129),
.ZN(net9903)
);

SDFFS_X1 merge9218(
.D(net4437),
.SE(net4431),
.SI(net3512),
.SN(net2629),
.CK(clk),
.Q(net9905),
.QN(net9904)
);

INV_X16 merge9219(
.A(net10213),
.ZN(net9906)
);

INV_X32 merge9220(
.A(net11252),
.ZN(net9907)
);

SDFFS_X2 merge9221(
.D(net8444),
.SE(net6541),
.SI(net4691),
.SN(net6462),
.CK(clk),
.Q(net9909),
.QN(net9908)
);

INV_X4 merge9222(
.A(net11223),
.ZN(net9910)
);

MUX2_X1 merge9223(
.A(net2600),
.B(net3690),
.S(net4588),
.Z(net9911)
);

INV_X1 merge9224(
.A(net10154),
.ZN(net9912)
);

INV_X2 merge9225(
.A(net10022),
.ZN(net9913)
);

DFFR_X1 merge9226(
.D(net410),
.RN(net640),
.CK(clk),
.Q(net9915),
.QN(net9914)
);

SDFFR_X1 merge9227(
.D(net5211),
.RN(net2294),
.SE(net5215),
.SI(net4321),
.CK(clk),
.Q(net9917),
.QN(net9916)
);

INV_X8 merge9228(
.A(net10146),
.ZN(net9918)
);

SDFFR_X2 merge9229(
.D(net4675),
.RN(net4726),
.SE(net2623),
.SI(net2863),
.CK(clk),
.Q(net9920),
.QN(net9919)
);

SDFF_X1 merge9230(
.D(net6052),
.SE(net5061),
.SI(net6028),
.CK(clk),
.Q(net9922),
.QN(net9921)
);

SDFFS_X1 merge9231(
.D(net8265),
.SE(net8228),
.SI(net7288),
.SN(net8215),
.CK(clk),
.Q(net9924),
.QN(net9923)
);

SDFFS_X2 merge9232(
.D(net7370),
.SE(net7356),
.SI(net6434),
.SN(net6437),
.CK(clk),
.Q(net9926),
.QN(net9925)
);

SDFFR_X1 merge9233(
.D(net3651),
.RN(net3529),
.SE(net1722),
.SI(net2501),
.CK(clk),
.Q(net9928),
.QN(net9927)
);

DFFR_X2 merge9234(
.D(net2986),
.RN(net1986),
.CK(clk),
.Q(net9930),
.QN(net9929)
);

SDFF_X2 merge9235(
.D(net8471),
.SE(net8235),
.SI(net8390),
.CK(clk),
.Q(net9932),
.QN(net9931)
);

DFFS_X1 merge9236(
.D(net1454),
.SN(net1484),
.CK(clk),
.Q(net9934),
.QN(net9933)
);

DFFS_X2 merge9237(
.D(net6822),
.SN(net5900),
.CK(clk),
.Q(net9936),
.QN(net9935)
);

AND2_X2 merge9238(
.A1(net457),
.A2(net1474),
.ZN(net9937)
);

SDFFR_X2 merge9239(
.D(net7459),
.RN(net5388),
.SE(net7295),
.SI(net6522),
.CK(clk),
.Q(net9939),
.QN(net9938)
);

DFFRS_X1 merge9240(
.D(net1436),
.RN(net2618),
.SN(net2617),
.CK(clk),
.Q(net9941),
.QN(net9940)
);

DFFR_X1 merge9241(
.D(net2967),
.RN(net3899),
.CK(clk),
.Q(net9943),
.QN(net9942)
);

SDFFS_X1 merge9242(
.D(net7970),
.SE(net6993),
.SI(net7227),
.SN(net7224),
.CK(clk),
.Q(net9945),
.QN(net9944)
);

DFFR_X2 merge9243(
.D(net7822),
.RN(net6822),
.CK(clk),
.Q(net9947),
.QN(net9946)
);

AOI22_X1 merge9244(
.A1(net2270),
.A2(net5134),
.B1(net4182),
.B2(net4130),
.ZN(net9948)
);

SDFFS_X2 merge9245(
.D(net7351),
.SE(net7348),
.SI(net9293),
.SN(net9047),
.CK(clk),
.Q(net9950),
.QN(net9949)
);

INV_X16 merge9246(
.A(net10133),
.ZN(net9951)
);

SDFFR_X1 merge9247(
.D(net6655),
.RN(net7642),
.SE(net5726),
.SI(net5662),
.CK(clk),
.Q(net9953),
.QN(net9952)
);

OAI21_X4 merge9248(
.A(net954),
.B1(net223),
.B2(net1292),
.ZN(net9954)
);

SDFFR_X2 merge9249(
.D(net8228),
.RN(net7287),
.SE(net6259),
.SI(net7292),
.CK(clk),
.Q(net9956),
.QN(net9955)
);

SDFFS_X1 merge9250(
.D(net1673),
.SE(net1680),
.SI(net3453),
.SN(net3528),
.CK(clk),
.Q(net9958),
.QN(net9957)
);

AND4_X4 merge9251(
.A1(net5599),
.A2(net6491),
.A3(net5629),
.A4(net5596),
.ZN(net9959)
);

XOR2_X1 merge9252(
.A(net6847),
.B(net5864),
.Z(net9960)
);

NAND4_X1 merge9253(
.A1(net2463),
.A2(net2358),
.A3(net2241),
.A4(net3173),
.ZN(net9961)
);

SDFFS_X2 merge9254(
.D(net7421),
.SE(net6616),
.SI(net9365),
.SN(net9253),
.CK(clk),
.Q(net9963),
.QN(net9962)
);

SDFFR_X1 merge9255(
.D(net5614),
.RN(net3497),
.SE(net6522),
.SI(net6472),
.CK(clk),
.Q(net9965),
.QN(net9964)
);

SDFFR_X2 merge9256(
.D(net1679),
.RN(net1692),
.SE(net744),
.SI(net86),
.CK(clk),
.Q(net9967),
.QN(net9966)
);

SDFFS_X1 merge9257(
.D(net8326),
.SE(net6238),
.SI(net8328),
.SN(net11560),
.CK(clk),
.Q(net9969),
.QN(net9968)
);

SDFFS_X2 merge9258(
.D(net2651),
.SE(net1690),
.SI(net1711),
.SN(net11149),
.CK(clk),
.Q(net9971),
.QN(net9970)
);

SDFFR_X1 merge9259(
.D(net5177),
.RN(net6132),
.SE(net3182),
.SI(net7037),
.CK(clk),
.Q(net9973),
.QN(net9972)
);

SDFFR_X2 merge9260(
.D(net7319),
.RN(net7903),
.SE(net6163),
.SI(net5413),
.CK(clk),
.Q(net9975),
.QN(net9974)
);

SDFFS_X1 merge9261(
.D(net8452),
.SE(net8469),
.SI(net4611),
.SN(net4620),
.CK(clk),
.Q(net9977),
.QN(net9976)
);

SDFFS_X2 merge9262(
.D(net7536),
.SE(net7627),
.SI(net7436),
.SN(net6418),
.CK(clk),
.Q(net9979),
.QN(net9978)
);

SDFFR_X1 merge9263(
.D(net8213),
.RN(net1288),
.SE(net4173),
.SI(net11478),
.CK(clk),
.Q(net9981),
.QN(net9980)
);

SDFFR_X2 merge9264(
.D(net6870),
.RN(net7376),
.SE(net7277),
.SI(net8382),
.CK(clk),
.Q(net9983),
.QN(net9982)
);

DFFS_X1 merge9265(
.D(net5843),
.SN(net2986),
.CK(clk),
.Q(net9985),
.QN(net9984)
);

OR4_X1 merge9266(
.A1(net3634),
.A2(net3612),
.A3(net3663),
.A4(net3354),
.ZN(net9986)
);

OAI22_X1 merge9267(
.A1(net6506),
.A2(net4534),
.B1(net8320),
.B2(net8002),
.ZN(net9987)
);

AND4_X2 merge9268(
.A1(net6172),
.A2(net6363),
.A3(net6292),
.A4(net6364),
.ZN(net9988)
);

SDFFS_X1 merge9269(
.D(net2537),
.SE(net2552),
.SI(net677),
.SN(net1624),
.CK(clk),
.Q(net9990),
.QN(net9989)
);

DFFRS_X2 merge9270(
.D(net2049),
.RN(net1130),
.SN(net3172),
.CK(clk),
.Q(net9992),
.QN(net9991)
);

DFFS_X2 merge9271(
.D(net1916),
.SN(net1947),
.CK(clk),
.Q(net9994),
.QN(net9993)
);

AND4_X1 merge9272(
.A1(net6573),
.A2(net6571),
.A3(net8108),
.A4(net8290),
.ZN(net9995)
);

AOI22_X4 merge9273(
.A1(net4349),
.A2(net2589),
.B1(net3393),
.B2(net4620),
.ZN(net9996)
);

OAI22_X4 merge9274(
.A1(net1723),
.A2(net1749),
.B1(net2662),
.B2(net1791),
.ZN(net9997)
);

SDFFS_X2 merge9275(
.D(net6509),
.SE(net6538),
.SI(net3622),
.SN(net3615),
.CK(clk),
.Q(net9999),
.QN(net9998)
);

AOI22_X2 merge9276(
.A1(net3676),
.A2(net3611),
.B1(net3677),
.B2(net4595),
.ZN(net10000)
);

SDFFR_X1 merge9277(
.D(net4136),
.RN(net4124),
.SE(net5120),
.SI(net10558),
.CK(clk),
.Q(net10002),
.QN(net10001)
);

NAND4_X4 merge9278(
.A1(net8501),
.A2(net4712),
.A3(net5652),
.A4(net11111),
.ZN(net10003)
);

OAI211_X2 merge9279(
.A(net316),
.B(net315),
.C1(net3096),
.C2(net3084),
.ZN(net10004)
);

SDFF_X1 merge9280(
.D(net7848),
.SE(net7987),
.SI(net5953),
.CK(clk),
.Q(net10006),
.QN(net10005)
);

OR4_X2 merge9281(
.A1(net560),
.A2(net523),
.A3(net463),
.A4(net11044),
.ZN(net10007)
);

AOI211_X1 merge9282(
.A(net63),
.B(net153),
.C1(net3099),
.C2(net1035),
.ZN(net10008)
);

SDFFR_X2 merge9283(
.D(net2679),
.RN(net3660),
.SE(net4613),
.SI(net4495),
.CK(clk),
.Q(net10010),
.QN(net10009)
);

NAND4_X2 merge9284(
.A1(net4065),
.A2(net4052),
.A3(net4212),
.A4(net10898),
.ZN(net10011)
);

OR4_X4 merge9285(
.A1(net760),
.A2(net1741),
.A3(net4627),
.A4(net3688),
.ZN(net10012)
);

SDFFS_X1 merge9286(
.D(net3368),
.SE(net2446),
.SI(net3416),
.SN(net2314),
.CK(clk),
.Q(net10014),
.QN(net10013)
);

OAI22_X2 merge9287(
.A1(net2127),
.A2(net1453),
.B1(net415),
.B2(net350),
.ZN(net10015)
);

SDFFS_X2 merge9288(
.D(net3149),
.SE(net4431),
.SI(net1427),
.SN(net1401),
.CK(clk),
.Q(net10017),
.QN(net10016)
);

OAI211_X4 merge9289(
.A(net132),
.B(net233),
.C1(net3985),
.C2(net4038),
.ZN(net10018)
);

SDFFR_X1 merge9290(
.D(net7183),
.RN(net6808),
.SE(net7098),
.SI(net4239),
.CK(clk),
.Q(net10020),
.QN(net10019)
);

SDFFR_X2 merge9291(
.D(net1777),
.RN(net744),
.SE(net828),
.SI(net833),
.CK(clk),
.Q(net10022),
.QN(net10021)
);

OAI211_X1 merge9292(
.A(net1210),
.B(net2220),
.C1(net1252),
.C2(net1036),
.ZN(net10023)
);

SDFFS_X1 merge9293(
.D(net3308),
.SE(net2585),
.SI(net523),
.SN(net520),
.CK(clk),
.Q(net10025),
.QN(net10024)
);

SDFFS_X2 merge9294(
.D(net5649),
.SE(net3810),
.SI(net7493),
.SN(net5551),
.CK(clk),
.Q(net10027),
.QN(net10026)
);

SDFFR_X1 merge9295(
.D(net3391),
.RN(net2318),
.SE(net4394),
.SI(net4028),
.CK(clk),
.Q(net10029),
.QN(net10028)
);

SDFFR_X2 merge9296(
.D(net6525),
.RN(net6333),
.SE(net8477),
.SI(net6472),
.CK(clk),
.Q(net10031),
.QN(net10030)
);

SDFFS_X1 merge9297(
.D(net6638),
.SE(net5646),
.SI(net6333),
.SN(net11342),
.CK(clk),
.Q(net10033),
.QN(net10032)
);

NOR4_X4 merge9298(
.A1(net8934),
.A2(net8922),
.A3(net8924),
.A4(net10967),
.ZN(net10034)
);

NOR4_X2 merge9299(
.A1(net7016),
.A2(net6989),
.A3(net6994),
.A4(net6996),
.ZN(net10035)
);

SDFFS_X2 merge9300(
.D(net7487),
.SE(net7376),
.SI(net7324),
.SN(net4205),
.CK(clk),
.Q(net10037),
.QN(net10036)
);

SDFFR_X1 merge9301(
.D(net4214),
.RN(net5137),
.SE(net5162),
.SI(net11040),
.CK(clk),
.Q(net10039),
.QN(net10038)
);

SDFFR_X2 merge9302(
.D(net5057),
.RN(net5120),
.SE(net6934),
.SI(net6982),
.CK(clk),
.Q(net10041),
.QN(net10040)
);

SDFFS_X1 merge9303(
.D(net7226),
.SE(net7215),
.SI(net6993),
.SN(net8197),
.CK(clk),
.Q(net10043),
.QN(net10042)
);

SDFFS_X2 merge9304(
.D(net6026),
.SE(net6028),
.SI(net3904),
.SN(net7075),
.CK(clk),
.Q(net10045),
.QN(net10044)
);

SDFFR_X1 merge9305(
.D(net5604),
.RN(net5652),
.SE(net8460),
.SI(net6616),
.CK(clk),
.Q(net10047),
.QN(net10046)
);

AOI211_X4 merge9306(
.A(net3646),
.B(net4620),
.C1(net1571),
.C2(net483),
.ZN(net10048)
);

SDFFR_X2 merge9307(
.D(net6076),
.RN(net6082),
.SE(net7028),
.SI(net6989),
.CK(clk),
.Q(net10050),
.QN(net10049)
);

NOR4_X1 merge9308(
.A1(net1526),
.A2(net1418),
.A3(net2536),
.A4(net2531),
.ZN(net10051)
);

AOI211_X2 merge9309(
.A(net5951),
.B(net5975),
.C1(net5856),
.C2(net3038),
.ZN(net10052)
);

SDFFS_X1 merge9310(
.D(net8849),
.SE(net8859),
.SI(net6939),
.SN(net6968),
.CK(clk),
.Q(net10054),
.QN(net10053)
);

SDFFS_X2 merge9311(
.D(net5928),
.SE(net3991),
.SI(net5017),
.SN(net4932),
.CK(clk),
.Q(net10056),
.QN(net10055)
);

SDFFR_X1 merge9312(
.D(net108),
.RN(net973),
.SE(net1056),
.SI(net1091),
.CK(clk),
.Q(net10058),
.QN(net10057)
);

SDFFR_X2 merge9313(
.D(net1864),
.RN(net1880),
.SE(net772),
.SI(net777),
.CK(clk),
.Q(net10060),
.QN(net10059)
);

SDFFS_X1 merge9314(
.D(net5245),
.SE(net3981),
.SI(net1402),
.SN(net1436),
.CK(clk),
.Q(net10062),
.QN(net10061)
);

AOI22_X1 merge9315(
.A1(net6302),
.A2(net7273),
.B1(net8117),
.B2(net11413),
.ZN(net10063)
);

AND4_X4 merge9316(
.A1(net2672),
.A2(net2685),
.A3(net3620),
.A4(net3496),
.ZN(net10064)
);

NAND4_X1 merge9317(
.A1(net6491),
.A2(net6195),
.A3(net5589),
.A4(net4495),
.ZN(net10065)
);

SDFFS_X2 merge9318(
.D(net4201),
.SE(net7056),
.SI(net8095),
.SN(net7796),
.CK(clk),
.Q(net10067),
.QN(net10066)
);

SDFFR_X1 merge9319(
.D(net461),
.RN(net465),
.SE(net2299),
.SI(net2241),
.CK(clk),
.Q(net10069),
.QN(net10068)
);

OR4_X1 merge9320(
.A1(net5328),
.A2(net5360),
.A3(net5357),
.A4(net6172),
.ZN(net10070)
);

OAI22_X1 merge9321(
.A1(net5258),
.A2(net6387),
.B1(net7083),
.B2(net6212),
.ZN(net10071)
);

AND4_X2 merge9322(
.A1(net8467),
.A2(net8336),
.A3(net7505),
.A4(net7508),
.ZN(net10072)
);

SDFFR_X2 merge9323(
.D(net6972),
.RN(net5028),
.SE(net5950),
.SI(net5880),
.CK(clk),
.Q(net10074),
.QN(net10073)
);

SDFFS_X1 merge9324(
.D(net6365),
.SE(net1546),
.SI(net559),
.SN(net10843),
.CK(clk),
.Q(net10076),
.QN(net10075)
);

AND4_X1 merge9325(
.A1(net6528),
.A2(net8366),
.A3(net9341),
.A4(net9397),
.ZN(net10077)
);

SDFFS_X2 merge9326(
.D(net2585),
.SE(net3446),
.SI(net1453),
.SN(net3593),
.CK(clk),
.Q(net10079),
.QN(net10078)
);

AOI22_X4 merge9327(
.A1(net3740),
.A2(net3704),
.B1(net2760),
.B2(net2773),
.ZN(net10080)
);

OAI22_X4 merge9328(
.A1(net7338),
.A2(net6555),
.B1(net6533),
.B2(net11013),
.ZN(net10081)
);

AOI22_X2 merge9329(
.A1(net4069),
.A2(net2135),
.B1(net5062),
.B2(net5094),
.ZN(net10082)
);

SDFFR_X1 merge9330(
.D(net275),
.RN(net25),
.SE(net1993),
.SI(net2135),
.CK(clk),
.Q(net10084),
.QN(net10083)
);

NAND4_X4 merge9331(
.A1(net6239),
.A2(net6238),
.A3(net1391),
.A4(net3257),
.ZN(net10085)
);

SDFFR_X2 merge9332(
.D(net7350),
.RN(net5458),
.SE(net2388),
.SI(net3226),
.CK(clk),
.Q(net10087),
.QN(net10086)
);

SDFFS_X1 merge9333(
.D(net6476),
.SE(net8418),
.SI(net7249),
.SN(net8131),
.CK(clk),
.Q(net10089),
.QN(net10088)
);

SDFFS_X2 merge9334(
.D(net5073),
.SE(net5089),
.SI(net5876),
.SN(net5117),
.CK(clk),
.Q(net10091),
.QN(net10090)
);

OAI211_X2 merge9335(
.A(net4714),
.B(net4595),
.C1(net5473),
.C2(net5474),
.ZN(net10092)
);

SDFFR_X1 merge9336(
.D(net5587),
.RN(net5602),
.SE(net3841),
.SI(net5763),
.CK(clk),
.Q(net10094),
.QN(net10093)
);

SDFFR_X2 merge9337(
.D(net6466),
.RN(net6678),
.SE(net5556),
.SI(net5553),
.CK(clk),
.Q(net10096),
.QN(net10095)
);

SDFFS_X1 merge9338(
.D(net3507),
.SE(net3463),
.SI(net592),
.SN(net554),
.CK(clk),
.Q(net10098),
.QN(net10097)
);

SDFFS_X2 merge9339(
.D(net3062),
.SE(net3060),
.SI(net3139),
.SN(net3133),
.CK(clk),
.Q(net10100),
.QN(net10099)
);

OR4_X2 merge9340(
.A1(net962),
.A2(net2077),
.A3(net153),
.A4(net2987),
.ZN(net10101)
);

SDFFR_X1 merge9341(
.D(net7366),
.RN(net7189),
.SE(net6532),
.SI(net6533),
.CK(clk),
.Q(net10103),
.QN(net10102)
);

SDFFR_X2 merge9342(
.D(net9224),
.RN(net8235),
.SE(net9283),
.SI(net9399),
.CK(clk),
.Q(net10105),
.QN(net10104)
);

AOI211_X1 merge9343(
.A(net1070),
.B(net1108),
.C1(net2022),
.C2(net2077),
.ZN(net10106)
);

SDFFS_X1 merge9344(
.D(net1193),
.SE(net4234),
.SI(net4273),
.SN(net4168),
.CK(clk),
.Q(net10108),
.QN(net10107)
);

SDFFS_X2 merge9345(
.D(net999),
.SE(net1310),
.SI(net1110),
.SN(net1298),
.CK(clk),
.Q(net10110),
.QN(net10109)
);

SDFFR_X1 merge9346(
.D(net1035),
.RN(net325),
.SE(net276),
.SI(net1132),
.CK(clk),
.Q(net10112),
.QN(net10111)
);

NAND4_X2 merge9347(
.A1(net5925),
.A2(net6262),
.A3(net8187),
.A4(net7093),
.ZN(net10113)
);

SDFFR_X2 merge9348(
.D(net4665),
.RN(net5545),
.SE(net4520),
.SI(net4702),
.CK(clk),
.Q(net10115),
.QN(net10114)
);

OR4_X4 merge9349(
.A1(net410),
.A2(net1418),
.A3(net6196),
.A4(net6198),
.ZN(net10116)
);

SDFFS_X1 merge9350(
.D(net4336),
.SE(net4595),
.SI(net2730),
.SN(net2695),
.CK(clk),
.Q(net10118),
.QN(net10117)
);

SDFFS_X2 merge9351(
.D(net1257),
.SE(net1250),
.SI(net1080),
.SN(net2180),
.CK(clk),
.Q(net10120),
.QN(net10119)
);

OAI22_X2 merge9352(
.A1(net3238),
.A2(net3246),
.B1(net1269),
.B2(net4160),
.ZN(net10121)
);

SDFFR_X1 merge9353(
.D(net6867),
.RN(net5092),
.SE(net6993),
.SI(net11185),
.CK(clk),
.Q(net10123),
.QN(net10122)
);

SDFFR_X2 merge9354(
.D(net6544),
.RN(net6384),
.SE(net2626),
.SI(net3508),
.CK(clk),
.Q(net10125),
.QN(net10124)
);

SDFFS_X1 merge9355(
.D(net8004),
.SE(net8860),
.SI(net8955),
.SN(net8924),
.CK(clk),
.Q(net10127),
.QN(net10126)
);

SDFFS_X2 merge9356(
.D(net7814),
.SE(net4038),
.SI(net7068),
.SN(net7066),
.CK(clk),
.Q(net10129),
.QN(net10128)
);

SDFFR_X1 merge9357(
.D(net2511),
.RN(net2491),
.SE(net3466),
.SI(net3308),
.CK(clk),
.Q(net10131),
.QN(net10130)
);

OAI211_X4 merge9358(
.A(net3635),
.B(net2726),
.C1(net2746),
.C2(net11268),
.ZN(net10132)
);

SDFFR_X2 merge9359(
.D(net2042),
.RN(net1944),
.SE(net2100),
.SI(net1140),
.CK(clk),
.Q(net10134),
.QN(net10133)
);

OAI211_X1 merge9360(
.A(net3577),
.B(net3565),
.C1(net4435),
.C2(net4557),
.ZN(net10135)
);

SDFFS_X1 merge9361(
.D(net6952),
.SE(net6980),
.SI(net5932),
.SN(net5947),
.CK(clk),
.Q(net10137),
.QN(net10136)
);

NOR4_X4 merge9362(
.A1(net5295),
.A2(net6199),
.A3(net2417),
.A4(net2416),
.ZN(net10138)
);

NOR4_X2 merge9363(
.A1(net1741),
.A2(net1737),
.A3(net3649),
.A4(net3633),
.ZN(net10139)
);

SDFFS_X2 merge9364(
.D(net5033),
.SE(net4117),
.SI(net6032),
.SN(net6028),
.CK(clk),
.Q(net10141),
.QN(net10140)
);

AOI211_X4 merge9365(
.A(net1812),
.B(net2735),
.C1(net903),
.C2(net925),
.ZN(net10142)
);

SDFFR_X1 merge9366(
.D(net5224),
.RN(net8185),
.SE(net9130),
.SI(net11124),
.CK(clk),
.Q(net10144),
.QN(net10143)
);

SDFFR_X2 merge9367(
.D(net483),
.RN(net675),
.SE(net3545),
.SI(net2459),
.CK(clk),
.Q(net10146),
.QN(net10145)
);

SDFFS_X1 merge9368(
.D(net6217),
.SE(net6259),
.SI(net5299),
.SN(net5170),
.CK(clk),
.Q(net10148),
.QN(net10147)
);

SDFFS_X2 merge9369(
.D(net6498),
.SE(net6493),
.SI(net7505),
.SN(net11373),
.CK(clk),
.Q(net10150),
.QN(net10149)
);

NOR4_X1 merge9370(
.A1(net421),
.A2(net875),
.A3(net3572),
.A4(net3445),
.ZN(net10151)
);

SDFFR_X1 merge9371(
.D(net4493),
.RN(net5500),
.SE(net5530),
.SI(net6418),
.CK(clk),
.Q(net10153),
.QN(net10152)
);

SDFFR_X2 merge9372(
.D(net3256),
.RN(net1341),
.SE(net417),
.SI(net461),
.CK(clk),
.Q(net10155),
.QN(net10154)
);

SDFFS_X1 merge9373(
.D(net5434),
.SE(net4445),
.SI(net2491),
.SN(net2351),
.CK(clk),
.Q(net10157),
.QN(net10156)
);

SDFFS_X2 merge9374(
.D(net4950),
.SE(net5098),
.SI(net5932),
.SN(net11548),
.CK(clk),
.Q(net10159),
.QN(net10158)
);

SDFFR_X1 merge9375(
.D(net7549),
.RN(net7536),
.SE(net7467),
.SI(net7518),
.CK(clk),
.Q(net10161),
.QN(net10160)
);

AOI211_X2 merge9376(
.A(net2403),
.B(net2417),
.C1(net4544),
.C2(net4488),
.ZN(net10162)
);

SDFFR_X2 merge9377(
.D(net4431),
.RN(net6418),
.SE(net8360),
.SI(net8345),
.CK(clk),
.Q(net10164),
.QN(net10163)
);

AOI22_X1 merge9378(
.A1(net5540),
.A2(net6515),
.B1(net7123),
.B2(net6238),
.ZN(net10165)
);

SDFFS_X1 merge9379(
.D(net7017),
.SE(net7059),
.SI(net6832),
.SN(net6956),
.CK(clk),
.Q(net10167),
.QN(net10166)
);

SDFFS_X2 merge9380(
.D(net6252),
.SE(net6367),
.SI(net8267),
.SN(net6165),
.CK(clk),
.Q(net10169),
.QN(net10168)
);

AND4_X4 merge9381(
.A1(net1456),
.A2(net1416),
.A3(net1604),
.A4(net2650),
.ZN(net10170)
);

SDFFR_X1 merge9382(
.D(net9399),
.RN(net5547),
.SE(net5627),
.SI(net10515),
.CK(clk),
.Q(net10172),
.QN(net10171)
);

SDFFR_X2 merge9383(
.D(net6227),
.RN(net6195),
.SE(net7499),
.SI(net7487),
.CK(clk),
.Q(net10174),
.QN(net10173)
);

SDFFS_X1 merge9384(
.D(net2185),
.SE(net1190),
.SI(net1036),
.SN(net10865),
.CK(clk),
.Q(net10176),
.QN(net10175)
);

SDFFS_X2 merge9385(
.D(net2643),
.SE(net2650),
.SI(net2367),
.SN(net2366),
.CK(clk),
.Q(net10178),
.QN(net10177)
);

SDFFR_X1 merge9386(
.D(net8261),
.RN(net8294),
.SE(net6482),
.SI(net6195),
.CK(clk),
.Q(net10180),
.QN(net10179)
);

NAND4_X1 merge9387(
.A1(net274),
.A2(net294),
.A3(net3092),
.A4(net3071),
.ZN(net10181)
);

OR4_X1 merge9388(
.A1(net5535),
.A2(net5551),
.A3(net4488),
.A4(net5383),
.ZN(net10182)
);

SDFFR_X2 merge9389(
.D(net3518),
.RN(net5394),
.SE(net5677),
.SI(net2772),
.CK(clk),
.Q(net10184),
.QN(net10183)
);

SDFFS_X1 merge9390(
.D(net2311),
.SE(net2321),
.SI(net218),
.SN(net1108),
.CK(clk),
.Q(net10186),
.QN(net10185)
);

SDFFS_X2 merge9391(
.D(net7999),
.SE(net7792),
.SI(net6060),
.SN(net7045),
.CK(clk),
.Q(net10188),
.QN(net10187)
);

OAI22_X1 merge9392(
.A1(net3023),
.A2(net3140),
.B1(net3164),
.B2(net3080),
.ZN(net10189)
);

AND4_X2 merge9393(
.A1(net2420),
.A2(net3340),
.A3(net3423),
.A4(net3429),
.ZN(net10190)
);

SDFFR_X1 merge9394(
.D(net8018),
.RN(net7958),
.SE(net8972),
.SI(net8808),
.CK(clk),
.Q(net10192),
.QN(net10191)
);

SDFFR_X2 merge9395(
.D(net6126),
.RN(net6115),
.SE(net4207),
.SI(net5206),
.CK(clk),
.Q(net10194),
.QN(net10193)
);

SDFFS_X1 merge9396(
.D(net3340),
.SE(net3362),
.SI(net3563),
.SN(net4558),
.CK(clk),
.Q(net10196),
.QN(net10195)
);

AND4_X1 merge9397(
.A1(net3644),
.A2(net2511),
.A3(net3654),
.A4(net2717),
.ZN(net10197)
);

AOI22_X4 merge9398(
.A1(net2634),
.A2(net3622),
.B1(net4688),
.B2(net1599),
.ZN(net10198)
);

OAI22_X4 merge9399(
.A1(net5056),
.A2(net5120),
.B1(net1469),
.B2(net3424),
.ZN(net10199)
);

SDFFS_X2 merge9400(
.D(net6269),
.SE(net5253),
.SI(net5306),
.SN(net5274),
.CK(clk),
.Q(net10201),
.QN(net10200)
);

AOI22_X2 merge9401(
.A1(net4099),
.A2(net4069),
.B1(net4068),
.B2(net3940),
.ZN(net10202)
);

SDFFR_X1 merge9402(
.D(net4124),
.RN(net5974),
.SE(net8009),
.SI(net8016),
.CK(clk),
.Q(net10204),
.QN(net10203)
);

NAND4_X4 merge9403(
.A1(net454),
.A2(net449),
.A3(net5276),
.A4(net6199),
.ZN(net10205)
);

SDFFR_X2 merge9404(
.D(net7117),
.RN(net7249),
.SE(net7051),
.SI(net7050),
.CK(clk),
.Q(net10207),
.QN(net10206)
);

SDFFS_X1 merge9405(
.D(net5285),
.SE(net6209),
.SI(net5297),
.SN(net5330),
.CK(clk),
.Q(net10209),
.QN(net10208)
);

OAI211_X2 merge9406(
.A(net7439),
.B(net6541),
.C1(net8996),
.C2(net9012),
.ZN(net10210)
);

OR4_X2 merge9407(
.A1(net554),
.A2(net559),
.A3(net561),
.A4(net1428),
.ZN(net10211)
);

SDFFS_X2 merge9408(
.D(net1502),
.SE(net634),
.SI(net1605),
.SN(net1576),
.CK(clk),
.Q(net10213),
.QN(net10212)
);

SDFFR_X1 merge9409(
.D(net4555),
.RN(net6506),
.SE(net6566),
.SI(net5545),
.CK(clk),
.Q(net10215),
.QN(net10214)
);

SDFFR_X2 merge9410(
.D(net4830),
.RN(net5483),
.SE(net3516),
.SI(net3582),
.CK(clk),
.Q(net10217),
.QN(net10216)
);

AOI211_X1 merge9411(
.A(net4075),
.B(net4069),
.C1(net4112),
.C2(net4094),
.ZN(net10218)
);

NAND4_X2 merge9412(
.A1(net764),
.A2(net766),
.A3(net1734),
.A4(net1635),
.ZN(net10219)
);

OR4_X4 merge9413(
.A1(net3237),
.A2(net4548),
.A3(net4557),
.A4(net11512),
.ZN(net10220)
);

OAI22_X2 merge9414(
.A1(net3132),
.A2(net4146),
.B1(net5151),
.B2(net5125),
.ZN(net10221)
);

OAI211_X4 merge9415(
.A(net4166),
.B(net3199),
.C1(net4219),
.C2(net5162),
.ZN(net10222)
);

MUX2_X2 merge9416(
.A(net1229),
.B(net3181),
.S(net4159),
.Z(net10223)
);

OAI211_X1 merge9417(
.A(net5848),
.B(net5853),
.C1(net6001),
.C2(net5999),
.ZN(net10224)
);

SDFFS_X1 merge9418(
.D(net1733),
.SE(net2661),
.SI(net2513),
.SN(net2650),
.CK(clk),
.Q(net10226),
.QN(net10225)
);

SDFFS_X2 merge9419(
.D(net1563),
.SE(net4514),
.SI(net3445),
.SN(net11516),
.CK(clk),
.Q(net10228),
.QN(net10227)
);

SDFFR_X1 merge9420(
.D(net6197),
.RN(net3295),
.SE(net7956),
.SI(net8117),
.CK(clk),
.Q(net10230),
.QN(net10229)
);

NOR4_X4 merge9421(
.A1(net1119),
.A2(net3085),
.A3(net3168),
.A4(net4167),
.ZN(net10231)
);

SDFF_X2 merge9422(
.D(net4644),
.SE(net1703),
.SI(net3622),
.CK(clk),
.Q(net10233),
.QN(net10232)
);

NOR4_X2 merge9423(
.A1(net2395),
.A2(net2487),
.A3(net511),
.A4(net1286),
.ZN(net10234)
);

DFFRS_X1 merge9424(
.D(net3226),
.RN(net428),
.SN(net3359),
.CK(clk),
.Q(net10236),
.QN(net10235)
);

AOI211_X4 merge9425(
.A(net4101),
.B(net3104),
.C1(net4160),
.C2(net4273),
.ZN(net10237)
);

NOR4_X1 merge9426(
.A1(net1961),
.A2(net3117),
.A3(net4049),
.A4(net3035),
.ZN(net10238)
);

SDFFR_X2 merge9427(
.D(net3948),
.RN(net4948),
.SE(net4048),
.SI(net4957),
.CK(clk),
.Q(net10240),
.QN(net10239)
);

AOI211_X2 merge9428(
.A(net7050),
.B(net7074),
.C1(net6331),
.C2(net6376),
.ZN(net10241)
);

SDFFS_X1 merge9429(
.D(net1781),
.SE(net1775),
.SI(net3674),
.SN(net4610),
.CK(clk),
.Q(net10243),
.QN(net10242)
);

SDFFS_X2 merge9430(
.D(net6164),
.SE(net6182),
.SI(net7118),
.Q(net7076),
.CK(clk),
.QN(net10244)
);

SDFFR_X1 merge9431(
.D(net7149),
.RN(net7169),
.SE(net5210),
.SI(net5258),
.CK(clk),
.Q(net10247),
.QN(net10246)
);

SDFFR_X2 merge9432(
.D(net5377),
.RN(net2520),
.SE(net682),
.SI(net723),
.CK(clk),
.Q(net10249),
.QN(net10248)
);

SDFFS_X1 merge9433(
.D(net5351),
.SE(net8252),
.SI(net8339),
.SN(net11439),
.CK(clk),
.Q(net10251),
.QN(net10250)
);

AOI22_X1 merge9434(
.A1(net367),
.A2(net403),
.B1(net1310),
.B2(net1362),
.ZN(net10252)
);

SDFFS_X2 merge9435(
.D(net4347),
.SE(net4525),
.SI(net4565),
.SN(net4558),
.CK(clk),
.Q(net10254),
.QN(net10253)
);

AND4_X4 merge9436(
.A1(net3435),
.A2(net559),
.A3(net1680),
.A4(net1672),
.ZN(net10255)
);

SDFFR_X1 merge9437(
.D(net2180),
.RN(net2050),
.SE(net2178),
.SI(net2077),
.CK(clk),
.Q(net10257),
.QN(net10256)
);

SDFFR_X2 merge9438(
.D(net592),
.RN(net495),
.SE(net920),
.SI(net890),
.CK(clk),
.Q(net10259),
.QN(net10258)
);

SDFFS_X1 merge9439(
.D(net4264),
.SE(net4281),
.SI(net488),
.SN(net465),
.CK(clk),
.Q(net10261),
.QN(net10260)
);

NAND4_X1 merge9440(
.A1(net3310),
.A2(net3308),
.A3(net4261),
.A4(net4160),
.ZN(net10262)
);

OR4_X1 merge9441(
.A1(net3117),
.A2(net2907),
.A3(net4105),
.A4(net2122),
.ZN(net10263)
);

SDFFS_X2 merge9442(
.D(net3158),
.SE(net3108),
.SI(net4980),
.SN(net4949),
.CK(clk),
.Q(net10265),
.QN(net10264)
);

SDFFR_X1 merge9443(
.D(net2846),
.RN(net2870),
.SE(net3736),
.SI(net10673),
.CK(clk),
.Q(net10267),
.QN(net10266)
);

OAI22_X1 merge9444(
.A1(net2561),
.A2(net1647),
.B1(net4547),
.B2(net4563),
.ZN(net10268)
);

SDFFR_X2 merge9445(
.D(net4755),
.RN(net5711),
.SE(net5403),
.SI(net5267),
.CK(clk),
.Q(net10270),
.QN(net10269)
);

SDFFS_X1 merge9446(
.D(net2445),
.SE(net1613),
.SI(net6705),
.SN(net10634),
.CK(clk),
.Q(net10272),
.QN(net10271)
);

AND4_X2 merge9447(
.A1(net4460),
.A2(net4525),
.A3(net3602),
.A4(net5525),
.ZN(net10273)
);

SDFFS_X2 merge9448(
.D(net7963),
.SE(net8938),
.SI(net5953),
.SN(net7860),
.CK(clk),
.Q(net10275),
.QN(net10274)
);

SDFFR_X1 merge9449(
.D(net6176),
.RN(net6156),
.SE(net7953),
.SI(net7918),
.CK(clk),
.Q(net10277),
.QN(net10276)
);

SDFFR_X2 merge9450(
.D(net7354),
.RN(net7371),
.SE(net2566),
.SI(net652),
.CK(clk),
.Q(net10279),
.QN(net10278)
);

SDFFS_X1 merge9451(
.D(net4249),
.SE(net5301),
.SI(net5358),
.SN(net5253),
.CK(clk),
.Q(net10281),
.QN(net10280)
);

SDFFS_X2 merge9452(
.D(net483),
.SE(net1646),
.SI(net1610),
.SN(net677),
.CK(clk),
.Q(net10283),
.QN(net10282)
);

AND4_X1 merge9453(
.A1(net276),
.A2(net274),
.A3(net2399),
.A4(net3192),
.ZN(net10284)
);

SDFFR_X1 merge9454(
.D(net8196),
.RN(net5235),
.SE(net3474),
.SI(net1399),
.CK(clk),
.Q(net10286),
.QN(net10285)
);

SDFFR_X2 merge9455(
.D(net8301),
.RN(net8338),
.SE(net8023),
.SI(net8933),
.CK(clk),
.Q(net10288),
.QN(net10287)
);

SDFFS_X1 merge9456(
.D(net7434),
.SE(net6365),
.SI(net6276),
.SN(net6391),
.CK(clk),
.Q(net10290),
.QN(net10289)
);

AOI22_X4 merge9457(
.A1(net1282),
.A2(net1306),
.B1(net3470),
.B2(net3497),
.ZN(net10291)
);

OAI22_X4 merge9458(
.A1(net7107),
.A2(net7022),
.B1(net6152),
.B2(net6134),
.ZN(net10292)
);

SDFFS_X2 merge9459(
.D(net5100),
.SE(net4780),
.SI(net8379),
.SN(net5482),
.CK(clk),
.Q(net10294),
.QN(net10293)
);

AOI22_X2 merge9460(
.A1(net7857),
.A2(net7958),
.B1(net8043),
.B2(net5120),
.ZN(net10295)
);

NAND4_X4 merge9461(
.A1(net1677),
.A2(net1680),
.A3(net3528),
.A4(net3632),
.ZN(net10296)
);

SDFFR_X1 merge9462(
.D(net3794),
.RN(net3621),
.SE(net3441),
.SI(net11118),
.CK(clk),
.Q(net10298),
.QN(net10297)
);

SDFFR_X2 merge9463(
.D(net166),
.RN(net1133),
.SE(net3999),
.SI(net3952),
.CK(clk),
.Q(net10300),
.QN(net10299)
);

SDFFS_X1 merge9464(
.D(net2145),
.SE(net2158),
.SI(net3921),
.SN(net3940),
.CK(clk),
.Q(net10302),
.QN(net10301)
);

SDFFS_X2 merge9465(
.D(net1080),
.SE(net1024),
.SI(net1008),
.SN(net1029),
.CK(clk),
.Q(net10304),
.QN(net10303)
);

OAI211_X2 merge9466(
.A(net1324),
.B(net1330),
.C1(net4416),
.C2(net4423),
.ZN(net10305)
);

SDFFR_X1 merge9467(
.D(net6216),
.RN(net4071),
.SE(net1421),
.SI(net1430),
.CK(clk),
.Q(net10307),
.QN(net10306)
);

SDFFR_X2 merge9468(
.D(net7646),
.RN(net6675),
.SE(net5240),
.SI(net5717),
.CK(clk),
.Q(net10309),
.QN(net10308)
);

SDFFS_X1 merge9469(
.D(net6848),
.SE(net6945),
.SI(net8097),
.SN(net8064),
.CK(clk),
.Q(net10311),
.QN(net10310)
);

OR4_X2 merge9470(
.A1(net4932),
.A2(net4958),
.A3(net4901),
.A4(net4957),
.ZN(net10312)
);

SDFFS_X2 merge9471(
.D(net3594),
.SE(net3586),
.SI(net6336),
.SN(net5530),
.CK(clk),
.Q(net10314),
.QN(net10313)
);

SDFFR_X1 merge9472(
.D(net6841),
.RN(net7239),
.SE(net7850),
.SI(net7066),
.CK(clk),
.Q(net10316),
.QN(net10315)
);

AOI211_X1 merge9473(
.A(net1742),
.B(net1753),
.C1(net5532),
.C2(net5566),
.ZN(net10317)
);

SDFFR_X2 merge9474(
.D(net4383),
.RN(net3341),
.SE(net3117),
.SI(net5064),
.CK(clk),
.Q(net10319),
.QN(net10318)
);

SDFFS_X1 merge9475(
.D(net1415),
.SE(net617),
.SI(net3491),
.SN(net3470),
.CK(clk),
.Q(net10321),
.QN(net10320)
);

NAND4_X2 merge9476(
.A1(net2729),
.A2(net2605),
.A3(net817),
.A4(net778),
.ZN(net10322)
);

OR4_X4 merge9477(
.A1(net3277),
.A2(net3355),
.A3(net5048),
.A4(net5061),
.ZN(net10323)
);

SDFFS_X2 merge9478(
.D(net6390),
.SE(net6315),
.SI(net639),
.SN(net586),
.CK(clk),
.Q(net10325),
.QN(net10324)
);

SDFFR_X1 merge9479(
.D(net293),
.RN(net298),
.SE(net7040),
.SI(net7054),
.CK(clk),
.Q(net10327),
.QN(net10326)
);

OAI22_X2 merge9480(
.A1(net148),
.A2(net1940),
.B1(net284),
.B2(net1319),
.ZN(net10328)
);

SDFFR_X2 merge9481(
.D(net3193),
.RN(net3155),
.SE(net1790),
.SI(net1816),
.CK(clk),
.Q(net10330),
.QN(net10329)
);

SDFFS_X1 merge9482(
.D(net6846),
.SE(net7075),
.SI(net8046),
.SN(net6097),
.CK(clk),
.Q(net10332),
.QN(net10331)
);

SDFFS_X2 merge9483(
.D(net1527),
.SE(net4431),
.SI(net3160),
.SN(net2144),
.CK(clk),
.Q(net10334),
.QN(net10333)
);

OAI211_X4 merge9484(
.A(net3209),
.B(net3181),
.C1(net5393),
.C2(net7397),
.ZN(net10335)
);

OAI211_X1 merge9485(
.A(net5149),
.B(net8177),
.C1(net11326),
.C2(net11431),
.ZN(net10336)
);

SDFFR_X1 merge9486(
.D(net3762),
.RN(net3756),
.SE(net885),
.SI(net870),
.CK(clk),
.Q(net10338),
.QN(net10337)
);

NOR4_X4 merge9487(
.A1(net268),
.A2(net309),
.A3(net3524),
.A4(net2606),
.ZN(net10339)
);

SDFFR_X2 merge9488(
.D(net2351),
.RN(net2371),
.SE(net3443),
.SI(net1400),
.CK(clk),
.Q(net10341),
.QN(net10340)
);

NOR4_X2 merge9489(
.A1(net3270),
.A2(net4357),
.A3(net425),
.A4(net1391),
.ZN(net10342)
);

AOI211_X4 merge9490(
.A(net4397),
.B(net4306),
.C1(net8117),
.C2(net11558),
.ZN(net10343)
);

SDFFS_X1 merge9491(
.D(net7996),
.SE(net7792),
.SI(net8905),
.SN(net8016),
.CK(clk),
.Q(net10345),
.QN(net10344)
);

SDFFS_X2 merge9492(
.D(net921),
.SE(net890),
.SI(net6452),
.SN(net6265),
.CK(clk),
.Q(net10347),
.QN(net10346)
);

NOR4_X1 merge9493(
.A1(net118),
.A2(net3139),
.A3(net3379),
.A4(net3345),
.ZN(net10348)
);

SDFFR_X1 merge9494(
.D(net3490),
.RN(net3462),
.SE(net296),
.SI(net3022),
.CK(clk),
.Q(net10350),
.QN(net10349)
);

AOI211_X2 merge9495(
.A(net3688),
.B(net4640),
.C1(net4541),
.C2(net4590),
.ZN(net10351)
);

AOI22_X1 merge9496(
.A1(net2224),
.A2(net1236),
.B1(net3192),
.B2(net11279),
.ZN(net10352)
);

AND4_X4 merge9497(
.A1(net805),
.A2(net800),
.A3(net7197),
.A4(net6506),
.ZN(net10353)
);

SDFFR_X2 merge9498(
.D(net4557),
.RN(net5454),
.SE(net559),
.SI(net3604),
.CK(clk),
.Q(net10355),
.QN(net10354)
);

NAND4_X1 merge9499(
.A1(net3423),
.A2(net2514),
.A3(net5141),
.A4(net5149),
.ZN(net10356)
);

OR4_X1 merge9500(
.A1(net5390),
.A2(net5288),
.A3(net1109),
.A4(net2527),
.ZN(net10357)
);

SDFFS_X1 merge9501(
.D(net5103),
.SE(net3413),
.SI(net4393),
.SN(net4396),
.CK(clk),
.Q(net10359),
.QN(net10358)
);

SDFFS_X2 merge9502(
.D(net4518),
.SE(net4520),
.SI(net9107),
.SN(net9077),
.CK(clk),
.Q(net10361),
.QN(net10360)
);

SDFFR_X1 merge9503(
.D(net3118),
.RN(net235),
.SE(net2386),
.SI(net1465),
.CK(clk),
.Q(net10363),
.QN(net10362)
);

OAI22_X1 merge9504(
.A1(net5518),
.A2(net5501),
.B1(net7416),
.B2(net5482),
.ZN(net10364)
);

SDFFR_X2 merge9505(
.D(net3608),
.RN(net2633),
.SE(net4210),
.SI(net5112),
.CK(clk),
.Q(net10366),
.QN(net10365)
);

AND4_X2 merge9506(
.A1(net5069),
.A2(net4076),
.A3(net4214),
.A4(net4157),
.ZN(net10367)
);

SDFFS_X1 merge9507(
.D(net9049),
.SE(net9026),
.SI(net8864),
.SN(net8113),
.CK(clk),
.Q(net10369),
.QN(net10368)
);

SDFFS_X2 merge9508(
.D(net2541),
.SE(net2484),
.SI(net162),
.SN(net284),
.CK(clk),
.Q(net10371),
.QN(net10370)
);

SDFFR_X1 merge9509(
.D(net7190),
.RN(net6364),
.SE(net6681),
.SI(net6640),
.CK(clk),
.Q(net10373),
.QN(net10372)
);

SDFFR_X2 merge9510(
.D(net2878),
.RN(net3794),
.SE(net6414),
.SI(net5351),
.CK(clk),
.Q(net10375),
.QN(net10374)
);

AND4_X1 merge9511(
.A1(net2540),
.A2(net2142),
.A3(net277),
.A4(net274),
.ZN(net10376)
);

SDFFS_X1 merge9512(
.D(net6484),
.SE(net6277),
.SI(net1553),
.SN(net1698),
.CK(clk),
.Q(net10378),
.QN(net10377)
);

AOI22_X4 merge9513(
.A1(net1334),
.A2(net3256),
.B1(net3232),
.B2(net3235),
.ZN(net10379)
);

SDFFS_X2 merge9514(
.D(net1207),
.SE(net2172),
.SI(net3086),
.SN(net1053),
.CK(clk),
.Q(net10381),
.QN(net10380)
);

SDFFR_X1 merge9515(
.D(net5949),
.RN(net5953),
.SE(net2286),
.SI(net2294),
.CK(clk),
.Q(net10383),
.QN(net10382)
);

SDFFR_X2 merge9516(
.D(net925),
.RN(net774),
.SE(net4541),
.SI(net10780),
.CK(clk),
.Q(net10385),
.QN(net10384)
);

SDFFS_X1 merge9517(
.D(net4128),
.SE(net4108),
.SI(net5239),
.SN(net5307),
.CK(clk),
.Q(net10387),
.QN(net10386)
);

SDFFS_X2 merge9518(
.D(net4090),
.SE(net5226),
.SI(net5994),
.SN(net5933),
.CK(clk),
.Q(net10389),
.QN(net10388)
);

SDFFR_X1 merge9519(
.D(net6150),
.RN(net6212),
.SE(net4262),
.SI(net6870),
.CK(clk),
.Q(net10391),
.QN(net10390)
);

SDFFR_X2 merge9520(
.D(net4589),
.RN(net4566),
.SE(net4862),
.SI(net5277),
.CK(clk),
.Q(net10393),
.QN(net10392)
);

SDFFS_X1 merge9521(
.D(net8081),
.SE(net8187),
.SI(net4517),
.SN(net5542),
.CK(clk),
.Q(net10395),
.QN(net10394)
);

SDFFS_X2 merge9522(
.D(net8161),
.SE(net8155),
.SI(net6384),
.SN(net4642),
.CK(clk),
.Q(net10397),
.QN(net10396)
);

SDFFR_X1 merge9523(
.D(net763),
.RN(net2620),
.SE(net2469),
.SI(net3526),
.CK(clk),
.Q(net10399),
.QN(net10398)
);

SDFFR_X2 merge9524(
.D(net5460),
.RN(net5396),
.SE(net2778),
.SI(net932),
.CK(clk),
.Q(net10401),
.QN(net10400)
);

OAI22_X4 merge9525(
.A1(net4499),
.A2(net5317),
.B1(net3217),
.B2(net7302),
.ZN(net10402)
);

AOI22_X2 merge9526(
.A1(net6914),
.A2(net6989),
.B1(net1458),
.B2(net1484),
.ZN(net10403)
);

SDFFS_X1 merge9527(
.D(net6364),
.SE(net7397),
.SI(net5303),
.SN(net2509),
.CK(clk),
.Q(net10405),
.QN(net10404)
);

SDFFS_X2 merge9528(
.D(net1895),
.SE(net2814),
.SI(net5520),
.SN(net5515),
.CK(clk),
.Q(net10407),
.QN(net10406)
);

NAND4_X4 merge9529(
.A1(net1404),
.A2(net465),
.A3(net4178),
.A4(net4357),
.ZN(net10408)
);

SDFFR_X1 merge9530(
.D(net9061),
.RN(net9057),
.SE(net4234),
.SI(net1217),
.CK(clk),
.Q(net10410),
.QN(net10409)
);

SDFFR_X2 merge9531(
.D(net6459),
.RN(net5502),
.SE(net691),
.SI(net514),
.CK(clk),
.Q(net10412),
.QN(net10411)
);

OAI211_X2 merge9532(
.A(net7420),
.B(net7315),
.C1(net5534),
.C2(net5525),
.ZN(net10413)
);

SDFFS_X1 merge9533(
.D(net2702),
.SE(net2692),
.SI(net3247),
.SN(net2220),
.CK(clk),
.Q(net10415),
.QN(net10414)
);

SDFFS_X2 merge9534(
.D(net342),
.SE(net333),
.SI(net4011),
.SN(net4023),
.CK(clk),
.Q(net10417),
.QN(net10416)
);

SDFFR_X1 merge9535(
.D(net5274),
.RN(net8165),
.SE(net8150),
.SI(net11352),
.CK(clk),
.Q(net10419),
.QN(net10418)
);

OR4_X2 merge9536(
.A1(net5596),
.A2(net5655),
.A3(net489),
.A4(net875),
.ZN(net10420)
);

SDFFR_X2 merge9537(
.D(net6301),
.RN(net6327),
.SE(net5337),
.SI(net4404),
.CK(clk),
.Q(net10422),
.QN(net10421)
);

SDFFS_X1 merge9538(
.D(net3174),
.SE(net3192),
.SI(net2724),
.SN(net1791),
.CK(clk),
.Q(net10424),
.QN(net10423)
);

AOI211_X1 merge9539(
.A(net5396),
.B(net5258),
.C1(net4476),
.C2(net3582),
.ZN(net10425)
);

SDFFS_X2 merge9540(
.D(net2470),
.SE(net2572),
.SI(net6537),
.SN(net6542),
.CK(clk),
.Q(net10427),
.QN(net10426)
);

SDFFR_X1 merge9541(
.D(net879),
.RN(net4780),
.SE(net5443),
.SI(net5469),
.CK(clk),
.Q(net10429),
.QN(net10428)
);

SDFFR_X2 merge9542(
.D(net3413),
.RN(net4265),
.SE(net7264),
.SI(net6259),
.CK(clk),
.Q(net10431),
.QN(net10430)
);

SDFFS_X1 merge9543(
.D(net3355),
.SE(net4458),
.SI(net1708),
.SN(net1713),
.CK(clk),
.Q(net10433),
.QN(net10432)
);

NAND4_X2 merge9544(
.A1(net1680),
.A2(net1667),
.A3(net7324),
.A4(net10640),
.ZN(net10434)
);

SDFFS_X2 merge9545(
.D(net7892),
.SE(net7909),
.SI(net232),
.SN(net221),
.CK(clk),
.Q(net10436),
.QN(net10435)
);

OR4_X4 merge9546(
.A1(net7290),
.A2(net7292),
.A3(net8246),
.A4(net6292),
.ZN(net10437)
);

SDFFR_X1 merge9547(
.D(net6195),
.RN(net8366),
.SE(net6369),
.SI(net6177),
.CK(clk),
.Q(net10439),
.QN(net10438)
);

SDFFR_X2 merge9548(
.D(net8206),
.RN(net9118),
.SE(net3422),
.SI(net4298),
.CK(clk),
.Q(net10441),
.QN(net10440)
);

OAI22_X2 merge9549(
.A1(net2635),
.A2(net2728),
.B1(net582),
.B2(net576),
.ZN(net10442)
);

SDFFS_X1 merge9550(
.D(net5925),
.SE(net2016),
.SI(net4160),
.SN(net11376),
.CK(clk),
.Q(net10444),
.QN(net10443)
);

SDFFS_X2 merge9551(
.D(net3661),
.SE(net2589),
.SI(net4165),
.SN(net4163),
.CK(clk),
.Q(net10446),
.QN(net10445)
);

SDFFR_X1 merge9552(
.D(net6213),
.RN(net6150),
.SE(net7182),
.SI(net7169),
.CK(clk),
.Q(net10448),
.QN(net10447)
);

OAI211_X4 merge9553(
.A(net4180),
.B(net4102),
.C1(net3992),
.C2(net3981),
.ZN(net10449)
);

OAI211_X1 merge9554(
.A(net208),
.B(net188),
.C1(net3297),
.C2(net4160),
.ZN(net10450)
);

SDFFR_X2 merge9555(
.D(net6129),
.RN(net5135),
.SE(net3667),
.SI(net3709),
.CK(clk),
.Q(net10452),
.QN(net10451)
);

NOR4_X4 merge9556(
.A1(net6080),
.A2(net6043),
.A3(net7808),
.A4(net7850),
.ZN(net10453)
);

NOR4_X2 merge9557(
.A1(net4108),
.A2(net4112),
.A3(net231),
.A4(net215),
.ZN(net10454)
);

SDFFS_X1 merge9558(
.D(net5979),
.SE(net6912),
.SI(net6149),
.SN(net6182),
.CK(clk),
.Q(net10456),
.QN(net10455)
);

SDFFS_X2 merge9559(
.D(net1810),
.SE(net2724),
.SI(net7557),
.SN(net7525),
.CK(clk),
.Q(net10458),
.QN(net10457)
);

AOI211_X4 merge9560(
.A(net5301),
.B(net5250),
.C1(net5306),
.C2(net10977),
.ZN(net10459)
);

NOR4_X1 merge9561(
.A1(net1742),
.A2(net1817),
.A3(net3687),
.A4(net2605),
.ZN(net10460)
);

SDFFR_X1 merge9562(
.D(net7803),
.RN(net7910),
.SE(net8862),
.SI(net7812),
.CK(clk),
.Q(net10462),
.QN(net10461)
);

SDFFR_X2 merge9563(
.D(net3440),
.RN(net3397),
.SE(net5079),
.SI(net5094),
.CK(clk),
.Q(net10464),
.QN(net10463)
);

SDFFS_X1 merge9564(
.D(net2625),
.SE(net2712),
.SI(net5149),
.SN(net10795),
.CK(clk),
.Q(net10466),
.QN(net10465)
);

AOI211_X2 merge9565(
.A(net1292),
.B(net2256),
.C1(net3038),
.C2(net6944),
.ZN(net10467)
);

SDFFS_X2 merge9566(
.D(net3169),
.SE(net4210),
.SI(net4018),
.SN(net3038),
.CK(clk),
.Q(net10469),
.QN(net10468)
);

SDFFR_X1 merge9567(
.D(net489),
.RN(net1487),
.SE(net3471),
.SI(net11075),
.CK(clk),
.Q(net10471),
.QN(net10470)
);

SDFFR_X2 merge9568(
.D(net517),
.RN(net489),
.SE(net5081),
.SI(net5075),
.CK(clk),
.Q(net10473),
.QN(net10472)
);

SDFFS_X1 merge9569(
.D(net6273),
.SE(net7224),
.SI(net2184),
.SN(net2176),
.CK(clk),
.Q(net10475),
.QN(net10474)
);

SDFFS_X2 merge9570(
.D(net7074),
.SE(net7348),
.SI(net5389),
.SN(net6509),
.CK(clk),
.Q(net10477),
.QN(net10476)
);

AOI22_X1 merge9571(
.A1(net3648),
.A2(net2735),
.B1(net3764),
.B2(net3757),
.ZN(net10478)
);

AND4_X4 merge9572(
.A1(net4393),
.A2(net3383),
.A3(net2125),
.A4(net2958),
.ZN(net10479)
);

SDFFR_X1 merge9573(
.D(net3977),
.RN(net4094),
.SE(net3165),
.SI(net4135),
.CK(clk),
.Q(net10481),
.QN(net10480)
);

NAND4_X1 merge9574(
.A1(net233),
.A2(net1132),
.A3(net2254),
.A4(net3247),
.ZN(net10482)
);

SDFFR_X2 merge9575(
.D(net3710),
.RN(net2703),
.SE(net2417),
.SI(net11138),
.CK(clk),
.Q(net10484),
.QN(net10483)
);

OR4_X1 merge9576(
.A1(net4626),
.A2(net2772),
.A3(net8144),
.A4(net7940),
.ZN(net10485)
);

OAI22_X1 merge9577(
.A1(net2083),
.A2(net2126),
.B1(net6036),
.B2(net6028),
.ZN(net10486)
);

SDFFS_X1 merge9578(
.D(net3184),
.SE(net2987),
.SI(net3004),
.SN(net5153),
.CK(clk),
.Q(net10488),
.QN(net10487)
);

SDFFS_X2 merge9579(
.D(net1339),
.SE(net1397),
.SI(net6418),
.SN(net7533),
.CK(clk),
.Q(net10490),
.QN(net10489)
);

SDFFR_X1 merge9580(
.D(net8427),
.RN(net8346),
.SE(net2773),
.SI(net5586),
.CK(clk),
.Q(net10492),
.QN(net10491)
);

AND4_X2 merge9581(
.A1(net6467),
.A2(net6462),
.A3(net9170),
.A4(net8207),
.ZN(net10493)
);

SDFFR_X2 merge9582(
.D(net1713),
.RN(net2583),
.SE(net2585),
.SI(net11299),
.CK(clk),
.Q(net10495),
.QN(net10494)
);

AND4_X1 merge9583(
.A1(net1175),
.A2(net1162),
.A3(net2497),
.A4(net1541),
.ZN(net10496)
);

SDFFS_X1 merge9584(
.D(net6629),
.SE(net6628),
.SI(net5226),
.SN(net33),
.CK(clk),
.Q(net10498),
.QN(net10497)
);

SDFFS_X2 merge9585(
.D(net7170),
.SE(net7169),
.SI(net9111),
.SN(net8860),
.CK(clk),
.Q(net10500),
.QN(net10499)
);

SDFFR_X1 merge9586(
.D(net5934),
.RN(net3038),
.SE(net4028),
.SI(net3978),
.CK(clk),
.Q(net10502),
.QN(net10501)
);

SDFFR_X2 merge9587(
.D(net4967),
.RN(net5953),
.SE(net4004),
.SI(net6867),
.CK(clk),
.Q(net10504),
.QN(net10503)
);

NOR2_X1 merge9588(
.A1(net3367),
.A2(net3385),
.ZN(net10505)
);

DFFR_X1 merge9589(
.D(net3569),
.RN(net3583),
.CK(clk),
.Q(net10507),
.QN(net10506)
);

OR2_X2 merge9590(
.A1(net1398),
.A2(net1432),
.ZN(net10508)
);

DFFR_X2 merge9591(
.D(net426),
.RN(net452),
.CK(clk),
.Q(net10510),
.QN(net10509)
);

DFFS_X1 merge9592(
.D(net7736),
.SN(net7772),
.CK(clk),
.Q(net10512),
.QN(net10511)
);

DFFS_X2 merge9593(
.D(net8693),
.SN(net8740),
.CK(clk),
.Q(net10514),
.QN(net10513)
);

DFFR_X1 merge9594(
.D(net9381),
.RN(net9370),
.CK(clk),
.Q(net10516),
.QN(net10515)
);

DFFR_X2 merge9595(
.D(net8183),
.RN(net8216),
.CK(clk),
.Q(net10518),
.QN(net10517)
);

DFFS_X1 merge9596(
.D(net5679),
.SN(net5725),
.CK(clk),
.Q(net10520),
.QN(net10519)
);

DFFS_X2 merge9597(
.D(net7913),
.SN(net7917),
.CK(clk),
.Q(net10522),
.QN(net10521)
);

NOR2_X4 merge9598(
.A1(net1700),
.A2(net1714),
.ZN(net10523)
);

DFFR_X1 merge9599(
.D(net2573),
.RN(net2588),
.CK(clk),
.Q(net10525),
.QN(net10524)
);

NOR2_X2 merge9600(
.A1(net4351),
.A2(net4352),
.ZN(net10526)
);

XOR2_X2 merge9601(
.A(net8341),
.B(net8407),
.Z(net10527)
);

DFFR_X2 merge9602(
.D(net3711),
.RN(net3771),
.CK(clk),
.Q(net10529),
.QN(net10528)
);

DFFS_X1 merge9603(
.D(net319),
.Q(net10531),
.CK(clk),
.QN(net10530)
);

DFFS_X2 merge9604(
.D(net1929),
.SN(net1943),
.CK(clk),
.Q(net10533),
.QN(net10532)
);

DFFR_X1 merge9605(
.D(net60),
.RN(net92),
.CK(clk),
.Q(net10535),
.QN(net10534)
);

DFFR_X2 merge9606(
.D(net2835),
.RN(net2897),
.CK(clk),
.Q(net10537),
.QN(net10536)
);

DFFS_X1 merge9607(
.D(net1226),
.SN(net1233),
.CK(clk),
.Q(net10539),
.QN(net10538)
);

XNOR2_X1 merge9608(
.A(net738),
.B(net765),
.ZN(net10540)
);

DFFS_X2 merge9609(
.D(net9203),
.SN(net9289),
.CK(clk),
.Q(net10542),
.QN(net10541)
);

OR2_X4 merge9610(
.A1(net8621),
.A2(net8657),
.ZN(net10543)
);

DFFR_X1 merge9611(
.D(net5514),
.RN(net5526),
.CK(clk),
.Q(net10545),
.QN(net10544)
);

DFFR_X2 merge9612(
.D(net850),
.RN(net807),
.CK(clk),
.Q(net10547),
.QN(net10546)
);

DFFS_X1 merge9613(
.D(net7807),
.SN(net7799),
.CK(clk),
.Q(net10549),
.QN(net10548)
);

DFFS_X2 merge9614(
.D(net8821),
.Q(net8825),
.CK(clk),
.QN(net10550)
);

DFFR_X1 merge9615(
.D(net6882),
.RN(net9960),
.CK(clk),
.Q(net10553),
.QN(net10552)
);

DFFR_X2 merge9616(
.D(net9196),
.RN(net9177),
.CK(clk),
.Q(net10555),
.QN(net10554)
);

DFFS_X1 merge9617(
.D(net8504),
.SN(net8578),
.CK(clk),
.Q(net10557),
.QN(net10556)
);

DFFS_X2 merge9618(
.D(net5080),
.SN(net5087),
.CK(clk),
.Q(net10559),
.QN(net10558)
);

OR2_X1 merge9619(
.A1(net4427),
.A2(net4496),
.ZN(net10560)
);

DFFR_X1 merge9620(
.D(net5897),
.RN(net5906),
.CK(clk),
.Q(net10562),
.QN(net10561)
);

DFFR_X2 merge9621(
.D(net867),
.RN(net908),
.CK(clk),
.Q(net10564),
.QN(net10563)
);

DFFS_X1 merge9622(
.D(net8000),
.SN(net8006),
.CK(clk),
.Q(net10566),
.QN(net10565)
);

XNOR2_X2 merge9623(
.A(net1906),
.B(net1832),
.ZN(net10567)
);

AND2_X4 merge9624(
.A1(net650),
.A2(net676),
.ZN(net10568)
);

DFFS_X2 merge9625(
.D(net5244),
.SN(net5247),
.CK(clk),
.Q(net10570),
.QN(net10569)
);

DFFR_X1 merge9626(
.D(net7524),
.RN(net7554),
.CK(clk),
.Q(net10572),
.QN(net10571)
);

DFFR_X2 merge9627(
.D(net5435),
.RN(net5456),
.CK(clk),
.Q(net10574),
.QN(net10573)
);

AND2_X1 merge9628(
.A1(net9468),
.A2(net9466),
.ZN(net10575)
);

NAND2_X1 merge9629(
.A1(net2113),
.A2(net2116),
.ZN(net10576)
);

DFFS_X1 merge9630(
.D(net7002),
.SN(net7032),
.CK(clk),
.Q(net10578),
.QN(net10577)
);

NAND2_X2 merge9631(
.A1(net7090),
.A2(net7162),
.ZN(net10579)
);

DFFS_X2 merge9632(
.D(net5936),
.SN(net6013),
.CK(clk),
.Q(net10581),
.QN(net10580)
);

DFFR_X1 merge9633(
.D(net6392),
.RN(net6455),
.CK(clk),
.Q(net10583),
.QN(net10582)
);

DFFR_X2 merge9634(
.D(net2642),
.RN(net2645),
.CK(clk),
.Q(net10585),
.QN(net10584)
);

NAND2_X4 merge9635(
.A1(net3479),
.A2(net3482),
.ZN(net10586)
);

DFFS_X1 merge9636(
.D(net395),
.SN(net396),
.CK(clk),
.Q(net10588),
.QN(net10587)
);

DFFS_X2 merge9637(
.D(net9697),
.SN(net9961),
.CK(clk),
.Q(net10590),
.QN(net10589)
);

DFFR_X1 merge9638(
.D(net1819),
.RN(net1771),
.CK(clk),
.Q(net10592),
.QN(net10591)
);

DFFR_X2 merge9639(
.D(net5034),
.RN(net5001),
.CK(clk),
.Q(net10594),
.QN(net10593)
);

DFFS_X1 merge9640(
.D(net4801),
.SN(net4836),
.CK(clk),
.Q(net10596),
.QN(net10595)
);

DFFS_X2 merge9641(
.D(net8457),
.SN(net8453),
.CK(clk),
.Q(net10598),
.QN(net10597)
);

DFFR_X1 merge9642(
.D(net9481),
.RN(net9565),
.CK(clk),
.Q(net10600),
.QN(net10599)
);

DFFR_X2 merge9643(
.D(net9567),
.RN(net9642),
.CK(clk),
.Q(net10602),
.QN(net10601)
);

DFFS_X1 merge9644(
.D(net8298),
.SN(net8319),
.CK(clk),
.Q(net10604),
.QN(net10603)
);

DFFS_X2 merge9645(
.D(net6288),
.SN(net6324),
.CK(clk),
.Q(net10606),
.QN(net10605)
);

AND2_X2 merge9646(
.A1(net3664),
.A2(net3685),
.ZN(net10607)
);

XOR2_X1 merge9647(
.A(net1481),
.B(net1539),
.Z(net10608)
);

DFFR_X1 merge9648(
.D(net3088),
.RN(net3134),
.CK(clk),
.Q(net10610),
.QN(net10609)
);

NOR2_X1 merge9649(
.A1(net6233),
.A2(net6255),
.ZN(net10611)
);

OR2_X2 merge9650(
.A1(net4174),
.A2(net4179),
.ZN(net10612)
);

DFFR_X2 merge9651(
.D(net4594),
.RN(net4669),
.CK(clk),
.Q(net10614),
.QN(net10613)
);

DFFS_X1 merge9652(
.D(net4724),
.SN(net4725),
.CK(clk),
.Q(net10616),
.QN(net10615)
);

DFFS_X2 merge9653(
.D(net6916),
.SN(net6929),
.CK(clk),
.Q(net10618),
.QN(net10617)
);

NOR2_X4 merge9654(
.A1(net6579),
.A2(net6603),
.ZN(net10619)
);

NOR2_X2 merge9655(
.A1(net8119),
.A2(net8125),
.ZN(net10620)
);

XOR2_X2 merge9656(
.A(net2762),
.B(net2779),
.Z(net10621)
);

DFFR_X1 merge9657(
.D(net2071),
.RN(net2099),
.CK(clk),
.Q(net10623),
.QN(net10622)
);

XNOR2_X1 merge9658(
.A(net5155),
.B(net5161),
.ZN(net10624)
);

DFFR_X2 merge9659(
.D(net1013),
.RN(net1014),
.CK(clk),
.Q(net10626),
.QN(net10625)
);

DFFS_X1 merge9660(
.D(net9030),
.SN(net9099),
.CK(clk),
.Q(net10628),
.QN(net10627)
);

DFFS_X2 merge9661(
.D(net8929),
.SN(net8995),
.CK(clk),
.Q(net10630),
.QN(net10629)
);

DFFR_X1 merge9662(
.D(net5750),
.RN(net5762),
.CK(clk),
.Q(net10632),
.QN(net10631)
);

DFFR_X2 merge9663(
.D(net6661),
.RN(net6673),
.CK(clk),
.Q(net10634),
.QN(net10633)
);

DFFS_X1 merge9664(
.D(net4248),
.SN(net4255),
.CK(clk),
.Q(net10636),
.QN(net10635)
);

DFFS_X2 merge9665(
.D(net5570),
.SN(net5591),
.CK(clk),
.Q(net10638),
.QN(net10637)
);

DFFR_X1 merge9666(
.D(net7278),
.RN(net7305),
.CK(clk),
.Q(net10640),
.QN(net10639)
);

DFFR_X2 merge9667(
.D(net217),
.RN(net222),
.CK(clk),
.Q(net10642),
.QN(net10641)
);

DFFS_X1 merge9668(
.D(net3887),
.SN(net3891),
.CK(clk),
.Q(net10644),
.QN(net10643)
);

OR2_X4 merge9669(
.A1(net6155),
.A2(net6174),
.ZN(net10645)
);

OR2_X1 merge9670(
.A1(net7369),
.A2(net7368),
.ZN(net10646)
);

XNOR2_X2 merge9671(
.A(net1608),
.B(net1614),
.ZN(net10647)
);

DFFS_X2 merge9672(
.D(net2994),
.SN(net2949),
.CK(clk),
.Q(net10649),
.QN(net10648)
);

AND2_X4 merge9673(
.A1(net7429),
.A2(net7437),
.ZN(net10650)
);

DFFR_X1 merge9674(
.D(net6084),
.RN(net6089),
.CK(clk),
.Q(net10652),
.QN(net10651)
);

DFFR_X2 merge9675(
.D(net7643),
.RN(net7645),
.CK(clk),
.Q(net10654),
.QN(net10653)
);

AND2_X1 merge9676(
.A1(net3273),
.A2(net3351),
.ZN(net10655)
);

DFFS_X1 merge9677(
.D(net6479),
.SN(net6527),
.CK(clk),
.Q(net10657),
.QN(net10656)
);

NAND2_X1 merge9678(
.A1(net2193),
.A2(net2228),
.ZN(net10658)
);

NAND2_X2 merge9679(
.A1(net4120),
.A2(net4077),
.ZN(net10659)
);

DFFS_X2 merge9680(
.D(net3018),
.SN(net3033),
.CK(clk),
.Q(net10661),
.QN(net10660)
);

DFFR_X1 merge9681(
.D(net2384),
.RN(net2372),
.CK(clk),
.Q(net10663),
.QN(net10662)
);

DFFR_X2 merge9682(
.D(net4921),
.RN(net4927),
.CK(clk),
.Q(net10665),
.QN(net10664)
);

NAND2_X4 merge9683(
.A1(net1196),
.A2(net1198),
.ZN(net10666)
);

DFFS_X1 merge9684(
.D(net3986),
.SN(net4006),
.CK(clk),
.Q(net10668),
.QN(net10667)
);

AND2_X2 merge9685(
.A1(net1032),
.A2(net1114),
.ZN(net10669)
);

DFFS_X2 merge9686(
.D(net7179),
.SN(net7223),
.CK(clk),
.Q(net10671),
.QN(net10670)
);

XOR2_X1 merge9687(
.A(net3197),
.B(net3186),
.Z(net10672)
);

DFFR_X1 merge9688(
.D(net3790),
.RN(net3786),
.CK(clk),
.Q(net10674),
.QN(net10673)
);

NOR2_X1 merge9689(
.A1(net5324),
.A2(net5385),
.ZN(net10675)
);

DFFR_X2 merge9690(
.D(net4502),
.RN(net4527),
.CK(clk),
.Q(net10677),
.QN(net10676)
);

DFFS_X1 merge9691(
.D(net6768),
.SN(net6795),
.CK(clk),
.Q(net10679),
.QN(net10678)
);

DFFS_X2 merge9692(
.D(net8856),
.SN(net8916),
.CK(clk),
.Q(net10681),
.QN(net10680)
);

DFFR_X1 merge9693(
.D(net544),
.RN(net547),
.CK(clk),
.Q(net10683),
.QN(net10682)
);

OR2_X2 merge9694(
.A1(net1337),
.A2(net1347),
.ZN(net10684)
);

NOR2_X4 merge9695(
.A1(net2302),
.A2(net2319),
.ZN(net10685)
);

DFFR_X2 merge9696(
.D(net4039),
.RN(net3152),
.CK(clk),
.Q(net10687),
.QN(net10686)
);

NOR2_X2 merge9697(
.A1(net4480),
.A2(net3404),
.ZN(net10688)
);

DFFS_X1 merge9698(
.D(net9590),
.SN(net9634),
.CK(clk),
.Q(net10690),
.QN(net10689)
);

DFFS_X2 merge9699(
.D(net2010),
.SN(net1098),
.CK(clk),
.Q(net10692),
.QN(net10691)
);

DFFR_X1 merge9700(
.D(net4225),
.RN(net4054),
.CK(clk),
.Q(net10694),
.QN(net10693)
);

DFFR_X2 merge9701(
.D(net1199),
.RN(net10328),
.CK(clk),
.Q(net10696),
.QN(net10695)
);

DFFS_X1 merge9702(
.D(net1641),
.SN(net1634),
.CK(clk),
.Q(net10698),
.QN(net10697)
);

DFFS_X2 merge9703(
.D(net1974),
.SN(net2004),
.CK(clk),
.Q(net10700),
.QN(net10699)
);

XOR2_X2 merge9704(
.A(net2631),
.B(net1533),
.Z(net10701)
);

XNOR2_X1 merge9705(
.A(net3755),
.B(net2800),
.ZN(net10702)
);

OR2_X4 merge9706(
.A1(net1507),
.A2(net1559),
.ZN(net10703)
);

DFFR_X1 merge9707(
.D(net1026),
.RN(net10669),
.CK(clk),
.Q(net10705),
.QN(net10704)
);

OR2_X1 merge9708(
.A1(net3260),
.A2(net2262),
.ZN(net10706)
);

DFFR_X2 merge9709(
.D(net4760),
.RN(net4838),
.CK(clk),
.Q(net10708),
.QN(net10707)
);

XNOR2_X2 merge9710(
.A(net3415),
.B(net3205),
.ZN(net10709)
);

DFFS_X1 merge9711(
.D(net1952),
.SN(net3082),
.CK(clk),
.Q(net10711),
.QN(net10710)
);

DFFS_X2 merge9712(
.D(net8602),
.SN(net8624),
.CK(clk),
.Q(net10713),
.QN(net10712)
);

DFFR_X1 merge9713(
.D(net3893),
.RN(net4056),
.CK(clk),
.Q(net10715),
.QN(net10714)
);

DFFR_X2 merge9714(
.D(net8397),
.RN(net8499),
.CK(clk),
.Q(net10717),
.QN(net10716)
);

DFFS_X1 merge9715(
.D(net9605),
.SN(net8713),
.CK(clk),
.Q(net10718),
.QN(out4)
);

DFFS_X2 merge9716(
.D(net7481),
.SN(net7330),
.CK(clk),
.Q(net10720),
.QN(net10719)
);

DFFR_X1 merge9717(
.D(net8476),
.RN(net8558),
.CK(clk),
.Q(net10722),
.QN(net10721)
);

DFFR_X2 merge9718(
.D(net7722),
.RN(net8598),
.CK(clk),
.Q(net10724),
.QN(net10723)
);

DFFS_X1 merge9719(
.D(net3519),
.SN(net3409),
.CK(clk),
.Q(net10726),
.QN(net10725)
);

DFFS_X2 merge9720(
.D(net3447),
.SN(net2452),
.CK(clk),
.Q(net10728),
.QN(net10727)
);

AND2_X4 merge9721(
.A1(net4216),
.A2(net2239),
.ZN(net10729)
);

DFFR_X1 merge9722(
.D(net5943),
.RN(net6973),
.CK(clk),
.Q(net10731),
.QN(net10730)
);

AND2_X1 merge9723(
.A1(net7101),
.A2(net7163),
.ZN(net10732)
);

NAND2_X1 merge9724(
.A1(net2258),
.A2(net3208),
.ZN(net10733)
);

DFFR_X2 merge9725(
.D(net7158),
.RN(net7120),
.CK(clk),
.Q(net10735),
.QN(net10734)
);

NAND2_X2 merge9726(
.A1(net2365),
.A2(net3514),
.ZN(net10736)
);

NAND2_X4 merge9727(
.A1(net3971),
.A2(net5029),
.ZN(net10737)
);

DFFS_X1 merge9728(
.D(net3869),
.SN(net4778),
.CK(clk),
.Q(net10739),
.QN(net10738)
);

DFFS_X2 merge9729(
.D(net7683),
.SN(net7712),
.CK(clk),
.Q(net10741),
.QN(net10740)
);

DFFR_X1 merge9730(
.D(net8159),
.RN(net9071),
.CK(clk),
.Q(net10743),
.QN(net10742)
);

DFFR_X2 merge9731(
.D(net5359),
.RN(net4567),
.CK(clk),
.Q(net10745),
.QN(net10744)
);

DFFS_X1 merge9732(
.D(net5984),
.SN(net7880),
.CK(clk),
.Q(net10747),
.QN(net10746)
);

DFFS_X2 merge9733(
.D(net5197),
.SN(net4305),
.CK(clk),
.Q(net10749),
.QN(net10748)
);

DFFR_X1 merge9734(
.D(net8221),
.RN(net7232),
.CK(clk),
.Q(net10751),
.QN(net10750)
);

DFFR_X2 merge9735(
.D(net6802),
.RN(net5728),
.CK(clk),
.Q(net10753),
.QN(net10752)
);

AND2_X2 merge9736(
.A1(net7410),
.A2(net8351),
.ZN(net10754)
);

XOR2_X1 merge9737(
.A(net2150),
.B(net1290),
.Z(net10755)
);

DFFS_X1 merge9738(
.D(net1884),
.SN(net1898),
.CK(clk),
.Q(net10757),
.QN(net10756)
);

DFFS_X2 merge9739(
.D(net470),
.SN(net1472),
.CK(clk),
.Q(net10759),
.QN(net10758)
);

NOR2_X1 merge9740(
.A1(net2419),
.A2(net2283),
.ZN(net10760)
);

DFFR_X1 merge9741(
.D(net8949),
.RN(net8037),
.CK(clk),
.Q(net10762),
.QN(net10761)
);

DFFR_X2 merge9742(
.D(net4041),
.RN(net4017),
.CK(clk),
.Q(net10764),
.QN(net10763)
);

DFFS_X1 merge9743(
.D(net9306),
.SN(net9383),
.CK(clk),
.Q(net10766),
.QN(net10765)
);

DFFS_X2 merge9744(
.D(net5281),
.SN(net3335),
.CK(clk),
.Q(net10768),
.QN(net10767)
);

DFFR_X1 merge9745(
.D(net8136),
.RN(net8914),
.CK(clk),
.Q(net10770),
.QN(net10769)
);

DFFR_X2 merge9746(
.D(net7484),
.RN(net5633),
.CK(clk),
.Q(net10772),
.QN(net10771)
);

DFFS_X1 merge9747(
.D(net1889),
.SN(net937),
.CK(clk),
.Q(net10774),
.QN(net10773)
);

OR2_X2 merge9748(
.A1(net1876),
.A2(net930),
.ZN(net10775)
);

NOR2_X4 merge9749(
.A1(net2324),
.A2(net2364),
.ZN(net10776)
);

DFFS_X2 merge9750(
.D(net4772),
.SN(net6750),
.CK(clk),
.Q(net10778),
.QN(net10777)
);

DFFR_X1 merge9751(
.D(net4576),
.RN(net4601),
.CK(clk),
.Q(net10780),
.QN(net10779)
);

NOR2_X2 merge9752(
.A1(net1285),
.A2(net2159),
.ZN(net10781)
);

XOR2_X2 merge9753(
.A(net2674),
.B(net2718),
.Z(net10782)
);

XNOR2_X1 merge9754(
.A(net8488),
.B(net6708),
.ZN(net10783)
);

OR2_X4 merge9755(
.A1(net1511),
.A2(net1459),
.ZN(net10784)
);

DFFR_X2 merge9756(
.D(net8915),
.RN(net6986),
.CK(clk),
.Q(net10786),
.QN(net10785)
);

DFFS_X1 merge9757(
.D(net2845),
.SN(net2888),
.CK(clk),
.Q(net10788),
.QN(net10787)
);

DFFS_X2 merge9758(
.D(net6366),
.SN(net6415),
.CK(clk),
.Q(net10790),
.QN(net10789)
);

OR2_X1 merge9759(
.A1(net2160),
.A2(net1380),
.ZN(net10791)
);

XNOR2_X2 merge9760(
.A(net7601),
.B(net7498),
.ZN(net10792)
);

DFFR_X1 merge9761(
.D(net3804),
.RN(net4648),
.CK(clk),
.Q(net10794),
.QN(net10793)
);

DFFR_X2 merge9762(
.D(net4190),
.RN(net4230),
.CK(clk),
.Q(net10796),
.QN(net10795)
);

DFFS_X1 merge9763(
.D(net5007),
.SN(net4145),
.CK(clk),
.Q(net10798),
.QN(net10797)
);

AND2_X4 merge9764(
.A1(net4533),
.A2(net6377),
.ZN(net10799)
);

AND2_X1 merge9765(
.A1(net5348),
.A2(net5178),
.ZN(net10800)
);

NAND2_X1 merge9766(
.A1(net4654),
.A2(net2667),
.ZN(net10801)
);

DFFS_X2 merge9767(
.D(net6443),
.SN(net5376),
.CK(clk),
.Q(net10803),
.QN(net10802)
);

DFFR_X1 merge9768(
.D(net936),
.RN(net1905),
.CK(clk),
.Q(net10805),
.QN(net10804)
);

DFFR_X2 merge9769(
.D(net2627),
.RN(net3515),
.CK(clk),
.Q(net10807),
.QN(net10806)
);

DFFS_X1 merge9770(
.D(net8643),
.SN(net8620),
.CK(clk),
.Q(net10809),
.QN(net10808)
);

DFFS_X2 merge9771(
.D(net4855),
.SN(net6605),
.CK(clk),
.Q(net10811),
.QN(net10810)
);

NAND2_X2 merge9772(
.A1(net6326),
.A2(net7116),
.ZN(net10812)
);

DFFR_X1 merge9773(
.D(net8828),
.RN(net8910),
.CK(clk),
.Q(net10814),
.QN(net10813)
);

DFFR_X2 merge9774(
.D(net6935),
.RN(net7973),
.CK(clk),
.Q(net10816),
.QN(net10815)
);

DFFS_X1 merge9775(
.D(net9350),
.SN(net8503),
.CK(clk),
.Q(net10818),
.QN(net10817)
);

NAND2_X4 merge9776(
.A1(net8324),
.A2(net9157),
.ZN(net10819)
);

DFFS_X2 merge9777(
.D(net2168),
.SN(net3070),
.CK(clk),
.Q(net10821),
.QN(net10820)
);

AND2_X2 merge9778(
.A1(net4543),
.A2(net5643),
.ZN(net10822)
);

DFFR_X1 merge9779(
.D(net6692),
.RN(net6460),
.CK(clk),
.Q(net10824),
.QN(net10823)
);

XOR2_X1 merge9780(
.A(net4622),
.B(net2699),
.Z(net10825)
);

DFFR_X2 merge9781(
.D(net1267),
.RN(net10018),
.CK(clk),
.Q(net10827),
.QN(net10826)
);

DFFS_X1 merge9782(
.D(net7114),
.SN(net6190),
.CK(clk),
.Q(net10829),
.QN(net10828)
);

DFFS_X2 merge9783(
.D(net6941),
.SN(net5011),
.CK(clk),
.Q(net10831),
.QN(net10830)
);

DFFR_X1 merge9784(
.D(net405),
.RN(net9864),
.CK(clk),
.Q(net10833),
.QN(net10832)
);

NOR2_X1 merge9785(
.A1(net3211),
.A2(net3255),
.ZN(net10834)
);

DFFR_X2 merge9786(
.D(net6977),
.RN(net8909),
.CK(clk),
.Q(net10836),
.QN(net10835)
);

DFFS_X1 merge9787(
.D(net6806),
.SN(net7658),
.CK(clk),
.Q(net10838),
.QN(net10837)
);

DFFS_X2 merge9788(
.D(net1441),
.SN(net1366),
.CK(clk),
.Q(net10840),
.QN(net10839)
);

OR2_X2 merge9789(
.A1(net7337),
.A2(net9185),
.ZN(net10841)
);

NOR2_X4 merge9790(
.A1(net9004),
.A2(net9133),
.ZN(net10842)
);

DFFR_X1 merge9791(
.D(net5546),
.RN(net6411),
.CK(clk),
.Q(net10844),
.QN(net10843)
);

DFFR_X2 merge9792(
.D(net4799),
.RN(net5767),
.CK(clk),
.Q(net10846),
.QN(net10845)
);

NOR2_X2 merge9793(
.A1(net9171),
.A2(net7307),
.ZN(net10847)
);

XOR2_X2 merge9794(
.A(net1509),
.B(net1537),
.Z(net10848)
);

XNOR2_X1 merge9795(
.A(net5199),
.B(net4226),
.ZN(net10849)
);

OR2_X4 merge9796(
.A1(net6361),
.A2(net5251),
.ZN(net10850)
);

DFFS_X1 merge9797(
.D(net7094),
.SN(net8028),
.CK(clk),
.Q(net10852),
.QN(net10851)
);

DFFS_X2 merge9798(
.D(net3766),
.SN(net2714),
.CK(clk),
.Q(net10854),
.QN(net10853)
);

DFFR_X1 merge9799(
.D(net8626),
.RN(net8670),
.CK(clk),
.Q(net10856),
.QN(net10855)
);

DFFR_X2 merge9800(
.D(net2233),
.RN(net2453),
.CK(clk),
.Q(net10858),
.QN(net10857)
);

DFFS_X1 merge9801(
.D(net5099),
.SN(net7129),
.CK(clk),
.Q(net10860),
.QN(net10859)
);

OR2_X1 merge9802(
.A1(net5088),
.A2(net6275),
.ZN(net10861)
);

DFFS_X2 merge9803(
.D(net9454),
.SN(net7679),
.CK(clk),
.Q(net10863),
.QN(net10862)
);

XNOR2_X2 merge9804(
.A(net8234),
.B(net8139),
.ZN(net10864)
);

DFFR_X1 merge9805(
.D(net1992),
.RN(net2032),
.CK(clk),
.Q(net10866),
.QN(net10865)
);

AND2_X4 merge9806(
.A1(net8053),
.A2(net7058),
.ZN(net10867)
);

DFFR_X2 merge9807(
.D(net9237),
.RN(net9255),
.CK(clk),
.Q(net10869),
.QN(net10868)
);

DFFS_X1 merge9808(
.D(net9563),
.SN(net6748),
.CK(clk),
.Q(net10871),
.QN(net10870)
);

AND2_X1 merge9809(
.A1(net5172),
.A2(net4471),
.ZN(net10872)
);

DFFS_X2 merge9810(
.D(net2397),
.SN(net1615),
.CK(clk),
.Q(net10874),
.QN(net10873)
);

DFFR_X1 merge9811(
.D(net4564),
.RN(net3605),
.CK(clk),
.Q(net10876),
.QN(net10875)
);

DFFR_X2 merge9812(
.D(net1873),
.RN(net3861),
.CK(clk),
.Q(net10878),
.QN(net10877)
);

DFFS_X1 merge9813(
.D(net3957),
.SN(net3956),
.CK(clk),
.Q(net10880),
.QN(net10879)
);

DFFS_X2 merge9814(
.D(net2872),
.SN(net4825),
.CK(clk),
.Q(net10882),
.QN(net10881)
);

DFFR_X1 merge9815(
.D(net5349),
.RN(net7425),
.CK(clk),
.Q(net10884),
.QN(net10883)
);

DFFR_X2 merge9816(
.D(net4223),
.RN(net3262),
.CK(clk),
.Q(net10886),
.QN(net10885)
);

NAND2_X1 merge9817(
.A1(net6092),
.A2(net8936),
.ZN(net10887)
);

DFFS_X1 merge9818(
.D(net5957),
.SN(net6003),
.CK(clk),
.Q(net10889),
.QN(net10888)
);

DFFS_X2 merge9819(
.D(net7423),
.SN(net9091),
.CK(clk),
.Q(net10891),
.QN(net10890)
);

DFFR_X1 merge9820(
.D(net10106),
.RN(net10450),
.CK(clk),
.Q(net10893),
.QN(net10892)
);

NAND2_X2 merge9821(
.A1(net7057),
.A2(net7070),
.ZN(net10894)
);

NAND2_X4 merge9822(
.A1(net8970),
.A2(net8036),
.ZN(net10895)
);

DFFR_X2 merge9823(
.D(net8148),
.RN(net7145),
.CK(clk),
.Q(net10897),
.QN(net10896)
);

DFFS_X1 merge9824(
.D(net4388),
.SN(net4224),
.CK(clk),
.Q(net10899),
.QN(net10898)
);

DFFS_X2 merge9825(
.D(net4744),
.SN(net4616),
.CK(clk),
.Q(net10901),
.QN(net10900)
);

DFFR_X1 merge9826(
.D(net4965),
.RN(net5122),
.CK(clk),
.Q(net10903),
.QN(net10902)
);

DFFR_X2 merge9827(
.D(net5781),
.RN(net3796),
.CK(clk),
.Q(net10905),
.QN(net10904)
);

AND2_X2 merge9828(
.A1(net5116),
.A2(net5293),
.ZN(net10906)
);

XOR2_X1 merge9829(
.A(net6179),
.B(net5192),
.Z(net10907)
);

NOR2_X1 merge9830(
.A1(net3701),
.A2(net3417),
.ZN(net10908)
);

DFFS_X1 merge9831(
.D(net9329),
.SN(net9160),
.CK(clk),
.Q(net10910),
.QN(net10909)
);

DFFS_X2 merge9832(
.D(net8146),
.SN(net5189),
.CK(clk),
.Q(net10912),
.QN(net10911)
);

DFFR_X1 merge9833(
.D(net8653),
.RN(net9512),
.CK(clk),
.Q(net10914),
.QN(net10913)
);

OR2_X2 merge9834(
.A1(net2337),
.A2(net2330),
.ZN(net10915)
);

NOR2_X4 merge9835(
.A1(net9541),
.A2(net9564),
.ZN(net10916)
);

NOR2_X2 merge9836(
.A1(net5554),
.A2(net6355),
.ZN(net10917)
);

DFFR_X2 merge9837(
.D(net7104),
.RN(net7110),
.CK(clk),
.Q(net10919),
.QN(net10918)
);

DFFS_X1 merge9838(
.D(net8404),
.SN(net6524),
.CK(clk),
.Q(net10921),
.QN(net10920)
);

XOR2_X2 merge9839(
.A(net8976),
.B(net8904),
.Z(net10922)
);

DFFS_X2 merge9840(
.D(net6005),
.SN(net6334),
.CK(clk),
.Q(net10924),
.QN(net10923)
);

XNOR2_X1 merge9841(
.A(net8954),
.B(net9172),
.ZN(net10925)
);

DFFR_X1 merge9842(
.D(net9056),
.RN(net9140),
.CK(clk),
.Q(net10927),
.QN(net10926)
);

OR2_X4 merge9843(
.A1(net5271),
.A2(net4485),
.ZN(net10928)
);

DFFR_X2 merge9844(
.D(net1847),
.RN(net1869),
.CK(clk),
.Q(net10930),
.QN(net10929)
);

DFFS_X1 merge9845(
.D(net2082),
.SN(net9844),
.CK(clk),
.Q(net10932),
.QN(net10931)
);

OR2_X1 merge9846(
.A1(net4415),
.A2(net4315),
.ZN(net10933)
);

XNOR2_X2 merge9847(
.A(net9455),
.B(net8676),
.ZN(net10934)
);

DFFS_X2 merge9848(
.D(net8687),
.SN(net4849),
.CK(clk),
.Q(net10936),
.QN(net10935)
);

DFFR_X1 merge9849(
.D(net6770),
.RN(net6784),
.CK(clk),
.Q(net10938),
.QN(net10937)
);

DFFR_X2 merge9850(
.D(net8494),
.RN(net8574),
.CK(clk),
.Q(net10940),
.QN(net10939)
);

DFFS_X1 merge9851(
.D(net5790),
.SN(net8665),
.CK(clk),
.Q(net10942),
.QN(net10941)
);

DFFS_X2 merge9852(
.D(net413),
.SN(net2267),
.CK(clk),
.Q(net10944),
.QN(net10943)
);

DFFR_X1 merge9853(
.D(net2803),
.RN(net6760),
.CK(clk),
.Q(net10946),
.QN(net10945)
);

DFFR_X2 merge9854(
.D(net2694),
.RN(net2690),
.CK(clk),
.Q(net10948),
.QN(net10947)
);

DFFS_X1 merge9855(
.D(net3853),
.SN(net4432),
.CK(clk),
.Q(net10950),
.QN(net10949)
);

DFFS_X2 merge9856(
.D(net4236),
.SN(net4319),
.CK(clk),
.Q(net10952),
.QN(net10951)
);

DFFR_X1 merge9857(
.D(net6778),
.RN(net5636),
.CK(clk),
.Q(net10954),
.QN(net10953)
);

DFFR_X2 merge9858(
.D(net7556),
.RN(net9453),
.CK(clk),
.Q(net10956),
.QN(net10955)
);

DFFS_X1 merge9859(
.D(net9414),
.SN(net9266),
.CK(clk),
.Q(net10958),
.QN(net10957)
);

DFFS_X2 merge9860(
.D(net10791),
.SN(net2151),
.CK(clk),
.Q(net10960),
.QN(net10959)
);

AND2_X4 merge9861(
.A1(net7237),
.A2(net7323),
.ZN(net10961)
);

DFFR_X1 merge9862(
.D(net8611),
.RN(net9558),
.CK(clk),
.Q(net10963),
.QN(net10962)
);

DFFR_X2 merge9863(
.D(net3400),
.RN(net10008),
.CK(clk),
.Q(net10965),
.QN(net10964)
);

DFFS_X1 merge9864(
.D(net8980),
.SN(net7967),
.CK(clk),
.Q(net10967),
.QN(net10966)
);

DFFS_X2 merge9865(
.D(net5096),
.SN(net5115),
.CK(clk),
.Q(net10969),
.QN(net10968)
);

DFFR_X1 merge9866(
.D(net4629),
.RN(net5350),
.CK(clk),
.Q(net10971),
.QN(net10970)
);

DFFR_X2 merge9867(
.D(net5814),
.RN(net4621),
.CK(clk),
.Q(net10973),
.QN(net10972)
);

DFFS_X1 merge9868(
.D(net9084),
.SN(net9139),
.CK(clk),
.Q(net10975),
.QN(net10974)
);

DFFS_X2 merge9869(
.D(net5342),
.SN(net9201),
.CK(clk),
.Q(net10977),
.QN(net10976)
);

DFFR_X1 merge9870(
.D(net6441),
.RN(net7596),
.CK(clk),
.Q(net10979),
.QN(net10978)
);

DFFR_X2 merge9871(
.D(net9278),
.RN(net9239),
.CK(clk),
.Q(net10981),
.QN(net10980)
);

DFFS_X1 merge9872(
.D(net4749),
.SN(net6360),
.CK(clk),
.Q(net10983),
.QN(net10982)
);

DFFS_X2 merge9873(
.D(net3502),
.SN(net3495),
.CK(clk),
.Q(net10985),
.QN(net10984)
);

DFFR_X1 merge9874(
.D(net6521),
.RN(net6426),
.CK(clk),
.Q(net10987),
.QN(net10986)
);

DFFR_X2 merge9875(
.D(net9554),
.RN(net9479),
.CK(clk),
.Q(net10989),
.QN(net10988)
);

DFFS_X1 merge9876(
.D(net2864),
.SN(net1826),
.CK(clk),
.Q(net10991),
.QN(net10990)
);

DFFS_X2 merge9877(
.D(net7701),
.SN(net6805),
.CK(clk),
.Q(net10993),
.QN(net10992)
);

DFFR_X1 merge9878(
.D(net7699),
.RN(net9601),
.CK(clk),
.Q(out15),
.QN(net10994)
);

DFFR_X2 merge9879(
.D(net1897),
.RN(net3877),
.CK(clk),
.Q(net10996),
.QN(net10995)
);

AND2_X1 merge9880(
.A1(net6622),
.A2(net5743),
.ZN(net10997)
);

DFFS_X1 merge9881(
.D(net9566),
.SN(net7775),
.CK(clk),
.Q(net10999),
.QN(net10998)
);

DFFS_X2 merge9882(
.D(net8606),
.SN(net9569),
.CK(clk),
.Q(net11001),
.QN(net11000)
);

DFFR_X1 merge9883(
.D(net10339),
.RN(net10486),
.CK(clk),
.Q(net11003),
.QN(net11002)
);

DFFR_X2 merge9884(
.D(net10701),
.RN(net10647),
.CK(clk),
.Q(net11005),
.QN(net11004)
);

DFFS_X1 merge9885(
.D(net9380),
.SN(net8350),
.CK(clk),
.Q(net11007),
.QN(net11006)
);

DFFS_X2 merge9886(
.D(net9073),
.SN(net5992),
.CK(clk),
.Q(net11009),
.QN(net11008)
);

DFFR_X1 merge9887(
.D(net6006),
.RN(net10224),
.CK(clk),
.Q(net11011),
.QN(net11010)
);

NAND2_X1 merge9888(
.A1(net4584),
.A2(net5336),
.ZN(net11012)
);

DFFR_X2 merge9889(
.D(net7143),
.RN(net7322),
.CK(clk),
.Q(net11014),
.QN(net11013)
);

DFFS_X1 merge9890(
.D(net10408),
.SN(net481),
.CK(clk),
.Q(net11016),
.QN(net11015)
);

DFFS_X2 merge9891(
.D(net658),
.SN(net10376),
.CK(clk),
.Q(net11018),
.QN(net11017)
);

DFFR_X1 merge9892(
.D(net10312),
.RN(net10737),
.CK(clk),
.Q(net11020),
.QN(net11019)
);

DFFR_X2 merge9893(
.D(net6399),
.RN(net6279),
.CK(clk),
.Q(net11022),
.QN(net11021)
);

DFFS_X1 merge9894(
.D(net4815),
.SN(net4809),
.CK(clk),
.Q(net11024),
.QN(net11023)
);

DFFS_X2 merge9895(
.D(net9074),
.SN(net9024),
.CK(clk),
.Q(net11026),
.QN(net11025)
);

DFFR_X1 merge9896(
.D(net8230),
.RN(net8367),
.CK(clk),
.Q(net11028),
.QN(net11027)
);

NAND2_X2 merge9897(
.A1(net9195),
.A2(net9267),
.ZN(net11029)
);

DFFR_X2 merge9898(
.D(net10012),
.RN(net3693),
.CK(clk),
.Q(net11031),
.QN(net11030)
);

DFFS_X1 merge9899(
.D(net9114),
.SN(net9183),
.CK(clk),
.Q(net11033),
.QN(net11032)
);

DFFS_X2 merge9900(
.D(net6783),
.SN(net5823),
.CK(clk),
.Q(net11035),
.QN(net11034)
);

NAND2_X4 merge9901(
.A1(net9451),
.A2(net9543),
.ZN(net11036)
);

DFFR_X1 merge9902(
.D(net4560),
.RN(net4759),
.CK(clk),
.Q(net11038),
.QN(net11037)
);

DFFR_X2 merge9903(
.D(net10849),
.RN(net10684),
.CK(clk),
.Q(net11040),
.QN(net11039)
);

DFFS_X1 merge9904(
.D(net9037),
.SN(net9105),
.CK(clk),
.Q(net11042),
.QN(net11041)
);

DFFS_X2 merge9905(
.D(net572),
.SN(net10116),
.CK(clk),
.Q(net11044),
.QN(net11043)
);

DFFR_X1 merge9906(
.D(net6686),
.RN(net5735),
.CK(clk),
.Q(net11046),
.QN(net11045)
);

DFFR_X2 merge9907(
.D(net10004),
.RN(net10576),
.CK(clk),
.Q(net11048),
.QN(net11047)
);

DFFS_X1 merge9908(
.D(net6969),
.SN(net10052),
.CK(clk),
.Q(net11050),
.QN(net11049)
);

DFFS_X2 merge9909(
.D(net10132),
.SN(net10322),
.CK(clk),
.Q(net11052),
.QN(net11051)
);

DFFR_X1 merge9910(
.D(net10496),
.RN(net292),
.CK(clk),
.Q(net11054),
.QN(net11053)
);

DFFR_X2 merge9911(
.D(net10449),
.RN(net10252),
.CK(clk),
.Q(net11056),
.QN(net11055)
);

DFFS_X1 merge9912(
.D(net10357),
.SN(net9656),
.CK(clk),
.Q(net11058),
.QN(net11057)
);

DFFS_X2 merge9913(
.D(net10915),
.SN(net1554),
.CK(clk),
.Q(net11060),
.QN(net11059)
);

DFFR_X1 merge9914(
.D(net10139),
.RN(net10775),
.CK(clk),
.Q(net11062),
.QN(net11061)
);

AND2_X2 merge9915(
.A1(net6617),
.A2(net6516),
.ZN(net11063)
);

DFFR_X2 merge9916(
.D(net8489),
.RN(net9334),
.CK(clk),
.Q(net11065),
.QN(net11064)
);

DFFS_X1 merge9917(
.D(net6793),
.SN(net9464),
.CK(clk),
.Q(net11067),
.QN(net11066)
);

DFFS_X2 merge9918(
.D(net10379),
.SN(net10685),
.CK(clk),
.Q(net11069),
.QN(net11068)
);

DFFR_X1 merge9919(
.D(net4798),
.RN(net4774),
.CK(clk),
.Q(net11071),
.QN(net11070)
);

DFFR_X2 merge9920(
.D(net9954),
.RN(net10467),
.CK(clk),
.Q(net11073),
.QN(net11072)
);

DFFS_X1 merge9921(
.D(net1483),
.SN(net10703),
.CK(clk),
.Q(net11075),
.QN(net11074)
);

DFFS_X2 merge9922(
.D(net8974),
.SN(net9117),
.CK(clk),
.Q(net11077),
.QN(net11076)
);

DFFR_X1 merge9923(
.D(net10323),
.RN(net10007),
.CK(clk),
.Q(net11079),
.QN(net11078)
);

DFFR_X2 merge9924(
.D(net6492),
.RN(net9903),
.CK(clk),
.Q(net11081),
.QN(net11080)
);

DFFS_X1 merge9925(
.D(net8699),
.SN(net8637),
.CK(clk),
.Q(net11083),
.QN(net11082)
);

DFFS_X2 merge9926(
.D(net9720),
.SN(net10238),
.CK(clk),
.Q(net11085),
.QN(net11084)
);

DFFR_X1 merge9927(
.D(net10402),
.RN(net2592),
.CK(clk),
.Q(net11087),
.QN(net11086)
);

DFFR_X2 merge9928(
.D(net6720),
.RN(net6712),
.CK(clk),
.Q(net11089),
.QN(net11088)
);

DFFS_X1 merge9929(
.D(net7516),
.SN(net7419),
.CK(clk),
.Q(net11091),
.QN(net11090)
);

DFFS_X2 merge9930(
.D(net10658),
.SN(net10335),
.CK(clk),
.Q(net11093),
.QN(net11092)
);

DFFR_X1 merge9931(
.D(net9277),
.RN(net9243),
.CK(clk),
.Q(net11095),
.QN(net11094)
);

DFFR_X2 merge9932(
.D(net9092),
.RN(net8902),
.CK(clk),
.Q(net11097),
.QN(net11096)
);

DFFS_X1 merge9933(
.D(net6804),
.SN(net9638),
.CK(clk),
.Q(net11099),
.QN(net11098)
);

DFFS_X2 merge9934(
.D(net10729),
.SN(net6183),
.CK(clk),
.Q(net11101),
.QN(net11100)
);

DFFR_X1 merge9935(
.D(net5010),
.RN(net4055),
.CK(clk),
.Q(net11103),
.QN(net11102)
);

DFFR_X2 merge9936(
.D(net8140),
.RN(net8142),
.CK(clk),
.Q(net11105),
.QN(net11104)
);

DFFS_X1 merge9937(
.D(net10189),
.SN(net10202),
.CK(clk),
.Q(net11107),
.QN(net11106)
);

XOR2_X1 merge9938(
.A(net8022),
.B(net8941),
.Z(net11108)
);

DFFS_X2 merge9939(
.D(net2313),
.SN(net10262),
.CK(clk),
.Q(net11110),
.QN(net11109)
);

DFFR_X1 merge9940(
.D(net7735),
.RN(net8524),
.CK(clk),
.Q(net11112),
.QN(net11111)
);

DFFR_X2 merge9941(
.D(net814),
.RN(net2802),
.CK(clk),
.Q(net11114),
.QN(net11113)
);

DFFS_X1 merge9942(
.D(net1463),
.SN(net10162),
.CK(clk),
.Q(net11116),
.QN(net11115)
);

DFFS_X2 merge9943(
.D(net3639),
.SN(net10607),
.CK(clk),
.Q(net11118),
.QN(net11117)
);

DFFR_X1 merge9944(
.D(net6702),
.RN(net1626),
.CK(clk),
.Q(net11120),
.QN(net11119)
);

DFFR_X2 merge9945(
.D(net9296),
.RN(net7719),
.CK(clk),
.Q(net11122),
.QN(net11121)
);

DFFS_X1 merge9946(
.D(net9156),
.SN(net8381),
.CK(clk),
.Q(net11124),
.QN(net11123)
);

DFFS_X2 merge9947(
.D(net9572),
.SN(net9366),
.CK(clk),
.Q(net11126),
.QN(net11125)
);

DFFR_X1 merge9948(
.D(net9251),
.RN(net9054),
.CK(clk),
.Q(net11128),
.QN(net11127)
);

DFFR_X2 merge9949(
.D(net10263),
.RN(net10666),
.CK(clk),
.Q(net11130),
.QN(net11129)
);

DFFS_X1 merge9950(
.D(net10453),
.SN(net1238),
.CK(clk),
.Q(net11132),
.QN(net11131)
);

DFFS_X2 merge9951(
.D(net10064),
.SN(net9703),
.CK(clk),
.Q(net11134),
.QN(net11133)
);

DFFR_X1 merge9952(
.D(net9562),
.RN(net9489),
.CK(clk),
.Q(net11136),
.QN(net11135)
);

DFFR_X2 merge9953(
.D(net6759),
.RN(net6790),
.CK(clk),
.Q(net11137),
.QN(out5)
);

DFFS_X1 merge9954(
.D(net10709),
.SN(net10760),
.CK(clk),
.Q(net11139),
.QN(net11138)
);

DFFS_X2 merge9955(
.D(net8683),
.SN(net9367),
.CK(clk),
.Q(net11141),
.QN(net11140)
);

DFFR_X1 merge9956(
.D(net9557),
.RN(net9502),
.CK(clk),
.Q(net11143),
.QN(net11142)
);

DFFR_X2 merge9957(
.D(net7694),
.RN(net7668),
.CK(clk),
.Q(net11145),
.QN(net11144)
);

NOR2_X1 merge9958(
.A1(net9406),
.A2(net9323),
.ZN(net11146)
);

DFFS_X1 merge9959(
.D(net9291),
.SN(net8575),
.CK(clk),
.Q(net11148),
.QN(net11147)
);

DFFS_X2 merge9960(
.D(net3656),
.SN(net2665),
.CK(clk),
.Q(net11150),
.QN(net11149)
);

DFFR_X1 merge9961(
.D(net9986),
.RN(net10434),
.CK(clk),
.Q(net11152),
.QN(net11151)
);

DFFR_X2 merge9962(
.D(net8559),
.RN(net9459),
.CK(clk),
.Q(net11154),
.QN(net11153)
);

DFFS_X1 merge9963(
.D(net8712),
.SN(net7759),
.CK(clk),
.Q(net11156),
.QN(net11155)
);

DFFS_X2 merge9964(
.D(net1278),
.SN(net10023),
.CK(clk),
.Q(net11158),
.QN(net11157)
);

OR2_X2 merge9965(
.A1(net9143),
.A2(net9176),
.ZN(net11159)
);

DFFR_X1 merge9966(
.D(net8708),
.RN(net7749),
.CK(clk),
.Q(net11161),
.QN(net11160)
);

DFFR_X2 merge9967(
.D(net9153),
.RN(net8973),
.CK(clk),
.Q(net11163),
.QN(net11162)
);

DFFS_X1 merge9968(
.D(net7780),
.SN(net7717),
.CK(clk),
.Q(net11165),
.QN(net11164)
);

DFFS_X2 merge9969(
.D(net7786),
.SN(net8359),
.CK(clk),
.Q(net11167),
.QN(net11166)
);

DFFR_X1 merge9970(
.D(net445),
.RN(net3294),
.CK(clk),
.Q(net11169),
.QN(net11168)
);

DFFR_X2 merge9971(
.D(net10861),
.RN(net10181),
.CK(clk),
.Q(net11171),
.QN(net11170)
);

DFFS_X1 merge9972(
.D(net8971),
.SN(net9141),
.CK(clk),
.Q(net11173),
.QN(net11172)
);

DFFS_X2 merge9973(
.D(net10317),
.SN(net3653),
.CK(clk),
.Q(net11175),
.QN(net11174)
);

DFFR_X1 merge9974(
.D(net4116),
.RN(net10659),
.CK(clk),
.Q(net11177),
.QN(net11176)
);

DFFR_X2 merge9975(
.D(net9786),
.RN(net671),
.CK(clk),
.Q(net11179),
.QN(net11178)
);

DFFS_X1 merge9976(
.D(net8325),
.SN(net9437),
.CK(clk),
.Q(net11181),
.QN(net11180)
);

DFFS_X2 merge9977(
.D(net4188),
.SN(net9948),
.CK(clk),
.Q(net11183),
.QN(net11182)
);

DFFR_X1 merge9978(
.D(net6181),
.RN(net10241),
.CK(clk),
.Q(net11185),
.QN(net11184)
);

DFFR_X2 merge9979(
.D(net8525),
.RN(net8554),
.CK(clk),
.Q(net11187),
.QN(net11186)
);

DFFS_X1 merge9980(
.D(net10825),
.SN(net10460),
.CK(clk),
.Q(net11189),
.QN(net11188)
);

DFFS_X2 merge9981(
.D(net10612),
.SN(net6180),
.CK(clk),
.Q(net11191),
.QN(net11190)
);

DFFR_X1 merge9982(
.D(net10234),
.RN(net10356),
.CK(clk),
.Q(net11193),
.QN(net11192)
);

DFFR_X2 merge9983(
.D(net9450),
.RN(net9274),
.CK(clk),
.Q(net11195),
.QN(net11194)
);

DFFS_X1 merge9984(
.D(net9252),
.SN(net9233),
.CK(clk),
.Q(net11197),
.QN(net11196)
);

DFFS_X2 merge9985(
.D(net7785),
.SN(net7748),
.CK(clk),
.Q(net11199),
.QN(net11198)
);

DFFR_X1 merge9986(
.D(net10867),
.RN(net3229),
.CK(clk),
.Q(net11201),
.QN(net11200)
);

DFFR_X2 merge9987(
.D(net9401),
.RN(net8570),
.CK(clk),
.Q(net11203),
.QN(net11202)
);

DFFS_X1 merge9988(
.D(net7626),
.SN(net7660),
.CK(clk),
.Q(net11205),
.QN(net11204)
);

DFFS_X2 merge9989(
.D(net9768),
.SN(net10284),
.CK(clk),
.Q(net11207),
.QN(net11206)
);

DFFR_X1 merge9990(
.D(net9352),
.RN(net10611),
.CK(clk),
.Q(net11209),
.QN(net11208)
);

DFFR_X2 merge9991(
.D(net8629),
.RN(net9547),
.CK(clk),
.Q(net11211),
.QN(net11210)
);

DFFS_X1 merge9992(
.D(net10540),
.SN(net2680),
.CK(clk),
.Q(net11213),
.QN(net11212)
);

DFFS_X2 merge9993(
.D(net9724),
.SN(net10190),
.CK(clk),
.Q(net11215),
.QN(net11214)
);

DFFR_X1 merge9994(
.D(net10624),
.RN(net10437),
.CK(clk),
.Q(net11217),
.QN(net11216)
);

DFFR_X2 merge9995(
.D(net9585),
.RN(net9550),
.CK(clk),
.Q(net11219),
.QN(net11218)
);

DFFS_X1 merge9996(
.D(net10305),
.SN(net4242),
.CK(clk),
.Q(net11221),
.QN(net11220)
);

DFFS_X2 merge9997(
.D(net10082),
.SN(net10199),
.CK(clk),
.Q(net11223),
.QN(net11222)
);

NOR2_X4 merge9998(
.A1(net9482),
.A2(net8515),
.ZN(net11224)
);

DFFR_X1 merge9999(
.D(net7663),
.RN(net7757),
.CK(clk),
.Q(net11226),
.QN(net11225)
);

DFFR_X2 merge10000(
.D(net10092),
.RN(net9901),
.CK(clk),
.Q(net11228),
.QN(net11227)
);

DFFS_X1 merge10001(
.D(net7773),
.SN(net9544),
.CK(clk),
.Q(net11230),
.QN(net11229)
);

DFFS_X2 merge10002(
.D(net4653),
.SN(net5628),
.CK(clk),
.Q(net11232),
.QN(net11231)
);

DFFR_X1 merge10003(
.D(net10508),
.RN(net10220),
.CK(clk),
.Q(net11234),
.QN(net11233)
);

DFFR_X2 merge10004(
.D(net8614),
.RN(net9556),
.CK(clk),
.Q(net11236),
.QN(net11235)
);

DFFS_X1 merge10005(
.D(net2154),
.SN(net238),
.CK(clk),
.Q(net11238),
.QN(net11237)
);

DFFS_X2 merge10006(
.D(net8500),
.SN(net10800),
.CK(clk),
.Q(net11240),
.QN(net11239)
);

DFFR_X1 merge10007(
.D(net10575),
.RN(net7777),
.CK(clk),
.Q(net11242),
.QN(net11241)
);

DFFR_X2 merge10008(
.D(net8932),
.RN(net8025),
.CK(clk),
.Q(net11244),
.QN(net11243)
);

DFFS_X1 merge10009(
.D(net3331),
.SN(net1371),
.CK(clk),
.Q(net11246),
.QN(net11245)
);

DFFS_X2 merge10010(
.D(net7009),
.SN(net8029),
.CK(clk),
.Q(net11248),
.QN(net11247)
);

DFFR_X1 merge10011(
.D(net9753),
.RN(net9712),
.CK(clk),
.Q(net11250),
.QN(net11249)
);

DFFR_X2 merge10012(
.D(net10420),
.RN(net10908),
.CK(clk),
.Q(net11252),
.QN(net11251)
);

DFFS_X1 merge10013(
.D(net9483),
.SN(net8564),
.CK(clk),
.Q(net11254),
.QN(net11253)
);

DFFS_X2 merge10014(
.D(net9765),
.SN(net10296),
.CK(clk),
.Q(net11256),
.QN(net11255)
);

DFFR_X1 merge10015(
.D(net9421),
.RN(net9467),
.CK(clk),
.Q(net11258),
.QN(net11257)
);

DFFR_X2 merge10016(
.D(net9560),
.RN(net8684),
.CK(clk),
.Q(net11260),
.QN(net11259)
);

DFFS_X1 merge10017(
.D(net8244),
.SN(net10819),
.CK(clk),
.Q(net11262),
.QN(net11261)
);

DFFS_X2 merge10018(
.D(net7767),
.SN(net9577),
.CK(clk),
.Q(net11264),
.QN(net11263)
);

DFFR_X1 merge10019(
.D(net8633),
.RN(net9871),
.CK(clk),
.Q(net11266),
.QN(net11265)
);

DFFR_X2 merge10020(
.D(net3686),
.RN(net10567),
.CK(clk),
.Q(net11268),
.QN(net11267)
);

DFFS_X1 merge10021(
.D(net10352),
.SN(net10672),
.CK(clk),
.Q(net11270),
.QN(net11269)
);

DFFS_X2 merge10022(
.D(net10348),
.SN(net2149),
.CK(clk),
.Q(net11272),
.QN(net11271)
);

DFFR_X1 merge10023(
.D(net8697),
.RN(net8703),
.CK(clk),
.Q(out23),
.QN(net11273)
);

DFFR_X2 merge10024(
.D(net1387),
.RN(net3364),
.CK(clk),
.Q(net11275),
.QN(net11274)
);

DFFS_X1 merge10025(
.D(net10121),
.SN(net10221),
.CK(clk),
.Q(net11277),
.QN(net11276)
);

DFFS_X2 merge10026(
.D(net10834),
.SN(net10872),
.CK(clk),
.Q(net11279),
.QN(net11278)
);

NOR2_X2 merge10027(
.A1(net9510),
.A2(net9535),
.ZN(net11280)
);

DFFR_X1 merge10028(
.D(net8731),
.RN(net8705),
.CK(clk),
.Q(net11282),
.QN(net11281)
);

DFFR_X2 merge10029(
.D(net10222),
.RN(net6191),
.CK(clk),
.Q(net11284),
.QN(net11283)
);

DFFS_X1 merge10030(
.D(net10015),
.SN(net10479),
.CK(clk),
.Q(net11286),
.QN(net11285)
);

DFFS_X2 merge10031(
.D(net7771),
.SN(net7774),
.CK(clk),
.Q(net11288),
.QN(net11287)
);

DFFR_X1 merge10032(
.D(net10526),
.RN(net10505),
.CK(clk),
.Q(net11290),
.QN(net11289)
);

DFFR_X2 merge10033(
.D(net9607),
.RN(net9534),
.CK(clk),
.Q(net11292),
.QN(net11291)
);

DFFS_X1 merge10034(
.D(net8735),
.SN(net8709),
.CK(clk),
.Q(net11294),
.QN(net11293)
);

DFFS_X2 merge10035(
.D(net10135),
.SN(net10736),
.CK(clk),
.Q(net11296),
.QN(net11295)
);

XOR2_X2 merge10036(
.A(net9599),
.B(net8716),
.Z(net11297)
);

DFFR_X1 merge10037(
.D(net10523),
.RN(net10198),
.CK(clk),
.Q(net11299),
.QN(net11298)
);

DFFR_X2 merge10038(
.D(net10367),
.RN(net10011),
.CK(clk),
.Q(net11301),
.QN(net11300)
);

DFFS_X1 merge10039(
.D(net10655),
.SN(net10291),
.CK(clk),
.Q(net11303),
.QN(net11302)
);

DFFS_X2 merge10040(
.D(net8704),
.Q(net11304),
.CK(clk),
.QN(out2)
);

DFFR_X1 merge10041(
.D(net10961),
.RN(net7250),
.CK(clk),
.Q(net11306),
.QN(net11305)
);

DFFR_X2 merge10042(
.D(net1538),
.RN(net10848),
.CK(clk),
.Q(net11308),
.QN(net11307)
);

DFFS_X1 merge10043(
.D(net10922),
.SN(net9695),
.CK(clk),
.Q(net11310),
.QN(net11309)
);

DFFS_X2 merge10044(
.D(net10675),
.SN(net4375),
.CK(clk),
.Q(net11312),
.QN(net11311)
);

DFFR_X1 merge10045(
.D(net10336),
.RN(net10907),
.CK(clk),
.Q(net11314),
.QN(net11313)
);

DFFR_X2 merge10046(
.D(net9600),
.RN(net9617),
.CK(clk),
.Q(net11316),
.QN(net11315)
);

DFFS_X1 merge10047(
.D(net10142),
.SN(net10478),
.CK(clk),
.Q(net11318),
.QN(net11317)
);

DFFS_X2 merge10048(
.D(net8714),
.SN(net8715),
.CK(clk),
.Q(out10),
.QN(net11319)
);

DFFR_X1 merge10049(
.D(net2221),
.RN(net10454),
.CK(clk),
.Q(net11321),
.QN(net11320)
);

DFFR_X2 merge10050(
.D(net4292),
.RN(net10776),
.CK(clk),
.Q(net11323),
.QN(net11322)
);

DFFS_X1 merge10051(
.D(net9632),
.SN(net9633),
.CK(clk),
.Q(net11325),
.QN(net11324)
);

DFFS_X2 merge10052(
.D(net10223),
.SN(net5158),
.CK(clk),
.Q(net11327),
.QN(net11326)
);

DFFR_X1 merge10053(
.D(net9639),
.RN(net8717),
.CK(clk),
.Q(net11328),
.QN(out7)
);

DFFR_X2 merge10054(
.D(net11159),
.RN(net9707),
.CK(clk),
.Q(net11330),
.QN(net11329)
);

DFFS_X1 merge10055(
.D(net10035),
.SN(net9892),
.CK(clk),
.Q(net11332),
.QN(net11331)
);

DFFS_X2 merge10056(
.D(net10077),
.SN(net10165),
.CK(clk),
.Q(net11334),
.QN(net11333)
);

DFFR_X1 merge10057(
.D(net9827),
.RN(net10733),
.CK(clk),
.Q(net11336),
.QN(net11335)
);

DFFR_X2 merge10058(
.D(net10237),
.RN(net2147),
.CK(clk),
.Q(net11338),
.QN(net11337)
);

DFFS_X1 merge10059(
.D(net9997),
.SN(net3776),
.CK(clk),
.Q(net11340),
.QN(net11339)
);

DFFS_X2 merge10060(
.D(net11224),
.SN(net6684),
.CK(clk),
.Q(net11342),
.QN(net11341)
);

DFFR_X1 merge10061(
.D(net10706),
.RN(net10812),
.CK(clk),
.Q(net11344),
.QN(net11343)
);

DFFR_X2 merge10062(
.D(net10255),
.RN(net10822),
.CK(clk),
.Q(net11346),
.QN(net11345)
);

DFFS_X1 merge10063(
.D(net10850),
.SN(net1476),
.CK(clk),
.Q(net11348),
.QN(net11347)
);

DFFS_X2 merge10064(
.D(net10080),
.SN(net2748),
.CK(clk),
.Q(net11350),
.QN(net11349)
);

DFFR_X1 merge10065(
.D(net10928),
.RN(net10113),
.CK(clk),
.Q(net11352),
.QN(net11351)
);

DFFR_X2 merge10066(
.D(net10493),
.RN(net6489),
.CK(clk),
.Q(net11354),
.QN(net11353)
);

DFFS_X1 merge10067(
.D(net10702),
.SN(net10621),
.CK(clk),
.Q(net11356),
.QN(net11355)
);

DFFS_X2 merge10068(
.D(net9704),
.SN(net2355),
.CK(clk),
.Q(net11358),
.QN(net11357)
);

DFFR_X1 merge10069(
.D(net10048),
.RN(net10782),
.CK(clk),
.Q(net11360),
.QN(net11359)
);

DFFR_X2 merge10070(
.D(net304),
.RN(net10781),
.CK(clk),
.Q(net11362),
.QN(net11361)
);

DFFS_X1 merge10071(
.D(net9893),
.SN(net9746),
.CK(clk),
.Q(net11364),
.QN(net11363)
);

DFFS_X2 merge10072(
.D(net7298),
.SN(net10459),
.CK(clk),
.Q(net11366),
.QN(net11365)
);

DFFR_X1 merge10073(
.D(net474),
.RN(net10170),
.CK(clk),
.Q(net11368),
.QN(net11367)
);

DFFR_X2 merge10074(
.D(net10586),
.RN(net10051),
.CK(clk),
.Q(net11370),
.QN(net11369)
);

DFFS_X1 merge10075(
.D(net4330),
.SN(net2162),
.CK(clk),
.Q(net11372),
.QN(net11371)
);

DFFS_X2 merge10076(
.D(net9822),
.SN(net10792),
.CK(clk),
.Q(net11374),
.QN(net11373)
);

DFFR_X1 merge10077(
.D(net10925),
.RN(net10034),
.CK(clk),
.Q(net11376),
.QN(net11375)
);

DFFR_X2 merge10078(
.D(net9866),
.RN(net10894),
.CK(clk),
.Q(net11378),
.QN(net11377)
);

DFFS_X1 merge10079(
.D(net10442),
.SN(net10485),
.CK(clk),
.Q(net11380),
.QN(net11379)
);

DFFS_X2 merge10080(
.D(net9959),
.SN(net9987),
.CK(clk),
.Q(net11382),
.QN(net11381)
);

DFFR_X1 merge10081(
.D(net10081),
.RN(net9988),
.CK(clk),
.Q(net11384),
.QN(net11383)
);

DFFR_X2 merge10082(
.D(net5283),
.RN(net10205),
.CK(clk),
.Q(net11386),
.QN(net11385)
);

DFFS_X1 merge10083(
.D(net10210),
.SN(net11297),
.CK(clk),
.Q(net11388),
.QN(net11387)
);

DFFS_X2 merge10084(
.D(net10065),
.SN(net7574),
.CK(clk),
.Q(net11390),
.QN(net11389)
);

DFFR_X1 merge10085(
.D(net10295),
.RN(net10895),
.CK(clk),
.Q(net11392),
.QN(net11391)
);

DFFR_X2 merge10086(
.D(net11012),
.RN(net10219),
.CK(clk),
.Q(net11394),
.QN(net11393)
);

DFFS_X1 merge10087(
.D(net11036),
.SN(net9433),
.CK(clk),
.Q(net11396),
.QN(net11395)
);

DFFS_X2 merge10088(
.D(net10755),
.SN(net10608),
.CK(clk),
.Q(net11398),
.QN(net11397)
);

DFFR_X1 merge10089(
.D(net6529),
.RN(net6261),
.CK(clk),
.Q(net11400),
.QN(net11399)
);

DFFR_X2 merge10090(
.D(net10292),
.RN(net10063),
.CK(clk),
.Q(net11402),
.QN(net11401)
);

DFFS_X1 merge10091(
.D(net9995),
.SN(net9671),
.CK(clk),
.Q(net11404),
.QN(net11403)
);

DFFS_X2 merge10092(
.D(net9748),
.SN(net4320),
.CK(clk),
.Q(net11406),
.QN(net11405)
);

DFFR_X1 merge10093(
.D(net9937),
.RN(net1501),
.CK(clk),
.Q(net11408),
.QN(net11407)
);

DFFR_X2 merge10094(
.D(net10342),
.RN(net11029),
.CK(clk),
.Q(net11410),
.QN(net11409)
);

DFFS_X1 merge10095(
.D(net10619),
.SN(net10000),
.CK(clk),
.Q(net11412),
.QN(net11411)
);

DFFS_X2 merge10096(
.D(net10732),
.SN(net10620),
.CK(clk),
.Q(net11414),
.QN(net11413)
);

DFFR_X1 merge10097(
.D(net10413),
.RN(net7428),
.CK(clk),
.Q(net11416),
.QN(net11415)
);

DFFR_X2 merge10098(
.D(net10101),
.RN(net10218),
.CK(clk),
.Q(net11418),
.QN(net11417)
);

DFFS_X1 merge10099(
.D(net10268),
.SN(net10273),
.CK(clk),
.Q(net11420),
.QN(net11419)
);

DFFS_X2 merge10100(
.D(net4125),
.SN(net10906),
.CK(clk),
.Q(net11422),
.QN(net11421)
);

DFFR_X1 merge10101(
.D(net10211),
.RN(net10784),
.CK(clk),
.Q(net11424),
.QN(net11423)
);

DFFR_X2 merge10102(
.D(net11146),
.RN(net9477),
.CK(clk),
.Q(net11426),
.QN(net11425)
);

DFFS_X1 merge10103(
.D(net9666),
.SN(net10916),
.CK(clk),
.Q(net11428),
.QN(net11427)
);

DFFS_X2 merge10104(
.D(net10072),
.SN(net10650),
.CK(clk),
.Q(net11430),
.QN(net11429)
);

DFFR_X1 merge10105(
.D(net10527),
.RN(net8357),
.CK(clk),
.Q(net11432),
.QN(net11431)
);

DFFR_X2 merge10106(
.D(net8317),
.RN(net10841),
.CK(clk),
.Q(net11434),
.QN(net11433)
);

DFFS_X1 merge10107(
.D(net6184),
.SN(net10579),
.CK(clk),
.Q(net11436),
.QN(net11435)
);

DFFS_X2 merge10108(
.D(net10847),
.SN(net10864),
.CK(clk),
.Q(net11438),
.QN(net11437)
);

DFFR_X1 merge10109(
.D(net10917),
.RN(net10799),
.CK(clk),
.Q(net11440),
.QN(net11439)
);

DFFR_X2 merge10110(
.D(net10364),
.RN(net10151),
.CK(clk),
.Q(net11442),
.QN(net11441)
);

DFFS_X1 merge10111(
.D(net10646),
.SN(net10543),
.CK(clk),
.Q(net11444),
.QN(net11443)
);

DFFS_X2 merge10112(
.D(net9698),
.SN(net9735),
.CK(clk),
.Q(net11446),
.QN(net11445)
);

DFFR_X1 merge10113(
.D(net10934),
.RN(net10783),
.CK(clk),
.Q(net11448),
.QN(net11447)
);

DFFR_X2 merge10114(
.D(net10568),
.RN(net9911),
.CK(clk),
.Q(net11450),
.QN(net11449)
);

DFFS_X1 merge10115(
.D(net10801),
.SN(net11063),
.CK(clk),
.Q(net11452),
.QN(net11451)
);

DFFS_X2 merge10116(
.D(net8323),
.SN(net9777),
.CK(clk),
.Q(net11454),
.QN(net11453)
);

DFFR_X1 merge10117(
.D(net9728),
.RN(net9810),
.CK(clk),
.Q(net11456),
.QN(net11455)
);

DFFR_X2 merge10118(
.D(net10071),
.RN(net10560),
.CK(clk),
.Q(net11458),
.QN(net11457)
);

DFFS_X1 merge10119(
.D(net10425),
.SN(net10343),
.CK(clk),
.Q(net11460),
.QN(net11459)
);

DFFS_X2 merge10120(
.D(net9784),
.SN(net7148),
.CK(clk),
.Q(net11462),
.QN(net11461)
);

DFFR_X1 merge10121(
.D(net10003),
.RN(net11280),
.CK(clk),
.Q(net11464),
.QN(net11463)
);

DFFR_X2 merge10122(
.D(net3754),
.RN(net10197),
.CK(clk),
.Q(net11466),
.QN(net11465)
);

DFFS_X1 merge10123(
.D(net2264),
.SN(net10933),
.CK(clk),
.Q(net11468),
.QN(net11467)
);

DFFS_X2 merge10124(
.D(net10997),
.SN(net10353),
.CK(clk),
.Q(out0),
.QN(net11469)
);

DFFR_X1 merge10125(
.D(net9996),
.RN(net2711),
.CK(clk),
.Q(net11471),
.QN(net11470)
);

DFFR_X2 merge10126(
.D(net10482),
.RN(net10231),
.CK(clk),
.Q(net11473),
.QN(net11472)
);

DFFS_X1 merge10127(
.D(net9787),
.SN(net10645),
.CK(clk),
.Q(net11475),
.QN(net11474)
);

DFFS_X2 merge10128(
.D(net10403),
.SN(net10688),
.CK(clk),
.Q(net11477),
.QN(net11476)
);

DFFR_X1 merge10129(
.D(net10070),
.RN(net10842),
.CK(clk),
.Q(net11479),
.QN(net11478)
);

DFFR_X2 merge10130(
.D(net10754),
.RN(net7415),
.CK(clk),
.Q(net11481),
.QN(net11480)
);

DFFS_X1 merge10131(
.D(net5280),
.SN(net10138),
.CK(clk),
.Q(net11483),
.QN(net11482)
);

DFFS_X2 merge10132(
.D(net4663),
.SN(net10182),
.CK(clk),
.Q(net11485),
.QN(net11484)
);

DFFR_X1 merge10133(
.D(net9687),
.RN(net10085),
.CK(clk),
.Q(net11487),
.QN(net11486)
);

DFFR_X2 merge10134(
.D(net10887),
.RN(net11108),
.CK(clk),
.Q(net11489),
.QN(net11488)
);

DFFS_X1 merge10135(
.D(net6619),
.SN(net10351),
.CK(clk),
.Q(net11491),
.QN(net11490)
);

DFF_X1 s10136(
.D(net228),
.CK(clk),
.Q(net11493),
.QN(net11492)
);

DFF_X2 s10137(
.D(net569),
.CK(clk),
.Q(net11495),
.QN(net11494)
);

DFF_X1 s10138(
.D(net590),
.CK(clk),
.Q(net11497),
.QN(net11496)
);

DFF_X2 s10139(
.D(net591),
.CK(clk),
.Q(net11499),
.QN(net11498)
);

DFF_X1 s10140(
.D(net1052),
.CK(clk),
.Q(net11501),
.QN(net11500)
);

DFF_X2 s10141(
.D(net1116),
.CK(clk),
.Q(net11503),
.QN(net11502)
);

DFF_X1 s10142(
.D(net1208),
.CK(clk),
.Q(net11505),
.QN(net11504)
);

DFF_X2 s10143(
.D(net1531),
.CK(clk),
.Q(net11507),
.QN(net11506)
);

DFF_X1 s10144(
.D(net1882),
.CK(clk),
.Q(net11509),
.QN(net11508)
);

DFF_X2 s10145(
.D(net2008),
.CK(clk),
.Q(net11511),
.QN(net11510)
);

DFF_X1 s10146(
.D(net2329),
.CK(clk),
.Q(net11513),
.QN(net11512)
);

DFF_X2 s10147(
.D(net2444),
.CK(clk),
.Q(net11515),
.QN(net11514)
);

DFF_X1 s10148(
.D(net2449),
.CK(clk),
.Q(net11517),
.QN(net11516)
);

DFF_X2 s10149(
.D(net2454),
.CK(clk),
.Q(net11519),
.QN(net11518)
);

DFF_X1 s10150(
.D(net2901),
.CK(clk),
.Q(net11521),
.QN(net11520)
);

DFF_X2 s10151(
.D(net3510),
.CK(clk),
.Q(net11523),
.QN(net11522)
);

DFF_X1 s10152(
.D(net3673),
.CK(clk),
.Q(net11525),
.QN(net11524)
);

DFF_X2 s10153(
.D(net3946),
.CK(clk),
.Q(net11527),
.QN(net11526)
);

DFF_X1 s10154(
.D(net4134),
.CK(clk),
.Q(net11529),
.QN(net11528)
);

DFF_X2 s10155(
.D(net4170),
.CK(clk),
.Q(net11531),
.QN(net11530)
);

DFF_X1 s10156(
.D(net4323),
.CK(clk),
.Q(net11533),
.QN(net11532)
);

DFF_X2 s10157(
.D(net4816),
.CK(clk),
.Q(net11535),
.QN(net11534)
);

DFF_X1 s10158(
.D(net4829),
.CK(clk),
.Q(net11537),
.QN(net11536)
);

DFF_X2 s10159(
.D(net4938),
.CK(clk),
.Q(net11539),
.QN(net11538)
);

DFF_X1 s10160(
.D(net5035),
.CK(clk),
.Q(net11541),
.QN(net11540)
);

DFF_X2 s10161(
.D(net5270),
.CK(clk),
.Q(net11543),
.QN(net11542)
);

DFF_X1 s10162(
.D(net5747),
.CK(clk),
.Q(net11545),
.QN(net11544)
);

DFF_X2 s10163(
.D(net5831),
.CK(clk),
.Q(net11547),
.QN(net11546)
);

DFF_X1 s10164(
.D(net5920),
.CK(clk),
.Q(net11549),
.QN(net11548)
);

DFF_X2 s10165(
.D(net6019),
.CK(clk),
.Q(net11551),
.QN(net11550)
);

DFF_X1 s10166(
.D(net6623),
.CK(clk),
.Q(net11553),
.QN(net11552)
);

DFF_X2 s10167(
.D(net6889),
.CK(clk),
.Q(net11555),
.QN(net11554)
);

DFF_X1 s10168(
.D(net6895),
.CK(clk),
.Q(net11557),
.QN(net11556)
);

DFF_X2 s10169(
.D(net7245),
.CK(clk),
.Q(net11559),
.QN(net11558)
);

DFF_X1 s10170(
.D(net7424),
.CK(clk),
.Q(net11561),
.QN(net11560)
);

DFF_X2 s10171(
.D(net7605),
.CK(clk),
.Q(net11563),
.QN(net11562)
);

DFF_X1 s10172(
.D(net7858),
.CK(clk),
.Q(net11565),
.QN(net11564)
);

DFF_X2 s10173(
.D(net7879),
.CK(clk),
.Q(net11567),
.QN(net11566)
);

DFF_X1 s10174(
.D(net8147),
.CK(clk),
.Q(net11569),
.QN(net11568)
);

DFF_X2 s10175(
.D(net8227),
.CK(clk),
.Q(net11571),
.QN(net11570)
);

DFF_X1 s10176(
.D(net8376),
.CK(clk),
.Q(net11573),
.QN(net11572)
);

DFF_X2 s10177(
.D(net8387),
.CK(clk),
.Q(net11575),
.QN(net11574)
);

DFF_X1 s10178(
.D(net8496),
.CK(clk),
.Q(net11577),
.QN(net11576)
);

DFF_X2 s10179(
.D(net8829),
.CK(clk),
.Q(net11579),
.QN(net11578)
);

DFF_X1 s10180(
.D(net9180),
.CK(clk),
.Q(net11581),
.QN(net11580)
);

DFF_X2 s10181(
.D(net9315),
.CK(clk),
.Q(net11583),
.QN(net11582)
);

DFF_X1 s10182(
.D(net9472),
.CK(clk),
.Q(net11585),
.QN(net11584)
);

DFF_X2 s10183(
.D(net9555),
.CK(clk),
.Q(net11587),
.QN(net11586)
);

DFF_X1 s10184(
.D(net9725),
.CK(clk),
.Q(net11589),
.QN(net11588)
);


endmodule
