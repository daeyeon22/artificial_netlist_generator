module test_circuit (
	input in0,
	input in1,
	input in2,
	input in3,
	input in4,
	input in5,
	input in6,
	input in7,
	input in8,
	input in9,
	input in10,
	input in11,
	input in12,
	input in13,
	input in14,
	input in15,
	input in16,
	input in17,
	input in18,
	input in19,
	input in20,
	input in21,
	input in22,
	input in23,
	input in24,
	input in25,
	input clk,
	input rst,
	output out0,
	output out1,
	output out2,
	output out3,
	output out4,
	output out5,
	output out6,
	output out7,
	output out8,
	output out9,
	output out10,
	output out11,
	output out12,
	output out13,
	output out14,
	output out15,
	output out16,
	output out17,
	output out18,
	output out19,
	output out20,
	output out21,
	output out22,
	output out23,
	output out24,
	output out25
);


wire net11237;
wire net11236;
wire net11235;
wire net11234;
wire net11233;
wire net11231;
wire net11230;
wire net11228;
wire net11227;
wire net11221;
wire net11220;
wire net11216;
wire net11215;
wire net11212;
wire net11210;
wire net11209;
wire net11208;
wire net11206;
wire net11205;
wire net11204;
wire net11203;
wire net11202;
wire net11201;
wire net11198;
wire net11197;
wire net11195;
wire net11194;
wire net11192;
wire net11191;
wire net11190;
wire net11188;
wire net11186;
wire net11185;
wire net11177;
wire net11174;
wire net11170;
wire net11168;
wire net11165;
wire net11163;
wire net11161;
wire net11160;
wire net11159;
wire net11158;
wire net11157;
wire net11156;
wire net11151;
wire net11150;
wire net11148;
wire net11144;
wire net11142;
wire net11137;
wire net11133;
wire net11132;
wire net11127;
wire net11126;
wire net11124;
wire net11123;
wire out0;
wire net11120;
wire net11116;
wire net11115;
wire net11112;
wire net11108;
wire net11107;
wire net11106;
wire net11102;
wire net11100;
wire net11099;
wire net11091;
wire net11090;
wire net11088;
wire net11086;
wire net11083;
wire net11082;
wire net11080;
wire net11078;
wire net11077;
wire net11073;
wire net11072;
wire net11069;
wire net11067;
wire net11065;
wire net11064;
wire net11063;
wire net11059;
wire net11058;
wire net11057;
wire net11056;
wire net11054;
wire net11062;
wire net11051;
wire net11049;
wire net11048;
wire net11046;
wire net11044;
wire net11042;
wire net11041;
wire net11040;
wire net11039;
wire net11036;
wire net11035;
wire net11034;
wire net11027;
wire net11026;
wire net11025;
wire net11023;
wire net11021;
wire net11016;
wire out7;
wire net11015;
wire out10;
wire net11010;
wire net11008;
wire net11007;
wire net11003;
wire net11189;
wire net11001;
wire out2;
wire net10997;
wire net10996;
wire net10992;
wire net10988;
wire net10981;
wire net10980;
wire net10979;
wire net10976;
wire net10968;
wire net10967;
wire net10965;
wire net10962;
wire net10961;
wire net10959;
wire net10957;
wire net10955;
wire net10954;
wire net10953;
wire net10945;
wire net10944;
wire net10943;
wire net10942;
wire net10938;
wire net10937;
wire net10936;
wire net10935;
wire net10934;
wire net10933;
wire net10932;
wire net10930;
wire net10928;
wire net10927;
wire net10924;
wire net10922;
wire net10921;
wire net10913;
wire net10912;
wire net10910;
wire net10908;
wire net10906;
wire net10905;
wire net10903;
wire net10902;
wire net10900;
wire net10899;
wire net10898;
wire net10896;
wire net10894;
wire net10893;
wire net10889;
wire net10887;
wire net10886;
wire net10885;
wire net10883;
wire net10874;
wire net10873;
wire out5;
wire net10871;
wire net10869;
wire net10866;
wire net10865;
wire net10864;
wire net10862;
wire net10861;
wire net10859;
wire net10858;
wire net10857;
wire net10855;
wire net10850;
wire net10848;
wire net10847;
wire net10843;
wire net10842;
wire net10841;
wire net10840;
wire net10839;
wire net10836;
wire net10835;
wire net10831;
wire net10830;
wire net10828;
wire net10827;
wire net10825;
wire net10824;
wire net10823;
wire net10821;
wire net10837;
wire net10820;
wire net10818;
wire net10817;
wire net10816;
wire net10815;
wire net10814;
wire net10812;
wire net10811;
wire net10808;
wire net10806;
wire net10804;
wire net10802;
wire net10801;
wire net10800;
wire net10798;
wire net10797;
wire net10796;
wire net10795;
wire net10793;
wire net10791;
wire net10789;
wire net10787;
wire net10786;
wire net10785;
wire net10782;
wire net10780;
wire net10779;
wire net10771;
wire net10767;
wire net10764;
wire net10762;
wire net10759;
wire net10758;
wire net10757;
wire net10755;
wire net10750;
wire net10749;
wire net10748;
wire net10747;
wire net10746;
wire net10745;
wire net10743;
wire net10742;
wire net10735;
wire net10734;
wire net10733;
wire net10730;
wire net10729;
wire net10727;
wire net10725;
wire net10724;
wire net10719;
wire net10718;
wire net10717;
wire net10715;
wire net10711;
wire net10710;
wire net10709;
wire net10705;
wire net10704;
wire net10703;
wire net10700;
wire net10699;
wire net10693;
wire net10692;
wire net10691;
wire net10690;
wire net10689;
wire net10687;
wire net10685;
wire net10683;
wire net10681;
wire net10679;
wire net10677;
wire net10675;
wire net10673;
wire net10672;
wire net10670;
wire net10669;
wire net10667;
wire net10666;
wire net10665;
wire net10664;
wire net10662;
wire net10658;
wire net10656;
wire net10652;
wire net10650;
wire net10648;
wire net10647;
wire net10646;
wire net10645;
wire net10640;
wire net10638;
wire net10637;
wire net10634;
wire net10631;
wire net10625;
wire net10623;
wire net10622;
wire net10621;
wire net10620;
wire net10619;
wire net10613;
wire net10610;
wire net10609;
wire net10607;
wire net10604;
wire net10602;
wire net10601;
wire net10600;
wire net10597;
wire net10595;
wire net10594;
wire net10592;
wire net10591;
wire net10585;
wire net10583;
wire net10580;
wire net10579;
wire net10578;
wire net10576;
wire net10575;
wire net10574;
wire net10572;
wire net10571;
wire net10567;
wire net10565;
wire net10564;
wire net10563;
wire net10736;
wire net10561;
wire net10559;
wire net10558;
wire net10553;
wire net11152;
wire net10552;
wire net10551;
wire net10549;
wire net10548;
wire net10546;
wire net10545;
wire net10544;
wire net10538;
wire net10535;
wire net10533;
wire net10532;
wire net10526;
wire net10524;
wire net10523;
wire net10522;
wire net10520;
wire net10519;
wire net10518;
wire net10517;
wire net10515;
wire net10511;
wire net10510;
wire net10509;
wire net10503;
wire net10498;
wire net10497;
wire net10494;
wire net10493;
wire net10492;
wire net10490;
wire net10487;
wire net10485;
wire net10482;
wire net10778;
wire net10479;
wire net10475;
wire net10474;
wire net10473;
wire net10472;
wire net10505;
wire net10469;
wire net10468;
wire net10461;
wire net10456;
wire net10455;
wire net10453;
wire net10451;
wire net10448;
wire net10446;
wire net10445;
wire net10440;
wire net10439;
wire net10438;
wire net10436;
wire net10435;
wire net10433;
wire net10431;
wire net10430;
wire net10428;
wire net10425;
wire net10424;
wire net10423;
wire net10422;
wire net10419;
wire net10416;
wire net10414;
wire net10413;
wire net10412;
wire net10411;
wire net10409;
wire net10408;
wire net10404;
wire net10403;
wire net10401;
wire net10400;
wire net10398;
wire net10395;
wire net10394;
wire net10385;
wire net10384;
wire net10382;
wire net10381;
wire net10379;
wire net10378;
wire net10377;
wire net10376;
wire net10375;
wire net10969;
wire net10368;
wire net10367;
wire net10364;
wire net10363;
wire net10358;
wire net10353;
wire net10348;
wire net10343;
wire net10341;
wire net10340;
wire net10339;
wire net10911;
wire net10335;
wire net10334;
wire net10333;
wire net10332;
wire net10330;
wire net10329;
wire net10328;
wire net10326;
wire net10323;
wire net10322;
wire net10321;
wire net10320;
wire net10318;
wire net10317;
wire net10311;
wire net10310;
wire net10307;
wire net10306;
wire net10305;
wire net10303;
wire net10301;
wire net10300;
wire net10299;
wire net10297;
wire net10295;
wire net10293;
wire net10292;
wire net10291;
wire net10290;
wire net10288;
wire net10286;
wire net10285;
wire net10283;
wire net11172;
wire net10280;
wire net10277;
wire net10276;
wire net10275;
wire net10274;
wire net10272;
wire net10271;
wire net10269;
wire net10268;
wire net10267;
wire net10266;
wire net10265;
wire net10260;
wire net10259;
wire net10257;
wire net11061;
wire net10256;
wire net10255;
wire net10253;
wire net10252;
wire net10249;
wire net11131;
wire net10248;
wire net10244;
wire net10242;
wire net10240;
wire net10239;
wire net10287;
wire net10238;
wire net10236;
wire net10235;
wire net10234;
wire net10232;
wire net10231;
wire net10229;
wire net10226;
wire net10225;
wire net10224;
wire net10222;
wire net10221;
wire net10219;
wire net10218;
wire net10216;
wire net10215;
wire net10214;
wire net10211;
wire net10210;
wire net10209;
wire net10204;
wire net10202;
wire net10201;
wire net10193;
wire net10190;
wire net10186;
wire net10185;
wire net10184;
wire net10183;
wire net10182;
wire net10181;
wire net10180;
wire net10179;
wire net10175;
wire net10174;
wire net10173;
wire net10169;
wire net10168;
wire net10167;
wire net10784;
wire net10164;
wire net10160;
wire net10155;
wire net10154;
wire net10152;
wire net10151;
wire net10149;
wire net10146;
wire net10145;
wire net10228;
wire net10144;
wire net10141;
wire net10138;
wire net10136;
wire net10135;
wire net10132;
wire net10131;
wire net10129;
wire net10127;
wire net10126;
wire net10125;
wire net10124;
wire net10118;
wire net10117;
wire net10116;
wire net10114;
wire net10109;
wire net10108;
wire net10107;
wire net10105;
wire net10104;
wire net10102;
wire net10099;
wire net10098;
wire net10096;
wire net10095;
wire net10092;
wire net10091;
wire net10089;
wire net10088;
wire net10582;
wire net10087;
wire net10086;
wire net10085;
wire net10082;
wire net10080;
wire net10075;
wire net10073;
wire net10324;
wire net10072;
wire net10071;
wire net10070;
wire net10067;
wire net10066;
wire net10064;
wire net10061;
wire net10053;
wire net10051;
wire net10048;
wire net10047;
wire net10046;
wire net10044;
wire net10043;
wire net10042;
wire net10041;
wire net10039;
wire net10033;
wire net10031;
wire net10030;
wire net10028;
wire net10027;
wire net10024;
wire net10022;
wire net10020;
wire net10017;
wire net10016;
wire net10015;
wire net10011;
wire net10009;
wire net10153;
wire net10008;
wire net10005;
wire net10001;
wire net10000;
wire net9997;
wire net9992;
wire net9991;
wire net9988;
wire net9987;
wire net9985;
wire net9983;
wire net9982;
wire net9980;
wire net9979;
wire net9978;
wire net9976;
wire net9975;
wire net9974;
wire net9973;
wire net9970;
wire net9968;
wire net10465;
wire net9966;
wire net9961;
wire net9960;
wire net9959;
wire net9958;
wire net9957;
wire net9953;
wire net10566;
wire net9951;
wire net9948;
wire net11146;
wire net9947;
wire net10845;
wire net9938;
wire net9937;
wire net9935;
wire net9934;
wire net9931;
wire net9927;
wire net9925;
wire net9924;
wire net9923;
wire net9922;
wire net9918;
wire net9917;
wire net9916;
wire net9912;
wire net9911;
wire net9995;
wire net9909;
wire net9908;
wire net10270;
wire net9907;
wire net9906;
wire net9905;
wire net9901;
wire net9900;
wire net9899;
wire net9898;
wire net9896;
wire net10464;
wire net9894;
wire net9893;
wire net9891;
wire net9887;
wire net9884;
wire net9883;
wire net9881;
wire net9879;
wire net9878;
wire net11141;
wire net9877;
wire net9876;
wire net9871;
wire net9870;
wire net10337;
wire net9869;
wire net9868;
wire net9865;
wire net9863;
wire net9862;
wire net10060;
wire net9861;
wire net9860;
wire net9859;
wire net9858;
wire net9857;
wire net10246;
wire net9856;
wire net9855;
wire net9852;
wire net9850;
wire net9847;
wire net9845;
wire net9843;
wire net10189;
wire net9932;
wire net9841;
wire net9839;
wire net9836;
wire net9833;
wire net9831;
wire net10489;
wire net9830;
wire net9826;
wire net9825;
wire net9823;
wire net9822;
wire net9821;
wire net9820;
wire net9816;
wire net9812;
wire net9809;
wire net9807;
wire net9805;
wire net10313;
wire net9803;
wire net10856;
wire net9802;
wire net9801;
wire net9798;
wire net9797;
wire net9796;
wire net9795;
wire net9791;
wire net9790;
wire net9789;
wire net10296;
wire net9788;
wire net9786;
wire net9785;
wire net9783;
wire net9781;
wire net9780;
wire net9778;
wire net9774;
wire net9773;
wire net9772;
wire net9769;
wire net9768;
wire net9766;
wire net10629;
wire net9765;
wire net9764;
wire net9761;
wire net9760;
wire net9759;
wire net9758;
wire net9757;
wire net9756;
wire net9755;
wire net9751;
wire net9750;
wire net9749;
wire net9748;
wire net9747;
wire net9746;
wire net9743;
wire net11176;
wire net9742;
wire net9741;
wire net9739;
wire net9738;
wire net9737;
wire net9735;
wire net9777;
wire net9734;
wire net9732;
wire net9731;
wire net9729;
wire net9727;
wire net9726;
wire net9724;
wire net9723;
wire net9721;
wire net9720;
wire net9715;
wire net9711;
wire net9709;
wire net9708;
wire net9704;
wire net9703;
wire net9700;
wire net9699;
wire net9696;
wire net9695;
wire net9694;
wire net9693;
wire net9692;
wire net9691;
wire net9690;
wire net9689;
wire net9688;
wire net9685;
wire net9683;
wire net9682;
wire net9680;
wire net9678;
wire net9677;
wire net9675;
wire net9673;
wire net9672;
wire net9671;
wire net10369;
wire net9668;
wire net9667;
wire net9665;
wire net10187;
wire net9663;
wire net9661;
wire net9660;
wire net9659;
wire net9657;
wire net9653;
wire net9651;
wire net9679;
wire net9650;
wire net9649;
wire net9648;
wire net9647;
wire net9645;
wire net9641;
wire net9640;
wire net9638;
wire net10282;
wire net9634;
wire net9631;
wire net9629;
wire net9628;
wire net9625;
wire net9623;
wire net9622;
wire net9621;
wire net9753;
wire net9618;
wire net10018;
wire net9617;
wire net9616;
wire net9613;
wire net9612;
wire net9610;
wire net9607;
wire net9606;
wire net9604;
wire net10162;
wire net9603;
wire net9602;
wire net9601;
wire net9600;
wire net9598;
wire net9597;
wire net9596;
wire net9594;
wire net9592;
wire net9591;
wire net9589;
wire net9588;
wire net9587;
wire net9585;
wire net10651;
wire net9583;
wire net9581;
wire net11011;
wire net10279;
wire net9580;
wire net9579;
wire net9578;
wire net9576;
wire net9575;
wire net9574;
wire net10142;
wire net9573;
wire net9571;
wire net9570;
wire net9568;
wire net9565;
wire net9561;
wire net9555;
wire net9548;
wire net9547;
wire net9545;
wire net9544;
wire net9538;
wire net9537;
wire net9535;
wire net9534;
wire net9533;
wire net9529;
wire net9528;
wire net9525;
wire net9524;
wire net9519;
wire net9518;
wire net9516;
wire net9515;
wire net9514;
wire net9513;
wire net9512;
wire net9511;
wire net9508;
wire net9507;
wire net10918;
wire net9506;
wire net10999;
wire net9505;
wire net9504;
wire net9503;
wire net9502;
wire net9500;
wire net9499;
wire net9496;
wire net9492;
wire net9484;
wire net10365;
wire net9483;
wire net9479;
wire net9474;
wire net9473;
wire net9470;
wire net9469;
wire net9467;
wire net9464;
wire net9462;
wire net10254;
wire net9459;
wire net9457;
wire net9455;
wire net11125;
wire net9454;
wire net9452;
wire net9449;
wire net10829;
wire net9448;
wire net11187;
wire net9444;
wire net9443;
wire net9439;
wire net9438;
wire net9437;
wire net9436;
wire net9434;
wire net10853;
wire net9432;
wire net9431;
wire net9430;
wire net9429;
wire net9427;
wire net9424;
wire net9423;
wire net9422;
wire net9421;
wire net9419;
wire net9418;
wire net9416;
wire net9415;
wire net9412;
wire net9411;
wire net9632;
wire net9407;
wire net9406;
wire net9405;
wire net9404;
wire net9399;
wire net9398;
wire net9394;
wire net10587;
wire net9393;
wire net9392;
wire net9390;
wire net9389;
wire net9387;
wire net9386;
wire net9385;
wire net9384;
wire net9383;
wire net9381;
wire net9378;
wire net9377;
wire net9376;
wire net9375;
wire net9373;
wire net9369;
wire net9364;
wire net9363;
wire net9362;
wire net9361;
wire net9360;
wire net9358;
wire net9357;
wire net9356;
wire net9352;
wire net9351;
wire net9350;
wire net10396;
wire net9349;
wire net10611;
wire net9347;
wire net9346;
wire net9344;
wire net9343;
wire net9342;
wire net9341;
wire net9338;
wire net9337;
wire net9336;
wire net9333;
wire net9332;
wire net9331;
wire net9330;
wire net9326;
wire net9325;
wire net9324;
wire net9323;
wire net9320;
wire net9316;
wire net10161;
wire net9315;
wire net9314;
wire net9313;
wire net9311;
wire net10712;
wire net9310;
wire net9309;
wire net9306;
wire net9305;
wire net9304;
wire net10525;
wire net9303;
wire net10094;
wire net9300;
wire net9299;
wire net9298;
wire net9294;
wire net9293;
wire net10663;
wire net9291;
wire net9290;
wire net9295;
wire net9289;
wire net9288;
wire net9283;
wire net9282;
wire net9281;
wire net9280;
wire net9278;
wire net9276;
wire net10956;
wire net9275;
wire net9269;
wire net9268;
wire net9266;
wire net9265;
wire net9263;
wire net9261;
wire net9256;
wire net9253;
wire net9252;
wire net9251;
wire net9250;
wire net9248;
wire net9244;
wire net9240;
wire net9239;
wire net9237;
wire net9236;
wire net9234;
wire net9231;
wire net9228;
wire net9227;
wire net9226;
wire net9339;
wire net9224;
wire net9222;
wire net9221;
wire net9220;
wire net9215;
wire net9213;
wire net9212;
wire net9211;
wire net9210;
wire net9209;
wire net9208;
wire net9207;
wire net9205;
wire net10176;
wire net9204;
wire net9200;
wire net9199;
wire net9197;
wire net9195;
wire net9194;
wire net9193;
wire net9190;
wire net9188;
wire net9185;
wire net9183;
wire net10506;
wire net9182;
wire net9536;
wire net9181;
wire net9180;
wire net9178;
wire net9176;
wire net9175;
wire net9171;
wire net9167;
wire net9166;
wire net9165;
wire net9164;
wire net9161;
wire net9160;
wire net9159;
wire net9158;
wire net9258;
wire net9157;
wire net9156;
wire net11103;
wire net9154;
wire net9153;
wire net9152;
wire net9151;
wire net9147;
wire net9146;
wire net9145;
wire net9144;
wire net10447;
wire net9142;
wire net9141;
wire net9139;
wire net9136;
wire net9133;
wire net9132;
wire net9131;
wire net9130;
wire net9967;
wire net9126;
wire net9116;
wire net9174;
wire net9114;
wire net9112;
wire net9108;
wire net9107;
wire net9106;
wire net9105;
wire net9103;
wire net9100;
wire net9099;
wire net9095;
wire net9091;
wire net9090;
wire net9089;
wire net9088;
wire net9087;
wire net9674;
wire net9086;
wire net9084;
wire net9083;
wire net9081;
wire net9080;
wire net9076;
wire net9075;
wire net9488;
wire net9074;
wire net9073;
wire net9071;
wire net9069;
wire net9068;
wire net9063;
wire net9061;
wire net9059;
wire net9058;
wire net9057;
wire net9056;
wire net9710;
wire net9054;
wire net9053;
wire net9052;
wire net9051;
wire net9050;
wire net9046;
wire net9989;
wire net9045;
wire net9040;
wire net9039;
wire net9038;
wire net9035;
wire net9032;
wire net9029;
wire net9027;
wire net9026;
wire net9020;
wire net9019;
wire net9018;
wire net9016;
wire net9015;
wire net10504;
wire net9014;
wire net9013;
wire net9011;
wire net9010;
wire net9007;
wire net9005;
wire net9463;
wire net9004;
wire net9003;
wire net9002;
wire net9001;
wire net9000;
wire net8998;
wire net10359;
wire net8997;
wire net8996;
wire net8995;
wire net8993;
wire net8992;
wire net8991;
wire net8989;
wire net8986;
wire net8984;
wire net8983;
wire net8982;
wire net8980;
wire net9475;
wire net8978;
wire net8976;
wire net8975;
wire net8974;
wire net8973;
wire net8972;
wire net10543;
wire net8970;
wire net8969;
wire net8968;
wire net8966;
wire net8965;
wire net8961;
wire net8959;
wire net8958;
wire net8956;
wire net8954;
wire net8953;
wire net8946;
wire net8945;
wire net8941;
wire net8940;
wire net8939;
wire net8937;
wire net10312;
wire net8934;
wire net8927;
wire net9630;
wire net8924;
wire net8921;
wire net9155;
wire net8920;
wire net8919;
wire net8917;
wire net8915;
wire net8913;
wire net8905;
wire net8903;
wire net8902;
wire net8901;
wire net8900;
wire net8899;
wire net8897;
wire net8895;
wire net8893;
wire net11038;
wire net8890;
wire net8889;
wire net8887;
wire net8885;
wire net8884;
wire net8882;
wire net9238;
wire net8880;
wire net8877;
wire net8876;
wire net8875;
wire net8873;
wire net8871;
wire net8870;
wire net8869;
wire net8868;
wire net8867;
wire net8865;
wire net8863;
wire net8862;
wire net8861;
wire net10958;
wire net8860;
wire net8858;
wire net10593;
wire net8857;
wire net8856;
wire net8864;
wire net8855;
wire net8854;
wire net8853;
wire net8852;
wire net8851;
wire net8850;
wire net8849;
wire net8845;
wire net8844;
wire net8838;
wire net8837;
wire net8836;
wire net9055;
wire net8831;
wire net9806;
wire net8827;
wire net8826;
wire net8822;
wire net8821;
wire net8820;
wire net8819;
wire net8816;
wire net10442;
wire net10241;
wire net8814;
wire net8812;
wire net8811;
wire net8810;
wire net8809;
wire net8808;
wire net8806;
wire net8803;
wire net11092;
wire net8802;
wire net8799;
wire net8798;
wire net8796;
wire net8795;
wire net10388;
wire net9043;
wire net8791;
wire net8787;
wire net8786;
wire net8785;
wire net8784;
wire net11085;
wire net8782;
wire net8780;
wire net8779;
wire net8777;
wire net10081;
wire net8776;
wire net8769;
wire net8768;
wire net8766;
wire net8764;
wire net8763;
wire net9752;
wire net8762;
wire net8761;
wire net8760;
wire net8758;
wire net8753;
wire net8751;
wire net8750;
wire net8749;
wire net8747;
wire net8746;
wire net8745;
wire net8744;
wire net8741;
wire net8740;
wire net8739;
wire net8738;
wire net8737;
wire net8736;
wire net8735;
wire net8733;
wire net8732;
wire net8731;
wire net8728;
wire net10140;
wire net8727;
wire net8726;
wire net10530;
wire net8725;
wire net10178;
wire net8724;
wire net8723;
wire net9828;
wire net8722;
wire net8721;
wire net8720;
wire net8719;
wire net8717;
wire net8715;
wire net8714;
wire net8713;
wire net8712;
wire net8805;
wire net8710;
wire net8708;
wire net8707;
wire net8705;
wire net8704;
wire net8702;
wire net8701;
wire net8699;
wire net8696;
wire net10963;
wire net8695;
wire net8693;
wire net8692;
wire net8691;
wire net8689;
wire net8918;
wire net8688;
wire net8686;
wire net8683;
wire net8682;
wire net9490;
wire net8681;
wire net8680;
wire net8678;
wire net8677;
wire net8675;
wire net8673;
wire net8672;
wire net8671;
wire net8669;
wire net8668;
wire net8667;
wire net8666;
wire net8665;
wire net8661;
wire net8660;
wire net10716;
wire net10084;
wire net8658;
wire net8653;
wire net8652;
wire net8651;
wire net8648;
wire net8646;
wire net9170;
wire net8644;
wire net8643;
wire net8642;
wire out12;
wire net8641;
wire net8639;
wire net10529;
wire net8638;
wire net8718;
wire net8637;
wire net8636;
wire out14;
wire net8635;
wire net8634;
wire net9192;
wire net8633;
wire net8632;
wire out22;
wire net8631;
wire net11028;
wire net8628;
wire net10660;
wire net8626;
wire net8625;
wire net10741;
wire net8624;
wire net8623;
wire net8621;
wire net8619;
wire net9784;
wire out18;
wire net8615;
wire net11183;
wire net8874;
wire net8613;
wire net8611;
wire out11;
wire net8981;
wire net8607;
wire net8606;
wire net8605;
wire net8600;
wire net8598;
wire net8597;
wire out6;
wire net8589;
wire net8588;
wire net10882;
wire net8587;
wire net10148;
wire net8585;
wire net8584;
wire net8971;
wire net8580;
wire net8579;
wire net8577;
wire net9875;
wire net8576;
wire net8574;
wire net8572;
wire net8571;
wire net8570;
wire net8569;
wire net8568;
wire net11098;
wire net8567;
wire net8564;
wire net8560;
wire net8558;
wire net8556;
wire net8555;
wire net8554;
wire net8553;
wire net8552;
wire net9892;
wire net8551;
wire net11145;
wire net8911;
wire net8549;
wire net8547;
wire net8546;
wire net11229;
wire net8545;
wire net8544;
wire net8929;
wire net8541;
wire net8539;
wire net8538;
wire net8534;
wire net8530;
wire net9371;
wire net8529;
wire net8528;
wire net8527;
wire net10012;
wire net8526;
wire net8525;
wire net8524;
wire net8815;
wire net8521;
wire net10437;
wire net8520;
wire net8519;
wire net8518;
wire net8513;
wire net8512;
wire net10345;
wire net9225;
wire net8510;
wire net8509;
wire net8507;
wire net8498;
wire net8497;
wire net9840;
wire net8495;
wire net8493;
wire net8492;
wire net11093;
wire net8489;
wire net8488;
wire net8486;
wire net8480;
wire net8479;
wire net10247;
wire net8478;
wire net8477;
wire net8475;
wire net11214;
wire net8474;
wire net8471;
wire net8469;
wire net8468;
wire net8466;
wire net8462;
wire net8460;
wire net11012;
wire net8459;
wire net8458;
wire net8456;
wire net8523;
wire net8455;
wire net8454;
wire net8453;
wire net8452;
wire net8450;
wire net8449;
wire net8444;
wire net8442;
wire net8438;
wire net8437;
wire net8434;
wire net8433;
wire net8432;
wire net8429;
wire net8842;
wire net8428;
wire net10586;
wire net8427;
wire net8426;
wire net8425;
wire net8423;
wire net8421;
wire net8418;
wire net8417;
wire net8414;
wire net8413;
wire net8412;
wire net8411;
wire net8410;
wire net8409;
wire net8781;
wire net8408;
wire net8407;
wire net8406;
wire net8405;
wire net8404;
wire net8400;
wire net8397;
wire net8396;
wire net8395;
wire net8394;
wire net8391;
wire net8390;
wire net8389;
wire net8388;
wire net8387;
wire net8382;
wire net8381;
wire net8378;
wire net9955;
wire net8377;
wire net8374;
wire net8372;
wire net8371;
wire net8369;
wire net8368;
wire net8367;
wire net8366;
wire net8365;
wire net8363;
wire net8362;
wire net8360;
wire net8358;
wire net8355;
wire net8353;
wire net10237;
wire net8350;
wire net8348;
wire net9522;
wire net8347;
wire net8685;
wire net8345;
wire net9374;
wire net8344;
wire net8343;
wire net8342;
wire net8341;
wire net8339;
wire net9111;
wire net8337;
wire net8335;
wire net10596;
wire net8332;
wire net9654;
wire net8331;
wire net8330;
wire net8329;
wire net8328;
wire net8326;
wire net8323;
wire net8322;
wire net8321;
wire out20;
wire net8319;
wire net8318;
wire net8317;
wire net8316;
wire net8314;
wire net9030;
wire net8312;
wire net8306;
wire net8304;
wire net8301;
wire net8300;
wire net8297;
wire net8296;
wire net8295;
wire net8292;
wire net8288;
wire net8286;
wire net8284;
wire net8283;
wire net8281;
wire net8280;
wire net8279;
wire net8276;
wire net8273;
wire net8272;
wire net8271;
wire net10230;
wire net8269;
wire net8266;
wire net8265;
wire net8264;
wire net8263;
wire net8261;
wire net9233;
wire net8260;
wire net8357;
wire net8257;
wire net8254;
wire net8253;
wire net8252;
wire net8249;
wire net10036;
wire net8247;
wire net8245;
wire net8244;
wire net8242;
wire net8241;
wire net8240;
wire net8239;
wire net8238;
wire net8236;
wire net8235;
wire net8234;
wire net8232;
wire net8231;
wire net10177;
wire net8227;
wire net8226;
wire net8225;
wire net8223;
wire net8222;
wire net8220;
wire net8219;
wire net8218;
wire net8217;
wire net8216;
wire net8213;
wire net8212;
wire net8210;
wire net9279;
wire net8209;
wire net8208;
wire net10386;
wire net8207;
wire net8206;
wire net8205;
wire net8203;
wire net8202;
wire net11128;
wire net8201;
wire net8199;
wire net8198;
wire net8754;
wire net8197;
wire net8196;
wire net8195;
wire net11169;
wire net8193;
wire net8191;
wire net8190;
wire net8188;
wire net8187;
wire net8186;
wire net10916;
wire net8185;
wire net8183;
wire net8179;
wire net8178;
wire net8175;
wire net9187;
wire net8172;
wire net8823;
wire net8168;
wire net8166;
wire net8165;
wire net8164;
wire net8161;
wire net8159;
wire net8158;
wire net9605;
wire net8157;
wire net8156;
wire net8155;
wire net8153;
wire net8516;
wire net8152;
wire net10338;
wire net8150;
wire net8149;
wire net8148;
wire net9713;
wire net8146;
wire net8145;
wire net8144;
wire net8143;
wire net8142;
wire net8140;
wire net8139;
wire net8138;
wire net9493;
wire net8136;
wire net8129;
wire net8128;
wire net8127;
wire net8125;
wire net8124;
wire net8123;
wire net8119;
wire net8118;
wire net8117;
wire net8114;
wire net10194;
wire net8113;
wire net8112;
wire net8448;
wire net8110;
wire net10618;
wire net8109;
wire net8106;
wire net8105;
wire net8101;
wire net8100;
wire net8097;
wire net8096;
wire net8095;
wire net8093;
wire net10486;
wire net8092;
wire net9366;
wire net8087;
wire net8084;
wire net9286;
wire net8083;
wire net8082;
wire net10844;
wire net9885;
wire net8081;
wire net10200;
wire net8080;
wire net8077;
wire net8076;
wire net9701;
wire net8075;
wire net8074;
wire net8073;
wire net8069;
wire net8068;
wire net8066;
wire net8063;
wire net8062;
wire net8060;
wire net8058;
wire net8057;
wire net8055;
wire net8051;
wire net8050;
wire net8049;
wire net8048;
wire net8047;
wire net8046;
wire net8044;
wire net8043;
wire net8042;
wire net8040;
wire net8039;
wire net8035;
wire net8034;
wire net8032;
wire net10415;
wire net8788;
wire net8030;
wire net8029;
wire net8028;
wire net8027;
wire net8026;
wire net9963;
wire net8025;
wire net8024;
wire net8023;
wire net8021;
wire net8018;
wire net8017;
wire net8016;
wire net8015;
wire net8012;
wire net8011;
wire net8009;
wire net8007;
wire net11094;
wire net10355;
wire net8006;
wire net8005;
wire net11110;
wire net8004;
wire net8003;
wire net8002;
wire net8001;
wire net7999;
wire net7997;
wire net7996;
wire net10123;
wire net8496;
wire net7994;
wire net7993;
wire net7991;
wire net10387;
wire net7990;
wire net7989;
wire net7988;
wire net7986;
wire net7985;
wire net7983;
wire net7980;
wire net7977;
wire net7974;
wire net7973;
wire net7970;
wire net7960;
wire net7958;
wire net7954;
wire net7953;
wire net7950;
wire net7949;
wire net9322;
wire net7948;
wire net11050;
wire net7944;
wire net8305;
wire net7943;
wire net7939;
wire net7937;
wire net7935;
wire net8354;
wire net7934;
wire net7933;
wire net7932;
wire net7930;
wire net7929;
wire net7928;
wire net7926;
wire net7925;
wire net7924;
wire net7923;
wire net7921;
wire net7920;
wire net7919;
wire net7917;
wire net7915;
wire net7914;
wire net7913;
wire net11217;
wire net9287;
wire net7912;
wire net7911;
wire net7910;
wire net9666;
wire net7909;
wire net10630;
wire net7908;
wire net7906;
wire net7905;
wire net11014;
wire net7902;
wire net7892;
wire net7891;
wire net7890;
wire net7889;
wire net7887;
wire net7884;
wire net7881;
wire net7879;
wire net8938;
wire net7878;
wire net7876;
wire net7874;
wire net7873;
wire net7871;
wire net9191;
wire net7870;
wire net7869;
wire out17;
wire net7865;
wire net7864;
wire net7863;
wire net7862;
wire net7861;
wire net8684;
wire net7860;
wire net7857;
wire net8091;
wire net7855;
wire net7852;
wire net7850;
wire net7849;
wire net7848;
wire net7847;
wire net7845;
wire net7843;
wire net7841;
wire net7840;
wire net7836;
wire net7833;
wire net7832;
wire net7824;
wire net7823;
wire net7822;
wire net7816;
wire net7814;
wire net7813;
wire net7812;
wire net7811;
wire net7810;
wire net7809;
wire net7806;
wire net7803;
wire net7802;
wire net7797;
wire net7796;
wire net7795;
wire net7794;
wire net10418;
wire net7791;
wire net7790;
wire net7789;
wire net7787;
wire net7786;
wire net7785;
wire net7781;
wire net7779;
wire net7777;
wire net7776;
wire net7772;
wire net7771;
wire net7770;
wire net7769;
wire net7767;
wire net7765;
wire net9633;
wire net7763;
wire net7762;
wire net7761;
wire net8916;
wire net7760;
wire net7759;
wire net9644;
wire net7758;
wire net7756;
wire net7755;
wire net7754;
wire net7753;
wire net10120;
wire net7752;
wire net7984;
wire net7751;
wire net7749;
wire net7748;
wire net7746;
wire net7745;
wire net7743;
wire net7742;
wire net7740;
wire net7737;
wire net7733;
wire net7732;
wire net7731;
wire net10458;
wire net7730;
wire net10951;
wire net7729;
wire net7726;
wire net7725;
wire net7724;
wire net7723;
wire net7721;
wire net7719;
wire net7715;
wire net7714;
wire net7712;
wire net7711;
wire net7710;
wire net7708;
wire net7707;
wire net7706;
wire net7704;
wire net7703;
wire net7699;
wire net9851;
wire net7696;
wire net7694;
wire net7693;
wire net7691;
wire net7688;
wire net7687;
wire net7686;
wire net7679;
wire net7678;
wire net7784;
wire net7675;
wire net7674;
wire net7671;
wire net7670;
wire net7669;
wire net7668;
wire net7666;
wire net7665;
wire net7663;
wire net7662;
wire net7660;
wire net7659;
wire net10470;
wire net7656;
wire net7655;
wire net7654;
wire net7653;
wire net7652;
wire net7651;
wire net8988;
wire net7648;
wire net9260;
wire net7647;
wire net7645;
wire net7644;
wire net7643;
wire net7642;
wire net10929;
wire net8550;
wire net7641;
wire net7640;
wire net7636;
wire net7634;
wire net7633;
wire net7632;
wire net7631;
wire net7629;
wire net10480;
wire net7628;
wire net7627;
wire net7626;
wire net7625;
wire net7624;
wire net10143;
wire net7621;
wire net7619;
wire net7617;
wire net7615;
wire net7614;
wire net9025;
wire net7609;
wire out19;
wire net7607;
wire net7605;
wire net8752;
wire net7603;
wire net7601;
wire net11109;
wire net7600;
wire net7598;
wire net7595;
wire net7594;
wire net7593;
wire net7592;
wire net7591;
wire net9771;
wire net7590;
wire net8385;
wire net7588;
wire net7587;
wire net7586;
wire net7585;
wire net7584;
wire net7582;
wire net7581;
wire net7579;
wire net9335;
wire net7577;
wire net7572;
wire net9113;
wire net7571;
wire net7570;
wire net7569;
wire net7568;
wire net7566;
wire net7565;
wire net7564;
wire net7562;
wire net7561;
wire net7560;
wire net7559;
wire net8131;
wire net7558;
wire net11181;
wire net7556;
wire net9705;
wire net7554;
wire net7553;
wire net7549;
wire net9717;
wire net7547;
wire net10639;
wire net7546;
wire net7545;
wire net7543;
wire net7541;
wire net7540;
wire net7539;
wire net9586;
wire net7538;
wire net7537;
wire net7956;
wire net7536;
wire net7535;
wire net7533;
wire net7531;
wire net10720;
wire net7530;
wire net7529;
wire net7527;
wire net9611;
wire net7526;
wire net7525;
wire net7523;
wire net7522;
wire net7521;
wire net7520;
wire net7519;
wire net9669;
wire net7518;
wire net7517;
wire net7516;
wire net7514;
wire net7510;
wire net7509;
wire net8102;
wire net7508;
wire net7507;
wire net7505;
wire net7503;
wire net7502;
wire net7501;
wire net7500;
wire net10147;
wire net8979;
wire net7499;
wire net7498;
wire net7657;
wire net7497;
wire net7493;
wire net11045;
wire net10488;
wire net7489;
wire net10678;
wire net7488;
wire net3712;
wire net10603;
wire net3650;
wire net5066;
wire net5427;
wire net3699;
wire net4859;
wire net3697;
wire net7427;
wire net10644;
wire net3692;
wire net3687;
wire net11095;
wire net3684;
wire net4757;
wire net3678;
wire net3673;
wire net2661;
wire net3672;
wire net4673;
wire net8338;
wire net5036;
wire net1050;
wire net3670;
wire net9022;
wire net3669;
wire net6666;
wire net3662;
wire net3657;
wire net10570;
wire net4219;
wire net8888;
wire net5980;
wire net7194;
wire net6390;
wire net3648;
wire net3641;
wire net1859;
wire net3637;
wire net4378;
wire net3635;
wire net8103;
wire net3622;
wire net324;
wire net3615;
wire net3609;
wire net649;
wire net6312;
wire net9079;
wire net3601;
wire net3597;
wire net3596;
wire net3590;
wire net3695;
wire net7859;
wire net4122;
wire net3588;
wire net3390;
wire net2119;
wire net3584;
wire net60;
wire net3582;
wire net3578;
wire net3575;
wire net3574;
wire net3570;
wire net4709;
wire net3567;
wire net3559;
wire net2665;
wire net3557;
wire net3556;
wire net1002;
wire net4495;
wire net3129;
wire net377;
wire net3548;
wire net8832;
wire net3660;
wire net5247;
wire net3546;
wire net2380;
wire net3545;
wire net9569;
wire net8104;
wire net3544;
wire net8593;
wire net6638;
wire net3543;
wire net7268;
wire net9933;
wire net3539;
wire net3538;
wire net3536;
wire net4159;
wire net8346;
wire net3535;
wire net3529;
wire net2047;
wire net3525;
wire net7410;
wire net3523;
wire net3521;
wire net10833;
wire net5119;
wire net3517;
wire net7271;
wire net7931;
wire net3512;
wire net3175;
wire net9138;
wire net3511;
wire net3509;
wire net4564;
wire net11053;
wire net6676;
wire net3508;
wire net3507;
wire net9740;
wire net3502;
wire net3500;
wire net3494;
wire net919;
wire net7196;
wire net8470;
wire net3493;
wire net5719;
wire net3491;
wire net3489;
wire net10007;
wire net329;
wire net3488;
wire net8908;
wire net7311;
wire net3487;
wire net3532;
wire net3486;
wire net3485;
wire net3484;
wire net3480;
wire net4321;
wire net3478;
wire net3476;
wire net10826;
wire net2043;
wire net9033;
wire net3473;
wire net571;
wire net3469;
wire net3466;
wire net3455;
wire net3451;
wire net8303;
wire net3260;
wire net3649;
wire net3449;
wire net5042;
wire net8022;
wire net5709;
wire net3444;
wire net2461;
wire net3442;
wire net3440;
wire net3439;
wire net144;
wire net3519;
wire net872;
wire net5099;
wire net6791;
wire net3426;
wire net8603;
wire net2003;
wire net6715;
wire net3427;
wire net3542;
wire net9328;
wire net3423;
wire net3419;
wire net4987;
wire net3688;
wire net171;
wire net4354;
wire net3638;
wire net11079;
wire net8536;
wire net3411;
wire net2884;
wire net3410;
wire net3408;
wire net1343;
wire net10555;
wire net10350;
wire net6850;
wire net3547;
wire net3406;
wire net8189;
wire net135;
wire net3401;
wire net7616;
wire net3396;
wire net3210;
wire net3394;
wire net3387;
wire net5745;
wire net3384;
wire net3382;
wire net3380;
wire net3377;
wire net7513;
wire net6701;
wire net9292;
wire net3376;
wire net3366;
wire net3370;
wire net7428;
wire net3369;
wire net10854;
wire net9124;
wire net3367;
wire net3363;
wire net1951;
wire net7285;
wire net9115;
wire net3360;
wire net621;
wire net5422;
wire net3354;
wire net1870;
wire net3350;
wire net3345;
wire net5930;
wire net9854;
wire net4533;
wire net3634;
wire net3341;
wire net7183;
wire net3339;
wire net5845;
wire net3336;
wire net10914;
wire net354;
wire net3330;
wire net3327;
wire net10636;
wire net1054;
wire net10212;
wire net6551;
wire net3326;
wire net3325;
wire net9148;
wire net3323;
wire net5533;
wire net3318;
wire net7804;
wire net4881;
wire net3316;
wire net1321;
wire net3314;
wire net1702;
wire net3302;
wire net3294;
wire net9273;
wire net3288;
wire net3286;
wire net3284;
wire net581;
wire net7415;
wire net3921;
wire net3280;
wire net2894;
wire net3589;
wire net3691;
wire net5590;
wire net8038;
wire net3278;
wire net2687;
wire net10738;
wire net3277;
wire net3275;
wire net4097;
wire net9541;
wire net3658;
wire net10499;
wire net3257;
wire net2284;
wire net7220;
wire net11213;
wire net3252;
wire net3246;
wire net3234;
wire net3240;
wire net3239;
wire net5808;
wire net7269;
wire in24;
wire net4645;
wire net7416;
wire net3235;
wire net6464;
wire net3232;
wire net3230;
wire net532;
wire net5925;
wire net3228;
wire net3149;
wire net3227;
wire net5044;
wire net3225;
wire net11068;
wire net3224;
wire net3438;
wire net10769;
wire net7695;
wire net1451;
wire net8793;
wire net3219;
wire net3218;
wire net5214;
wire net5183;
wire net3211;
wire net3352;
wire net8336;
wire net5697;
wire net7075;
wire net3207;
wire net2852;
wire net9919;
wire net7286;
wire net11196;
wire net3198;
wire net3193;
wire net11118;
wire net6500;
wire net3191;
wire net10635;
wire net3186;
wire net3184;
wire net4949;
wire net3180;
wire net7267;
wire net3647;
wire net3177;
wire net3173;
wire net7727;
wire net3169;
wire net9972;
wire net9810;
wire net1060;
wire net3165;
wire net3498;
wire net3157;
wire net8833;
wire net3375;
wire net8472;
wire net147;
wire net3145;
wire net3143;
wire net3141;
wire net3140;
wire net3137;
wire net3134;
wire net3130;
wire net3126;
wire net8771;
wire net2091;
wire net533;
wire net10615;
wire net5789;
wire net6923;
wire net7018;
wire net3160;
wire net6275;
wire net3121;
wire net1918;
wire net10756;
wire net3112;
wire net126;
wire net3111;
wire net8663;
wire net7511;
wire net3067;
wire net2981;
wire net8839;
wire net3110;
wire net5123;
wire net3109;
wire net3102;
wire net224;
wire net836;
wire net5999;
wire net5375;
wire net3097;
wire net9684;
wire net3321;
wire net3096;
wire net8542;
wire net8464;
wire net749;
wire net2783;
wire net7998;
wire net3459;
wire net5815;
wire net7006;
wire net3088;
wire net7242;
wire net10895;
wire net7567;
wire net3125;
wire net3526;
wire net7927;
wire net5683;
wire net3085;
wire net1175;
wire net2560;
wire net3083;
wire net8215;
wire net2435;
wire net10641;
wire net3808;
wire net3698;
wire net3082;
wire net3081;
wire net2565;
wire net3076;
wire net3215;
wire net7151;
wire net3071;
wire net9382;
wire net3949;
wire net3070;
wire net3068;
wire net4842;
wire net6767;
wire net3600;
wire net7306;
wire net3058;
wire net2138;
wire net3057;
wire net2211;
wire net9129;
wire net574;
wire net3431;
wire net3055;
wire net3492;
wire net3053;
wire net5876;
wire net3049;
wire net3047;
wire net8532;
wire net7244;
wire net9217;
wire net3042;
wire net11105;
wire net3039;
wire net6528;
wire net9214;
wire net3036;
wire net3035;
wire net3099;
wire net1258;
wire net3034;
wire net3032;
wire net3030;
wire net10023;
wire net7524;
wire net1080;
wire net3029;
wire net10308;
wire net3028;
wire net3023;
wire net2962;
wire net3021;
wire net3017;
wire net1663;
wire net3016;
wire net9355;
wire net5554;
wire net8932;
wire net3015;
wire net847;
wire net11087;
wire net3014;
wire net4414;
wire net9450;
wire net3011;
wire net3077;
wire net10904;
wire net3010;
wire net5794;
wire net8649;
wire net3006;
wire net411;
wire net10372;
wire net6852;
wire net3005;
wire net3004;
wire net3003;
wire net1704;
wire net11143;
wire net9064;
wire net3002;
wire net3000;
wire net2996;
wire net3158;
wire net7131;
wire net1525;
wire net916;
wire net2989;
wire net9767;
wire net3187;
wire net2022;
wire net5200;
wire net6740;
wire out8;
wire net2987;
wire net1830;
wire net6770;
wire net6251;
wire net2979;
wire net2978;
wire net159;
wire net2975;
wire net10984;
wire net10728;
wire net2972;
wire net2730;
wire net326;
wire net10263;
wire net6700;
wire net7684;
wire net2971;
wire net4955;
wire net3562;
wire net4191;
wire net2969;
wire net3481;
wire net2968;
wire net2967;
wire net1022;
wire net287;
wire net3059;
wire net3118;
wire net10994;
wire net7176;
wire net2954;
wire net2863;
wire net10360;
wire net9247;
wire net2509;
wire net6044;
wire net2950;
wire net2058;
wire net5520;
wire net3458;
wire net2949;
wire net792;
wire net2946;
wire net2714;
wire net2681;
wire net6721;
wire net2941;
wire net2940;
wire net8251;
wire net2939;
wire net11006;
wire net2938;
wire net11135;
wire net2936;
wire net7894;
wire net753;
wire net2932;
wire net2930;
wire net6782;
wire net11232;
wire net6858;
wire net2928;
wire net9245;
wire net5767;
wire net2923;
wire net2921;
wire net2918;
wire net2917;
wire net2915;
wire net1442;
wire net3679;
wire net6584;
wire net2913;
wire net3859;
wire net7155;
wire net5225;
wire net8964;
wire net4032;
wire net2908;
wire net4094;
wire net2903;
wire net4135;
wire net2902;
wire net9122;
wire net2436;
wire net5492;
wire net7918;
wire net4096;
wire net5265;
wire net534;
wire net10421;
wire net3616;
wire net3533;
wire net2891;
wire net11154;
wire net6354;
wire net2886;
wire net5222;
wire net1664;
wire net2878;
wire net2195;
wire net1705;
wire net2877;
wire net8923;
wire net8514;
wire net6667;
wire net10941;
wire net6895;
wire net2875;
wire net1256;
wire net3074;
wire net2872;
wire net7250;
wire net10032;
wire net2870;
wire net4238;
wire net2869;
wire net4437;
wire net4475;
wire net4560;
wire net2595;
wire net8610;
wire net2516;
wire net1992;
wire net9085;
wire net6657;
wire net2847;
wire net461;
wire net6897;
wire net2836;
wire net35;
wire net5199;
wire net4652;
wire net5548;
wire net2988;
wire net2871;
wire net2834;
wire net10753;
wire net8262;
wire net2832;
wire net2831;
wire net4978;
wire net7309;
wire net2829;
wire net3447;
wire net2752;
wire net9097;
wire net5368;
wire net2826;
wire net2818;
wire net3714;
wire net6357;
wire net2817;
wire net4128;
wire net7971;
wire net2811;
wire net3116;
wire net2807;
wire net5561;
wire net7900;
wire net5735;
wire net2806;
wire net6496;
wire net3467;
wire net8494;
wire net2705;
wire net2801;
wire net2800;
wire net5443;
wire net9203;
wire net2798;
wire net2796;
wire net9813;
wire net3655;
wire net2793;
wire net9567;
wire net3342;
wire net7107;
wire net2790;
wire net8379;
wire net1631;
wire net3710;
wire net1568;
wire net4512;
wire net3995;
wire net3133;
wire net7310;
wire net2784;
wire net2781;
wire net8907;
wire net3831;
wire net4138;
wire net2402;
wire net2777;
wire net3162;
wire net2145;
wire net9270;
wire net146;
wire net2952;
wire net11211;
wire net11104;
wire net802;
wire net2767;
wire net2766;
wire net5588;
wire net3306;
wire net9639;
wire net6689;
wire net9577;
wire net6806;
wire net2763;
wire net945;
wire net4085;
wire net5372;
wire net5432;
wire net2758;
wire net2756;
wire net2749;
wire net923;
wire net3961;
wire net2747;
wire net9465;
wire net9267;
wire net690;
wire net3203;
wire net9249;
wire net1601;
wire net2743;
wire net10761;
wire net3950;
wire net6240;
wire net5193;
wire net6601;
wire net2742;
wire net4666;
wire net8620;
wire net5801;
wire net6272;
wire net3388;
wire net2368;
wire net3528;
wire net585;
wire net3212;
wire net5397;
wire net2738;
wire net2495;
wire net1173;
wire net4323;
wire net10606;
wire net7324;
wire net2733;
wire net6028;
wire net7701;
wire net2000;
wire net3276;
wire net7372;
wire net2723;
wire net8912;
wire net2722;
wire net2720;
wire net10573;
wire net1215;
wire net5480;
wire net11222;
wire net2707;
wire net5675;
wire net6569;
wire net2700;
wire net777;
wire net3980;
wire net2694;
wire net3516;
wire net1508;
wire net9965;
wire net2622;
wire net7354;
wire net1197;
wire net2691;
wire net2689;
wire out4;
wire net795;
wire net2684;
wire net10196;
wire net8508;
wire net2680;
wire net3348;
wire net2497;
wire net2679;
wire net2674;
wire net1459;
wire net2873;
wire net2760;
wire net2666;
wire net10034;
wire net3612;
wire net3221;
wire net5313;
wire net2663;
wire net3811;
wire net9426;
wire net105;
wire net2659;
wire net10731;
wire net2658;
wire net10026;
wire net407;
wire net3268;
wire net4808;
wire net2657;
wire net2653;
wire net2381;
wire net2652;
wire net2650;
wire net1934;
wire net2649;
wire net9023;
wire net2648;
wire net1786;
wire net1037;
wire net2791;
wire net2642;
wire net454;
wire net4528;
wire net2634;
wire net4608;
wire net2631;
wire net2626;
wire net2772;
wire net2625;
wire net6280;
wire net10920;
wire net6302;
wire net3202;
wire net4113;
wire net10351;
wire net6979;
wire net4964;
wire net9620;
wire net2620;
wire net9745;
wire net3199;
wire net2618;
wire net626;
wire net6673;
wire net1800;
wire net3346;
wire net231;
wire net3251;
wire net3964;
wire net7034;
wire net9446;
wire net6600;
wire net9137;
wire net2782;
wire net2610;
wire net2603;
wire net11164;
wire net361;
wire net4086;
wire net2601;
wire net2600;
wire net662;
wire net8778;
wire net2596;
wire net3802;
wire net2591;
wire net9530;
wire net276;
wire net8828;
wire net2588;
wire net4819;
wire net2586;
wire net2014;
wire net9451;
wire net2232;
wire net2375;
wire net6123;
wire net2583;
wire net2581;
wire net3775;
wire in17;
wire net9990;
wire net4650;
wire net2579;
wire net2695;
wire net5839;
wire net7961;
wire net3579;
wire net2960;
wire net2576;
wire net2574;
wire net9799;
wire net6922;
wire net2571;
wire net2569;
wire net10851;
wire net9491;
wire net3031;
wire net2568;
wire net1575;
wire net7799;
wire net3153;
wire net10775;
wire net10540;
wire net2655;
wire net4907;
wire net8765;
wire net7623;
wire net6843;
wire net2566;
wire net2563;
wire net10810;
wire net5332;
wire net2561;
wire net6644;
wire net7476;
wire net2557;
wire net2555;
wire net1597;
wire net6793;
wire net2543;
wire net2672;
wire net2542;
wire net2541;
wire net1241;
wire net7612;
wire net5883;
wire net2538;
wire net1544;
wire net5457;
wire net8325;
wire net2536;
wire net7801;
wire net5933;
wire net2535;
wire net1563;
wire net5098;
wire net10405;
wire net2534;
wire net2532;
wire net2208;
wire net2527;
wire net9904;
wire net1688;
wire net10783;
wire net7965;
wire net3624;
wire net10752;
wire net7898;
wire net2524;
wire net8891;
wire net4747;
wire net6618;
wire net6545;
wire net2521;
wire net2520;
wire net4532;
wire net2519;
wire net2518;
wire net2241;
wire net2517;
wire net3586;
wire net2504;
wire net3247;
wire net1203;
wire net2502;
wire net2500;
wire net2499;
wire net3581;
wire net8543;
wire net3392;
wire net5312;
wire net2491;
wire net2487;
wire net2482;
wire net2956;
wire net5093;
wire net9733;
wire net3560;
wire net6660;
wire net5692;
wire net6542;
wire net2480;
wire net2479;
wire net2478;
wire net7750;
wire net2476;
wire net1592;
wire net8987;
wire net65;
wire net2645;
wire net5245;
wire net1613;
wire net5690;
wire net6619;
wire net5238;
wire net9687;
wire net8485;
wire net2469;
wire net2115;
wire net2896;
wire net734;
wire net2460;
wire net2459;
wire net7302;
wire net2453;
wire net2452;
wire net5022;
wire net2448;
wire net1460;
wire net2660;
wire net8711;
wire net2444;
wire net7938;
wire net2442;
wire net2233;
wire net2440;
wire net2439;
wire net8935;
wire net2438;
wire net3470;
wire net2842;
wire net2951;
wire net2498;
wire net2033;
wire net2431;
wire net8457;
wire net1888;
wire net8948;
wire net870;
wire net2429;
wire net6532;
wire net2810;
wire net4108;
wire net2425;
wire net2424;
wire net2422;
wire net8825;
wire net4444;
wire net10998;
wire net3155;
wire net208;
wire net4180;
wire net8614;
wire net2421;
wire net604;
wire net10632;
wire net3300;
wire net178;
wire net6745;
wire net2416;
wire net2525;
wire net5067;
wire net2413;
wire net1446;
wire net2412;
wire net2411;
wire net7182;
wire net2408;
wire net7972;
wire net2407;
wire net1914;
wire net912;
wire net2404;
wire net2401;
wire net2400;
wire net4607;
wire net6249;
wire net2399;
wire net2397;
wire net2391;
wire net1477;
wire net2390;
wire net10055;
wire net2389;
wire net2388;
wire net6522;
wire net2386;
wire net2385;
wire net10294;
wire net5806;
wire net1181;
wire net2379;
wire net10872;
wire net2378;
wire net1848;
wire net2377;
wire net3619;
wire net2840;
wire net2271;
wire net1611;
wire net7895;
wire net6720;
wire net2370;
wire net2364;
wire net8578;
wire net1520;
wire net10417;
wire net2362;
wire net4204;
wire net2361;
wire net3850;
wire net7431;
wire net2356;
wire net2353;
wire net2724;
wire net10508;
wire net3803;
wire net2352;
wire net3148;
wire net1139;
wire net10990;
wire net10223;
wire net2351;
wire net9104;
wire net6705;
wire net9714;
wire net2349;
wire net7085;
wire net8293;
wire net2718;
wire net8501;
wire net2347;
wire net2383;
wire net2345;
wire net2858;
wire net2344;
wire net2343;
wire net4250;
wire net8756;
wire net7387;
wire net2338;
wire net5430;
wire net2335;
wire net2334;
wire net9368;
wire net3163;
wire net9425;
wire net2006;
wire net1463;
wire net8465;
wire net3541;
wire net8033;
wire net7738;
wire net7281;
wire net9782;
wire net2326;
wire net9041;
wire net2325;
wire net2317;
wire net5091;
wire net1747;
wire net10289;
wire net8990;
wire net8169;
wire net138;
wire net365;
wire net2312;
wire net9060;
wire net2309;
wire net3413;
wire net7009;
wire net1640;
wire net3668;
wire net4457;
wire net2302;
wire net1118;
wire net390;
wire net2528;
wire net2296;
wire net10302;
wire net1738;
wire net1030;
wire net10925;
wire net10507;
wire net2292;
wire net10261;
wire net3124;
wire net2291;
wire net6097;
wire net11031;
wire net2290;
wire net762;
wire net5890;
wire net6968;
wire net2307;
wire net6281;
wire net2287;
wire net8361;
wire net5202;
wire net9096;
wire net1909;
wire net3885;
wire net133;
wire net216;
wire net1261;
wire net7417;
wire net2716;
wire net2280;
wire net2846;
wire net2279;
wire net2426;
wire net164;
wire net8067;
wire net2830;
wire net2275;
wire net4011;
wire net2274;
wire net2719;
wire net3269;
wire net5030;
wire net3623;
wire net2276;
wire net2272;
wire net3305;
wire net6714;
wire net2269;
wire net1596;
wire net2735;
wire net3307;
wire net2263;
wire net5075;
wire net10770;
wire net5670;
wire net2904;
wire net4118;
wire net2262;
wire net2259;
wire net7193;
wire net2252;
wire net2251;
wire net2249;
wire net5984;
wire net2248;
wire net4790;
wire net2247;
wire net1116;
wire net11199;
wire net11147;
wire net2245;
wire net10880;
wire net2765;
wire net2244;
wire net2243;
wire net6625;
wire net2242;
wire net2240;
wire net3295;
wire net1713;
wire net2238;
wire net2237;
wire net7221;
wire net8789;
wire net179;
wire net1571;
wire net2230;
wire net2229;
wire net8930;
wire net4272;
wire net2277;
wire net7690;
wire net5572;
wire net3066;
wire net5626;
wire net3554;
wire net2226;
wire net4116;
wire net5499;
wire net3310;
wire net2224;
wire net10476;
wire net2222;
wire net11002;
wire net1865;
wire net6178;
wire net2219;
wire net10483;
wire net8504;
wire net2313;
wire net4206;
wire net1822;
wire net6485;
wire net1975;
wire net2204;
wire net10714;
wire net3527;
wire net4196;
wire net5105;
wire net2192;
wire net2191;
wire net2187;
wire net4006;
wire net2184;
wire net5908;
wire net7483;
wire net2182;
wire net2741;
wire net7975;
wire net327;
wire net9065;
wire net3103;
wire net3291;
wire net4844;
wire net2174;
wire net2172;
wire net3836;
wire net7300;
wire net10198;
wire net3522;
wire net2171;
wire net2165;
wire net2164;
wire net2163;
wire net4775;
wire net2162;
wire net5017;
wire net2161;
wire net1340;
wire net9274;
wire net5607;
wire net6579;
wire net2160;
wire net1208;
wire net9312;
wire net2157;
wire in5;
wire net396;
wire net2154;
wire net7899;
wire net7231;
wire net7184;
wire net2152;
wire net2151;
wire net3890;
wire net2149;
wire net2144;
wire net10357;
wire net7358;
wire net9482;
wire net2493;
wire net6435;
wire net2142;
wire net9554;
wire net8370;
wire net6595;
wire net2135;
wire net10684;
wire net2134;
wire net9017;
wire net7551;
wire net853;
wire net8461;
wire net3250;
wire net5382;
wire net8645;
wire net8467;
wire net2354;
wire net2822;
wire net2693;
wire net8403;
wire net5638;
wire net2137;
wire net3643;
wire net2129;
wire net4315;
wire net10158;
wire net9890;
wire net3120;
wire net2126;
wire net5891;
wire net2125;
wire net3436;
wire net1876;
wire net1741;
wire net2123;
wire net219;
wire net2120;
wire net3752;
wire net794;
wire net4363;
wire net1069;
wire net8957;
wire net1365;
wire net6606;
wire net10970;
wire net10614;
wire net7866;
wire net2114;
wire net2113;
wire net2111;
wire net10696;
wire net2108;
wire net2106;
wire net2710;
wire net343;
wire net2105;
wire net8120;
wire net2270;
wire net1809;
wire net10556;
wire net2102;
wire net292;
wire net2881;
wire net3496;
wire net9994;
wire net2101;
wire net2959;
wire net2097;
wire net2708;
wire net2096;
wire net330;
wire net1219;
wire net5507;
wire net2474;
wire net2094;
wire net9557;
wire net6868;
wire net9956;
wire net2088;
wire net2086;
wire net8380;
wire net3267;
wire net8960;
wire net2508;
wire net10500;
wire net2085;
wire net2215;
wire net6537;
wire net2570;
wire net655;
wire net2084;
wire net2041;
wire net503;
wire net2078;
wire net6248;
wire net2180;
wire net3989;
wire net9523;
wire net8730;
wire net6946;
wire net3237;
wire net2073;
wire net2393;
wire net2072;
wire net2970;
wire net2068;
wire net2064;
wire net5702;
wire net9929;
wire net212;
wire net2061;
wire net9034;
wire net7853;
wire net2060;
wire net4319;
wire net9520;
wire net3308;
wire net2057;
wire net3626;
wire net8627;
wire net2054;
wire net425;
wire net3381;
wire net2769;
wire net1796;
wire net2010;
wire net4329;
wire net2859;
wire net2048;
wire net515;
wire net2045;
wire net2265;
wire net6350;
wire net6908;
wire net2042;
wire net7969;
wire net2039;
wire net2037;
wire net1958;
wire net2032;
wire net2246;
wire net1155;
wire net1429;
wire net7716;
wire net2026;
wire net1170;
wire net4754;
wire net2023;
wire net2725;
wire net177;
wire net2021;
wire net10100;
wire net2210;
wire net1368;
wire net7968;
wire net4415;
wire net6395;
wire net10076;
wire net7867;
wire net2019;
wire net6594;
wire net2018;
wire net2016;
wire net2332;
wire net211;
wire net11070;
wire net6226;
wire net2015;
wire net2776;
wire net8445;
wire net7359;
wire net2007;
wire net9162;
wire net2005;
wire net3248;
wire net2001;
wire net430;
wire net2098;
wire net1998;
wire net1997;
wire net1853;
wire net750;
wire net5278;
wire net2948;
wire net6708;
wire net1994;
wire net3762;
wire net6194;
wire net2040;
wire net1993;
wire net2009;
wire net310;
wire net10150;
wire net8311;
wire net6727;
wire net2506;
wire net1991;
wire net6892;
wire net10983;
wire net2104;
wire net763;
wire net3738;
wire net1190;
wire net1989;
wire net6776;
wire net4922;
wire net3080;
wire net1985;
wire net8392;
wire net744;
wire net9941;
wire net1984;
wire net350;
wire net3726;
wire net8951;
wire net4254;
wire net1983;
wire net1291;
wire net3955;
wire net1977;
wire net1308;
wire net1974;
wire net1754;
wire net4034;
wire net11122;
wire net8174;
wire net255;
wire net11114;
wire net2792;
wire net5576;
wire net2255;
wire net2572;
wire net1466;
wire net2890;
wire net3967;
wire net2505;
wire net5367;
wire net5369;
wire net1967;
wire net1964;
wire net2985;
wire net1961;
wire net2845;
wire net1960;
wire net9481;
wire net6332;
wire net1959;
wire net1956;
wire net2197;
wire net2471;
wire net3416;
wire net6025;
wire net10278;
wire net9173;
wire net2974;
wire net4137;
wire net1948;
wire net1946;
wire net10950;
wire net2510;
wire net1945;
wire net2567;
wire net1943;
wire net1942;
wire net1940;
wire net1939;
wire net10909;
wire net6218;
wire net9624;
wire net8447;
wire net2841;
wire net10768;
wire net1937;
wire net4937;
wire net861;
wire net9036;
wire net3338;
wire net2823;
wire net2545;
wire net1931;
wire net5031;
wire net9417;
wire net6115;
wire net8134;
wire net5493;
wire net6598;
wire net1923;
wire net1922;
wire net970;
wire net1921;
wire net9485;
wire net5558;
wire net6316;
wire net2214;
wire net1913;
wire net1912;
wire net7378;
wire net4812;
wire net1767;
wire net2933;
wire net8654;
wire net2888;
wire net1903;
wire net8925;
wire net1899;
wire net1897;
wire net8327;
wire net999;
wire net10931;
wire net6429;
wire net1896;
wire net3705;
wire net1555;
wire net4107;
wire net1895;
wire net3090;
wire net1894;
wire net10052;
wire net1889;
wire net6166;
wire net2257;
wire net7606;
wire net7259;
wire net3337;
wire net2585;
wire net1293;
wire net8608;
wire net3279;
wire net2036;
wire net1887;
wire net10617;
wire net10399;
wire net4647;
wire net2398;
wire net1884;
wire net1883;
wire net294;
wire net5749;
wire net1864;
wire net1861;
wire net500;
wire net1857;
wire net1856;
wire net1855;
wire net172;
wire net9028;
wire net4174;
wire net3681;
wire net1854;
wire net10599;
wire net2599;
wire net10868;
wire net1850;
wire net4570;
wire net4948;
wire net2337;
wire net1849;
wire net10393;
wire net10206;
wire net686;
wire net7290;
wire net3371;
wire net1846;
wire net904;
wire net442;
wire net10319;
wire net5192;
wire net1842;
wire net1841;
wire net3209;
wire net4044;
wire net1908;
wire net11111;
wire net1840;
wire net6462;
wire net11140;
wire net1838;
wire net10926;
wire net7573;
wire net1851;
wire net1837;
wire net2503;
wire net5678;
wire net6907;
wire net8994;
wire net1835;
wire net8773;
wire net4422;
wire net1826;
wire net6058;
wire net1556;
wire net5253;
wire net5612;
wire net10281;
wire net1819;
wire net10792;
wire net1817;
wire net3530;
wire net340;
wire net3194;
wire net1813;
wire net3652;
wire net3378;
wire net3084;
wire net1501;
wire net5756;
wire net2261;
wire net3242;
wire net10986;
wire net4839;
wire net2110;
wire net1029;
wire net4802;
wire net3884;
wire net4846;
wire net1811;
wire net313;
wire net4172;
wire net3317;
wire net10661;
wire net2076;
wire net1806;
wire net5508;
wire net2628;
wire net776;
wire net10491;
wire net2740;
wire net2575;
wire net1802;
wire net5989;
wire net10197;
wire net6467;
wire net3349;
wire net9497;
wire net2494;
wire net1795;
wire net1318;
wire net6297;
wire net2305;
wire net1792;
wire net9409;
wire net8430;
wire net977;
wire net1791;
wire net2761;
wire net4700;
wire net335;
wire net9367;
wire net6934;
wire net4229;
wire net5823;
wire net5924;
wire net3105;
wire net5556;
wire net7922;
wire net4684;
wire net4863;
wire net7955;
wire net6555;
wire net2704;
wire net9787;
wire net6159;
wire net8151;
wire net1780;
wire net1775;
wire net6976;
wire net3593;
wire net3195;
wire net1654;
wire net1774;
wire net9636;
wire net3503;
wire net2754;
wire net1987;
wire net5674;
wire net10901;
wire net1771;
wire net7335;
wire net1770;
wire net11113;
wire net3362;
wire net1769;
wire net5172;
wire net1768;
wire net8830;
wire net6197;
wire net6960;
wire net8356;
wire net1766;
wire net9800;
wire net1763;
wire net10452;
wire net2816;
wire net2329;
wire net1759;
wire net9143;
wire net4236;
wire net1757;
wire net2481;
wire net2874;
wire net2753;
wire net3233;
wire net1749;
wire net7374;
wire net5621;
wire net4618;
wire net6531;
wire net2295;
wire net1372;
wire net8170;
wire net114;
wire net8111;
wire net5914;
wire net1742;
wire net5768;
wire net1739;
wire net6451;
wire net4815;
wire net9517;
wire net6574;
wire net3462;
wire net1734;
wire net1733;
wire net2640;
wire net1732;
wire net483;
wire net7916;
wire net1731;
wire net6664;
wire net5288;
wire net1730;
wire net8840;
wire net4280;
wire net4813;
wire net1729;
wire net2731;
wire net1726;
wire net5147;
wire net1725;
wire net4803;
wire net1724;
wire net9942;
wire net5446;
wire net9494;
wire net1723;
wire net116;
wire net28;
wire net1722;
wire net22;
wire net10588;
wire net6838;
wire net7744;
wire net1721;
wire net9272;
wire net8602;
wire net8086;
wire net2892;
wire net1720;
wire net11032;
wire net1716;
wire net578;
wire net11178;
wire net1179;
wire net8070;
wire net5858;
wire net5816;
wire net1040;
wire net3220;
wire net246;
wire net783;
wire net1828;
wire net43;
wire net541;
wire net6604;
wire net4828;
wire net3693;
wire net3037;
wire net8107;
wire net2253;
wire net1941;
wire net6651;
wire net772;
wire net7059;
wire net10751;
wire net2643;
wire net761;
wire net8952;
wire net478;
wire net15;
wire net8383;
wire net4301;
wire net9397;
wire net5025;
wire net746;
wire net168;
wire net2827;
wire net6160;
wire net738;
wire net10713;
wire net1938;
wire net5560;
wire net3204;
wire net9435;
wire net9285;
wire net1638;
wire net737;
wire net1125;
wire net10819;
wire net2879;
wire net3293;
wire net10972;
wire net5458;
wire net4904;
wire net7327;
wire net9993;
wire net736;
wire net11076;
wire net1785;
wire net414;
wire net5344;
wire net1122;
wire net2696;
wire net7078;
wire net2559;
wire net7462;
wire net730;
wire net4917;
wire net3146;
wire out9;
wire net2617;
wire net728;
wire net3599;
wire net406;
wire net9396;
wire net5624;
wire net1999;
wire net4156;
wire net725;
wire net4517;
wire net808;
wire net2732;
wire net2392;
wire net724;
wire net6546;
wire net1526;
wire net2787;
wire net2220;
wire net721;
wire net10946;
wire net9889;
wire net7315;
wire net3632;
wire net7661;
wire net1315;
wire net1814;
wire net797;
wire net7548;
wire net1502;
wire net4756;
wire net1475;
wire net715;
wire net1100;
wire net1689;
wire net4316;
wire net9461;
wire net1178;
wire net4708;
wire net3046;
wire net703;
wire net1519;
wire net679;
wire net9550;
wire net1265;
wire net9928;
wire net3552;
wire net700;
wire net4170;
wire net3666;
wire net699;
wire net1075;
wire net706;
wire net4789;
wire net596;
wire net25;
wire net691;
wire net1488;
wire net5351;
wire net2906;
wire net10037;
wire net676;
wire net3078;
wire net7683;
wire net2258;
wire net6107;
wire net1051;
wire net960;
wire net8894;
wire net8274;
wire net2887;
wire net6641;
wire net693;
wire net2515;
wire net914;
wire net1264;
wire net7379;
wire net2446;
wire net670;
wire net7672;
wire net397;
wire net5387;
wire net7054;
wire net6940;
wire net2668;
wire net1218;
wire net6954;
wire net1656;
wire net4962;
wire net1660;
wire net1773;
wire net648;
wire net842;
wire net153;
wire net644;
wire net1418;
wire net5248;
wire net3008;
wire net1373;
wire net640;
wire net4841;
wire net1827;
wire net5348;
wire net5070;
wire net3389;
wire net1797;
wire net282;
wire net6311;
wire net10541;
wire net7166;
wire net637;
wire net2692;
wire net3977;
wire net2038;
wire net1947;
wire net7261;
wire net238;
wire net1383;
wire net7349;
wire net3024;
wire net579;
wire net2604;
wire net713;
wire net4766;
wire net2083;
wire net707;
wire net559;
wire net5884;
wire net632;
wire net8299;
wire net770;
wire net8949;
wire net2188;
wire net3409;
wire net1331;
wire net4499;
wire net2578;
wire net2651;
wire net631;
wire net611;
wire net9793;
wire net4899;
wire net1146;
wire net617;
wire net986;
wire net1615;
wire net6368;
wire net6816;
wire net7109;
wire net817;
wire net4176;
wire net3504;
wire net3355;
wire net2409;
wire net2544;
wire net603;
wire net9202;
wire net4290;
wire net3063;
wire net1153;
wire net599;
wire net8439;
wire net328;
wire net766;
wire net6707;
wire net3454;
wire net7026;
wire net1573;
wire net2608;
wire net591;
wire net996;
wire net6373;
wire net2260;
wire net2973;
wire net4591;
wire net1113;
wire net2475;
wire net587;
wire net934;
wire net1863;
wire net3920;
wire net9401;
wire net1415;
wire net10701;
wire net7698;
wire net6205;
wire net8419;
wire net3608;
wire net5881;
wire net7868;
wire net1560;
wire net650;
wire net7877;
wire net6824;
wire net58;
wire net8484;
wire net3217;
wire net9241;
wire net8843;
wire net5268;
wire net85;
wire net3027;
wire net4266;
wire net9615;
wire net4927;
wire net4347;
wire net7363;
wire net4143;
wire net186;
wire net8259;
wire net3073;
wire net1882;
wire net1393;
wire net9853;
wire net4348;
wire net710;
wire net3249;
wire net4529;
wire net1976;
wire net612;
wire net1010;
wire net957;
wire net5236;
wire net573;
wire net864;
wire net4998;
wire net3060;
wire net4745;
wire net3056;
wire net357;
wire net1965;
wire net768;
wire net1014;
wire net1681;
wire net8977;
wire net247;
wire net1687;
wire net5889;
wire net4282;
wire net564;
wire net3914;
wire net4577;
wire net6879;
wire net2020;
wire net1772;
wire net4498;
wire net189;
wire net5191;
wire net383;
wire net2788;
wire net1673;
wire net3782;
wire net555;
wire net1379;
wire net3737;
wire net553;
wire net2205;
wire net6826;
wire net9044;
wire net2636;
wire net7294;
wire net551;
wire net10407;
wire net8130;
wire net4390;
wire net1063;
wire net549;
wire net10258;
wire net3595;
wire net1428;
wire net6792;
wire net6363;
wire net546;
wire net2580;
wire net6680;
wire net5961;
wire net544;
wire net6353;
wire net3262;
wire net11184;
wire net9410;
wire net4896;
wire net3661;
wire net1;
wire net7385;
wire net10923;
wire net2602;
wire in3;
wire net1270;
wire net4584;
wire net10879;
wire net2584;
wire net896;
wire net7402;
wire net2029;
wire net535;
wire net3168;
wire net1552;
wire net9453;
wire net2729;
wire net2726;
wire net642;
wire net2159;
wire net659;
wire net830;
wire net3610;
wire net4431;
wire net729;
wire net3379;
wire net823;
wire net1250;
wire net2117;
wire net10726;
wire net1695;
wire net3860;
wire net1886;
wire net1468;
wire net7830;
wire net3445;
wire net98;
wire net524;
wire net4001;
wire net876;
wire net1052;
wire net3587;
wire net3333;
wire net5180;
wire net2079;
wire net9509;
wire net2953;
wire net297;
wire net10006;
wire net8729;
wire net5055;
wire net516;
wire net2779;
wire net1472;
wire net1793;
wire net6982;
wire net8290;
wire net7552;
wire net514;
wire net10732;
wire net8942;
wire net511;
wire net4685;
wire net3618;
wire net1335;
wire net5148;
wire net4151;
wire net685;
wire net107;
wire net2539;
wire net3881;
wire net269;
wire net9652;
wire net346;
wire net8575;
wire net510;
wire net7122;
wire net1233;
wire net1025;
wire net506;
wire net927;
wire net3100;
wire net333;
wire net9466;
wire net3062;
wire net3214;
wire net1927;
wire net975;
wire net1952;
wire net505;
wire net2864;
wire net9804;
wire net8629;
wire net8256;
wire net3550;
wire net6150;
wire net1376;
wire net2630;
wire net1409;
wire net3696;
wire net1437;
wire net1829;
wire net1032;
wire net9595;
wire net8255;
wire net3086;
wire net501;
wire net2931;
wire net3407;
wire net1481;
wire net652;
wire net495;
wire net7364;
wire net494;
wire net988;
wire net492;
wire net2143;
wire net489;
wire net485;
wire net2745;
wire net985;
wire net488;
wire net10878;
wire net646;
wire net838;
wire net5396;
wire net2170;
wire net475;
wire net6502;
wire net8275;
wire net2209;
wire net639;
wire net674;
wire net525;
wire net3400;
wire net7875;
wire net474;
wire net3094;
wire net4975;
wire net1867;
wire net8834;
wire net473;
wire net10822;
wire net6157;
wire net2955;
wire net1145;
wire net4658;
wire net472;
wire net3331;
wire net3340;
wire net1347;
wire net3101;
wire net3958;
wire net3707;
wire net2616;
wire net3061;
wire net2331;
wire net967;
wire net5346;
wire net6035;
wire net3646;
wire net7051;
wire net1057;
wire net2675;
wire net1567;
wire net1272;
wire net2176;
wire net10410;
wire net4372;
wire net8014;
wire net780;
wire net7202;
wire net364;
wire net3395;
wire net1266;
wire net8121;
wire net7904;
wire net5097;
wire net6057;
wire net4099;
wire net5582;
wire net283;
wire net6856;
wire net9353;
wire net3289;
wire net10208;
wire net6002;
wire net2737;
wire net3127;
wire net1114;
wire net9066;
wire net3972;
wire net1295;
wire net10444;
wire net2056;
wire net3832;
wire net9408;
wire net3965;
wire net3159;
wire net459;
wire net545;
wire net6003;
wire net4225;
wire net453;
wire net624;
wire net629;
wire net731;
wire net450;
wire net7946;
wire net448;
wire net5559;
wire net1196;
wire net2122;
wire net5363;
wire net5;
wire net10649;
wire net8898;
wire net1012;
wire net4443;
wire net10884;
wire net3285;
wire net3944;
wire net9006;
wire net1074;
wire net2216;
wire net3704;
wire net561;
wire net7484;
wire net444;
wire net8656;
wire net2638;
wire net2071;
wire net1374;
wire net3621;
wire net10389;
wire net8950;
wire net8904;
wire net504;
wire net2997;
wire net336;
wire net280;
wire net8881;
wire net969;
wire net437;
wire net4483;
wire net7764;
wire net3064;
wire net3631;
wire net8926;
wire net162;
wire net1017;
wire net4787;
wire net10315;
wire net718;
wire net10772;
wire net6725;
wire net2430;
wire net4893;
wire net3095;
wire net5764;
wire net3900;
wire net10383;
wire net8612;
wire net432;
wire net1761;
wire net5294;
wire net8706;
wire net2118;
wire net1645;
wire net428;
wire net774;
wire net556;
wire net3312;
wire net2706;
wire net7487;
wire net771;
wire net5184;
wire net5648;
wire net928;
wire net1336;
wire net1220;
wire net5235;
wire net3033;
wire net293;
wire net2324;
wire net2107;
wire net5829;
wire net689;
wire net7218;
wire net422;
wire net1743;
wire clk;
wire net5308;
wire net2637;
wire net3122;
wire net6691;
wire net3576;
wire net4327;
wire net382;
wire net563;
wire net5841;
wire net1188;
wire net3663;
wire net5465;
wire net758;
wire net8650;
wire net2746;
wire net1625;
wire net417;
wire net901;
wire net10547;
wire net2030;
wire net3791;
wire net415;
wire net4389;
wire net5217;
wire net3142;
wire net4781;
wire net412;
wire net748;
wire net1224;
wire net2299;
wire net9118;
wire net702;
wire net5077;
wire net7425;
wire net634;
wire net1981;
wire net3838;
wire net7610;
wire net5879;
wire net554;
wire net4216;
wire net9725;
wire net1192;
wire net6786;
wire net7583;
wire net2597;
wire net3939;
wire net10846;
wire net8071;
wire net3026;
wire net3721;
wire net4454;
wire net680;
wire net2677;
wire net6442;
wire net6797;
wire net403;
wire net4296;
wire net2066;
wire net2943;
wire net4852;
wire net8878;
wire net7053;
wire net1330;
wire net3216;
wire net3274;
wire net9128;
wire net5131;
wire net854;
wire net10722;
wire net8922;
wire net2656;
wire net4833;
wire net5512;
wire net8320;
wire net1678;
wire net1236;
wire net3397;
wire net166;
wire net1621;
wire net6466;
wire net388;
wire net402;
wire net387;
wire net2924;
wire net1097;
wire net3565;
wire net4489;
wire net4243;
wire net1874;
wire net385;
wire in21;
wire net10671;
wire net10304;
wire net9818;
wire net5303;
wire net2825;
wire net384;
wire net2050;
wire net2456;
wire net885;
wire net2234;
wire net3639;
wire net2156;
wire net8655;
wire net207;
wire net317;
wire net7528;
wire net3273;
wire net1089;
wire net4610;
wire net5482;
wire net6548;
wire net10078;
wire net1666;
wire net4400;
wire net1277;
wire net2298;
wire net155;
wire net1087;
wire net2070;
wire net3858;
wire net3344;
wire net3568;
wire net5048;
wire net2934;
wire net1034;
wire in8;
wire net4370;
wire net4449;
wire net10361;
wire net4818;
wire net6296;
wire net759;
wire net10892;
wire net1518;
wire net2089;
wire net3399;
wire net5358;
wire net152;
wire net139;
wire net5987;
wire net895;
wire net1249;
wire net3651;
wire net742;
wire net8947;
wire net2759;
wire net2893;
wire net4689;
wire net9642;
wire net5682;
wire net2533;
wire net3680;
wire net2025;
wire net10834;
wire net132;
wire net7713;
wire net1221;
wire net862;
wire net131;
wire net6498;
wire net733;
wire net2673;
wire net129;
wire net2529;
wire net4453;
wire net5780;
wire net10513;
wire net7044;
wire net3418;
wire net633;
wire net318;
wire net2304;
wire net9486;
wire net8772;
wire net7029;
wire net810;
wire net6735;
wire net6853;
wire net6986;
wire net258;
wire net10207;
wire net2789;
wire net3115;
wire net5563;
wire net123;
wire net592;
wire net7466;
wire net117;
wire net3973;
wire net9553;
wire net121;
wire net10721;
wire net5976;
wire net1297;
wire net0;
wire net3167;
wire net4303;
wire net8985;
wire net1982;
wire net10130;
wire net3403;
wire net462;
wire net653;
wire net3682;
wire net5759;
wire net1617;
wire net4306;
wire net285;
wire net600;
wire net5877;
wire net1234;
wire net7821;
wire net2236;
wire net1043;
wire net8020;
wire net4579;
wire net2995;
wire net11004;
wire net9936;
wire net73;
wire net10947;
wire net4401;
wire net825;
wire net4402;
wire net10019;
wire net1765;
wire net113;
wire net2550;
wire net6089;
wire net752;
wire net3290;
wire net1332;
wire net309;
wire net791;
wire net4218;
wire net7370;
wire net538;
wire net833;
wire net8592;
wire in13;
wire net10065;
wire net4239;
wire net311;
wire net362;
wire net1226;
wire net978;
wire net2712;
wire net110;
wire net949;
wire net886;
wire net8618;
wire net2374;
wire net890;
wire net4075;
wire net2709;
wire net6153;
wire net69;
wire net8502;
wire net793;
wire net2167;
wire net9779;
wire net846;
wire net1569;
wire net4041;
wire net10374;
wire net627;
wire net59;
wire net717;
wire net3443;
wire net874;
wire net7622;
wire net695;
wire net7467;
wire net1658;
wire net5258;
wire net513;
wire net9946;
wire net6147;
wire net3372;
wire net3113;
wire net6652;
wire net463;
wire net751;
wire net1551;
wire net915;
wire net7145;
wire net103;
wire net5609;
wire net2848;
wire net44;
wire net11166;
wire net849;
wire net100;
wire net97;
wire net2964;
wire net4411;
wire net6095;
wire net1878;
wire net394;
wire net4866;
wire net4993;
wire net3311;
wire net8537;
wire net787;
wire net2819;
wire net239;
wire net10002;
wire net27;
wire net195;
wire net1929;
wire net657;
wire net3945;
wire net94;
wire net1185;
wire net8487;
wire net2067;
wire net6663;
wire in12;
wire net9402;
wire net409;
wire net482;
wire net264;
wire net209;
wire net4683;
wire net582;
wire net3332;
wire net2646;
wire net8694;
wire net6530;
wire net5379;
wire net971;
wire net6921;
wire net88;
wire net1900;
wire net4553;
wire net9403;
wire net3164;
wire net5893;
wire net5243;
wire net735;
wire net99;
wire net3505;
wire net925;
wire net9984;
wire net7880;
wire net5406;
wire net2485;
wire net826;
wire net3179;
wire net199;
wire net2318;
wire net458;
wire net6760;
wire net678;
wire net262;
wire net1287;
wire net4759;
wire net3633;
wire net3571;
wire net1789;
wire net5407;
wire net10852;
wire net87;
wire net11033;
wire net7177;
wire net5568;
wire net290;
wire net66;
wire net8963;
wire net5473;
wire net6737;
wire net5112;
wire net1710;
wire net486;
wire net9969;
wire net9012;
wire net7278;
wire net2357;
wire net1046;
wire net10550;
wire net6360;
wire net857;
wire net81;
wire net3298;
wire net9420;
wire net3420;
wire net2264;
wire net2514;
wire net7216;
wire net6596;
wire net9962;
wire net202;
wire net5040;
wire net2339;
wire net572;
wire net3795;
wire net7728;
wire net1212;
wire net1545;
wire net2428;
wire net11;
wire net3322;
wire net1448;
wire in7;
wire net374;
wire net9296;
wire net4447;
wire net799;
wire net1486;
wire net1707;
wire net4162;
wire net7982;
wire net6356;
wire net2074;
wire net2100;
wire net889;
wire net8835;
wire net877;
wire net490;
wire net1064;
wire net2647;
wire net8640;
wire net298;
wire net467;
wire net241;
wire net851;
wire net9;
wire net1028;
wire net6017;
wire net998;
wire net9943;
wire net3166;
wire net11223;
wire net4373;
wire net160;
wire net1223;
wire net765;
wire net2853;
wire net252;
wire net10101;
wire net8287;
wire net7470;
wire net1603;
wire net31;
wire net288;
wire net2200;
wire net441;
wire net673;
wire net1314;
wire net3402;
wire net2155;
wire net6957;
wire net3236;
wire net2283;
wire net3686;
wire net773;
wire net3391;
wire net4653;
wire net7092;
wire net3303;
wire in6;
wire net4619;
wire net167;
wire net1414;
wire net9712;
wire net2876;
wire net2750;
wire net2189;
wire net9255;
wire net7320;
wire net2330;
wire net891;
wire net5617;
wire net8221;
wire net3304;
wire net8422;
wire net6381;
wire net75;
wire net2053;
wire net2513;
wire net8308;
wire net523;
wire net9082;
wire net2983;
wire net45;
wire net5488;
wire net3171;
wire net4979;
wire net935;
wire net3468;
wire net5603;
wire net4;
wire net9110;
wire net334;
wire net2268;
wire net477;
wire net9844;
wire net1489;
wire net2522;
wire net481;
wire net11175;
wire net3299;
wire net6;
wire net8531;
wire net5913;
wire net665;
wire net2371;
wire net10863;
wire net9609;
wire net1788;
wire net9093;
wire net4362;
wire net5602;
wire net379;
wire net197;
wire net6612;
wire net1387;
wire net10380;
wire net779;
wire net10467;
wire net3414;
wire net106;
wire net8896;
wire net6509;
wire net5350;
wire net995;
wire net7575;
wire net3876;
wire net2451;
wire net566;
wire net1210;
wire net1172;
wire net1498;
wire net7788;
wire net2621;
wire net1419;
wire net2670;
wire net68;
wire net6400;
wire net1405;
wire net7406;
wire net723;
wire net1177;
wire net6344;
wire net1110;
wire net696;
wire net4074;
wire net2008;
wire net8511;
wire net1632;
wire net7069;
wire net8177;
wire net7825;
wire net245;
wire net3192;
wire net1834;
wire net2839;
wire net2396;
wire net6079;
wire net3592;
wire net667;
wire net3452;
wire net18;
wire net1214;
wire net7061;
wire net90;
wire net10165;
wire net5947;
wire net1425;
wire net8;
wire net8609;
wire net1677;
wire net1727;
wire net3460;
wire net2849;
wire net10867;
wire net2688;
wire net2804;
wire net2082;
wire net1443;
wire in23;
wire net3558;
wire net5866;
wire net7907;
wire net7630;
wire net4017;
wire net9646;
wire net9608;
wire net163;
wire net3170;
wire net7414;
wire net51;
wire net5680;
wire net10371;
wire net2034;
wire net5800;
wire net2285;
wire net726;
wire net1165;
wire net11009;
wire net5577;
wire net5748;
wire net7132;
wire net10496;
wire net7800;
wire net347;
wire net5090;
wire net1007;
wire net1408;
wire net6909;
wire net2526;
wire net9637;
wire net4910;
wire net84;
wire net2577;
wire net2667;
wire net6122;
wire net398;
wire net1610;
wire net2363;
wire net7966;
wire net6188;
wire net3128;
wire in4;
wire net3309;
wire net1971;
wire net9526;
wire net240;
wire net9379;
wire net4799;
wire net1885;
wire net175;
wire net682;
wire net570;
wire net1777;
wire net7805;
wire net274;
wire in16;
wire net1549;
wire net4497;
wire net5886;
wire net2308;
wire net1252;
wire net1503;
wire net1676;
wire net5216;
wire net2633;
wire net496;
wire net1055;
wire net426;
wire net8441;
wire net348;
wire net1668;
wire net962;
wire net10420;
wire net36;
wire net4441;
wire net507;
wire net5673;
wire net1338;
wire net2201;
wire net671;
wire net7381;
wire net7491;
wire net3383;
wire net8595;
wire net21;
wire net143;
wire net609;
wire net1421;
wire net920;
wire net6911;
wire net3450;
wire net625;
wire net393;
wire net522;
wire net2463;
wire net1745;
wire in20;
wire net491;
wire net10838;
wire net818;
wire net4988;
wire net300;
wire net157;
wire net2081;
wire net10336;
wire net1935;
wire net95;
wire net7596;
wire net79;
wire net835;
wire net20;
wire net4002;
wire net10079;
wire net86;
wire net601;
wire net2256;
wire net3361;
wire net1530;
wire net3983;
wire net154;
wire net1006;
wire net9930;
wire net4260;
wire net6706;
wire net7658;
wire net1893;
wire net10991;
wire net251;
wire net1420;
wire net5449;
wire in18;
wire net6484;
wire net775;
wire net10989;
wire net10527;
wire net3364;
wire net254;
wire net7646;
wire net64;
wire net8013;
wire net408;
wire net4063;
wire net2530;
wire net2049;
wire net951;
wire net12;
wire net536;
wire net7897;
wire net83;
wire net33;
wire net4167;
wire net1011;
wire net9873;
wire net2150;
wire net185;
wire net5637;
wire net10347;
wire net4738;
wire net5792;
wire net3200;
wire net1820;
wire net10763;
wire net5699;
wire net638;
wire net10698;
wire net8755;
wire net128;
wire net5392;
wire net3176;
wire net2866;
wire net7818;
wire net2980;
wire net4326;
wire net1205;
wire net37;
wire net2384;
wire net7124;
wire net4184;
wire net530;
wire net9391;
wire net5117;
wire net6156;
wire net1511;
wire net38;
wire net3569;
wire net11119;
wire net3630;
wire net127;
wire net7257;
wire net1346;
wire net2814;
wire net569;
wire net10707;
wire net502;
wire net158;
wire net6458;
wire net6724;
wire net3428;
wire net145;
wire net8194;
wire net213;
wire net5936;
wire net7834;
wire net499;
wire net6278;
wire net50;
wire net2128;
wire net6069;
wire net2103;
wire net4945;
wire net7355;
wire net229;
wire net732;
wire net4869;
wire net457;
wire net645;
wire net4668;
wire net1636;
wire net479;
wire net149;
wire net10316;
wire net57;
wire net6006;
wire net984;
wire net8126;
wire net3495;
wire net2838;
wire net3845;
wire net3172;
wire net9284;
wire net137;
wire net2203;
wire net3182;
wire net4960;
wire net7494;
wire net5024;
wire net5436;
wire net5481;
wire net11017;
wire net10809;
wire net9480;
wire net6303;
wire net1586;
wire net3843;
wire net1148;
wire net1168;
wire net10460;
wire net2346;
wire net380;
wire net3197;
wire net359;
wire net993;
wire net191;
wire net755;
wire net47;
wire net5013;
wire net3625;
wire net10971;
wire net1104;
wire net5834;
wire net512;
wire net7282;
wire net3052;
wire net2415;
wire net8743;
wire net7074;
wire net1305;
wire net10760;
wire net13;
wire net3899;
wire net3001;
wire net3421;
wire net89;
wire net2942;
wire net741;
wire net3534;
wire net10063;
wire net3446;
wire net6818;
wire net944;
wire net1714;
wire net5177;
wire net5267;
wire net9489;
wire net3465;
wire net6885;
wire net1213;
wire net1410;
wire net3188;
wire net395;
wire net6733;
wire net2992;
wire net2387;
wire net49;
wire net6702;
wire net7021;
wire net664;
wire net9866;
wire net7618;
wire net296;
wire net10171;
wire net855;
wire net55;
wire net134;
wire net3474;
wire net3585;
wire net1182;
wire net4054;
wire net5928;
wire net6941;
wire net6717;
wire net2212;
wire in1;
wire net74;
wire net4692;
wire net2077;
wire net210;
wire net3254;
wire net4098;
wire net1954;
wire net4211;
wire net1237;
wire net10220;
wire net1317;
wire net9119;
wire net7331;
wire net5977;
wire net176;
wire net80;
wire net756;
wire net1970;
wire net10915;
wire net1858;
wire net9277;
wire net1243;
wire net1284;
wire net2857;
wire net5306;
wire net1639;
wire net852;
wire net3683;
wire net1465;
wire net6064;
wire net3642;
wire net445;
wire net7490;
wire net3785;
wire net5053;
wire net5661;
wire net9686;
wire net8617;
wire net70;
wire net2193;
wire net279;
wire net11173;
wire net3453;
wire net2;
wire net2468;
wire net192;
wire net594;
wire net174;
wire net6092;
wire net560;
wire net1755;
wire net225;
wire net1653;
wire net7705;
wire net265;
wire net6474;
wire net10948;
wire net9186;
wire net1804;
wire net2437;
wire net96;
wire net8230;
wire net3513;
wire net4939;
wire in2;
wire net610;
wire net180;
wire net4252;
wire net550;
wire net4520;
wire net3694;
wire net1542;
wire net3434;
wire net4153;
wire net5132;
wire net1447;
wire net9582;
wire net101;
wire net3784;
wire net3711;
wire net281;
wire net181;
wire net698;
wire net3510;
wire net1986;
wire net2278;
wire net182;
wire net3201;
wire net641;
wire net7604;
wire net6990;
wire net1033;
wire net10919;
wire net7613;
wire net785;
wire net701;
wire net286;
wire net5221;
wire net8742;
wire net2547;
wire net3139;
wire net476;
wire net3393;
wire net722;
wire net1095;
wire net4832;
wire net1803;
wire net301;
wire net1683;
wire net3315;
wire net8573;
wire net2427;
wire net345;
wire net3461;
wire net537;
wire net1881;
wire net10342;
wire net5373;
wire net8759;
wire net7429;
wire net2703;
wire net4460;
wire net966;
wire net4924;
wire net2333;
wire net1016;
wire net8099;
wire net193;
wire net1348;
wire net7042;
wire net48;
wire net8774;
wire net2627;
wire net194;
wire net3927;
wire net4337;
wire net5628;
wire net198;
wire net360;
wire net2833;
wire net2012;
wire net8841;
wire net6549;
wire net6881;
wire net236;
wire net9445;
wire net320;
wire net4304;
wire net295;
wire net204;
wire net3620;
wire net8824;
wire net3174;
wire net3613;
wire net7942;
wire net7692;
wire net3747;
wire net589;
wire net53;
wire net583;
wire net214;
wire net3665;
wire net9882;
wire net6994;
wire net7441;
wire net1262;
wire net10985;
wire net8010;
wire net767;
wire net3797;
wire net7147;
wire net237;
wire net4255;
wire net9848;
wire net480;
wire net5681;
wire net8282;
wire net1901;
wire net924;
wire net9127;
wire net2701;
wire net3898;
wire net3320;
wire net233;
wire net6744;
wire net8482;
wire net3718;
wire net220;
wire net6131;
wire net520;
wire net981;
wire net3892;
wire net7440;
wire net366;
wire net607;
wire net7080;
wire net651;
wire net7768;
wire net620;
wire net6997;
wire net939;
wire net3347;
wire net10454;
wire net4586;
wire net3773;
wire net5152;
wire net1614;
wire net2486;
wire net452;
wire net2372;
wire net2592;
wire net63;
wire net2227;
wire net7139;
wire net10264;
wire net1371;
wire net613;
wire net6914;
wire net760;
wire net7303;
wire net223;
wire net5362;
wire net4996;
wire net897;
wire net908;
wire net438;
wire net10362;
wire net9134;
wire net2994;
wire net2678;
wire net10074;
wire net6517;
wire net8690;
wire net227;
wire net3611;
wire net9021;
wire net7346;
wire in9;
wire net660;
wire net6036;
wire net6414;
wire net542;
wire net2702;
wire net1326;
wire net628;
wire net2914;
wire net9184;
wire net5518;
wire net1748;
wire net526;
wire net1495;
wire net2573;
wire net4605;
wire net10309;
wire net230;
wire net10754;
wire net1492;
wire net3755;
wire net3297;
wire net5186;
wire net577;
wire net5095;
wire net661;
wire net1910;
wire net1467;
wire net10049;
wire net7469;
wire net10897;
wire net4773;
wire net3147;
wire net8167;
wire net2202;
wire net8398;
wire net5061;
wire net4774;
wire net418;
wire net323;
wire net11047;
wire net10245;
wire net552;
wire net2899;
wire net244;
wire net3701;
wire net7782;
wire net7219;
wire net2773;
wire net905;
wire net10686;
wire net338;
wire net672;
wire net3098;
wire net4273;
wire net2865;
wire net1790;
wire net24;
wire net1602;
wire net3640;
wire net801;
wire net2147;
wire net10773;
wire net5087;
wire net249;
wire net8436;
wire net7550;
wire net5218;
wire net8132;
wire net1593;
wire net9246;
wire net3417;
wire net5943;
wire net9619;
wire net6070;
wire net5696;
wire net2132;
wire net10134;
wire net9257;
wire net3915;
wire net5610;
wire net8859;
wire net3463;
wire net518;
wire net3848;
wire net10356;
wire net1499;
wire net2911;
wire net7792;
wire net3605;
wire net5952;
wire net6198;
wire net183;
wire net1434;
wire net272;
wire net1558;
wire net902;
wire net10612;
wire net200;
wire net635;
wire net8829;
wire net8243;
wire net5195;
wire net6256;
wire net3771;
wire net234;
wire net4545;
wire net598;
wire net1538;
wire net4130;
wire net4798;
wire net961;
wire net884;
wire net6277;
wire net487;
wire net6743;
wire net261;
wire net7515;
wire net1253;
wire net315;
wire net9775;
wire net1137;
wire net3441;
wire net1426;
wire net5586;
wire net7680;
wire net493;
wire net263;
wire net2221;
wire net4384;
wire net10059;
wire net8594;
wire net8359;
wire net112;
wire net3923;
wire net6094;
wire net1396;
wire net8906;
wire net2916;
wire net2477;
wire net4120;
wire net2654;
wire net2199;
wire net6423;
wire net5460;
wire net6647;
wire net8386;
wire net663;
wire net10598;
wire net1821;
wire net6421;
wire net372;
wire net8277;
wire net2419;
wire net10156;
wire net7396;
wire net443;
wire net17;
wire net10590;
wire net270;
wire net8616;
wire net7820;
wire net3689;
wire net757;
wire net9635;
wire net1384;
wire net6951;
wire net997;
wire net7962;
wire net5309;
wire net3;
wire net2293;
wire net4636;
wire net727;
wire net10870;
wire net344;
wire net9259;
wire net6063;
wire net9380;
wire net3770;
wire net5906;
wire net9903;
wire net3475;
wire net4763;
wire net1643;
wire net2778;
wire net10973;
wire net5341;
wire net878;
wire net593;
wire net10907;
wire net278;
wire net7700;
wire net3685;
wire net1163;
wire in10;
wire net4961;
wire net436;
wire net10860;
wire net2140;
wire net3374;
wire net4930;
wire net1001;
wire net4179;
wire net7084;
wire net2861;
wire net161;
wire net7544;
wire net5639;
wire net291;
wire net9098;
wire net5966;
wire net11162;
wire net9880;
wire net1595;
wire net1836;
wire net588;
wire net529;
wire net376;
wire net1359;
wire net10122;
wire net4317;
wire net370;
wire net3617;
wire net19;
wire net4884;
wire net5159;
wire net306;
wire net4944;
wire net1717;
wire net1778;
wire net8914;
wire net1026;
wire net10327;
wire net1009;
wire net446;
wire net141;
wire net9940;
wire net8909;
wire net7162;
wire net3009;
wire net1684;
wire net784;
wire net1696;
wire net7775;
wire net3245;
wire net10514;
wire net5108;
wire net1862;
wire net130;
wire net1204;
wire net4821;
wire net9658;
wire net932;
wire net7156;
wire net217;
wire net312;
wire net1018;
wire net332;
wire net1158;
wire net93;
wire net9949;
wire net5315;
wire net7;
wire net10;
wire net2327;
wire net9235;
wire net8734;
wire in22;
wire net2935;
wire net7127;
wire net3007;
wire net2365;
wire net10891;
wire net4868;
wire net9317;
wire net3531;
wire net455;
wire net2855;
wire net423;
wire net958;
wire net3185;
wire net976;
wire net4633;
wire net8503;
wire net2289;
wire net72;
wire net3132;
wire net7858;
wire net221;
wire net965;
wire net337;
wire net4568;
wire net968;
wire net7246;
wire net4507;
wire net7408;
wire net9318;
wire net3577;
wire net1452;
wire net5965;
wire net3676;
wire net2554;
wire net3667;
wire net3270;
wire net3573;
wire net1440;
wire net367;
wire net2821;
wire net597;
wire net3229;
wire net704;
wire net349;
wire net8399;
wire net2556;
wire net1200;
wire net2002;
wire net5497;
wire net9676;
wire net2552;
wire net2805;
wire net10624;
wire net4455;
wire net464;
wire net6712;
wire net1635;
wire net356;
wire net9177;
wire net2815;
wire net8463;
wire net2093;
wire net1823;
wire net9478;
wire net1693;
wire net8054;
wire net2764;
wire net4213;
wire net371;
wire net1756;
wire net859;
wire net4750;
wire net6490;
wire net11130;
wire net4451;
wire net3969;
wire net373;
wire net7936;
wire net4202;
wire net800;
wire net9149;
wire net3628;
wire net2629;
wire net3913;
wire net807;
wire net811;
wire net8505;
wire net812;
wire net9722;
wire net5953;
wire net1059;
wire net813;
wire net5326;
wire net1588;
wire net275;
wire net6019;
wire net7361;
wire net5292;
wire net196;
wire net1925;
wire net3119;
wire net10121;
wire net4840;
wire net6580;
wire net816;
wire net6703;
wire net8591;
wire net2473;
wire net1310;
wire net819;
wire net3745;
wire net822;
wire net1528;
wire net3238;
wire net824;
wire net3769;
wire net2639;
wire net1462;
wire net6441;
wire net2736;
wire net3435;
wire net6307;
wire net4696;
wire net831;
wire net3760;
wire net832;
wire net3856;
wire net7368;
wire net9926;
wire net7072;
wire net3702;
wire net2069;
wire in25;
wire net4542;
wire net102;
wire net5349;
wire net841;
wire net1369;
wire net843;
wire net844;
wire net10877;
wire net5536;
wire net2231;
wire net71;
wire net2235;
wire net845;
wire net4330;
wire net7245;
wire net839;
wire net3356;
wire net894;
wire net1068;
wire net6237;
wire net1892;
wire net5882;
wire net1832;
wire net10995;
wire net368;
wire net1159;
wire net7031;
wire net1839;
wire net856;
wire net10097;
wire net3244;
wire net809;
wire net858;
wire net2728;
wire net1449;
wire net1021;
wire net4190;
wire net1736;
wire net860;
wire net972;
wire net10633;
wire net2813;
wire net863;
wire net5712;
wire net4737;
wire net3908;
wire net7967;
wire net2507;
wire net1482;
wire net3471;
wire net2062;
wire net866;
wire net868;
wire net10056;
wire net5279;
wire net2031;
wire net4500;
wire net1507;
wire net5525;
wire net869;
wire net5084;
wire net5399;
wire net6088;
wire net1450;
wire net6799;
wire net871;
wire net1968;
wire net1367;
wire net873;
wire net2698;
wire net5874;
wire net989;
wire net7260;
wire net2458;
wire net6832;
wire net3561;
wire net10119;
wire net4972;
wire net879;
wire net8770;
wire net3852;
wire net9327;
wire net5010;
wire net6861;
wire net3398;
wire net1401;
wire net1083;
wire net10739;
wire net259;
wire net1065;
wire net881;
wire net5335;
wire net2927;
wire net1930;
wire net1973;
wire net6948;
wire net887;
wire net656;
wire net5993;
wire net892;
wire net7872;
wire net4487;
wire net893;
wire net10344;
wire net7326;
wire net6149;
wire net898;
wire net6404;
wire net3266;
wire net6956;
wire net903;
wire net4521;
wire net2889;
wire net5283;
wire net1259;
wire net7798;
wire net3753;
wire net906;
wire net9824;
wire net378;
wire net4111;
wire net955;
wire net6170;
wire net910;
wire net8557;
wire net3432;
wire net1329;
wire net5019;
wire net911;
wire net2697;
wire net4309;
wire net608;
wire net913;
wire net4855;
wire net2447;
wire net714;
wire net922;
wire net3873;
wire net2457;
wire net4973;
wire net2311;
wire net1207;
wire net10050;
wire net926;
wire net5864;
wire net7249;
wire net9365;
wire net616;
wire net1608;
wire net6566;
wire net584;
wire net7314;
wire net930;
wire net2131;
wire net5946;
wire net3089;
wire net5833;
wire net2323;
wire net933;
wire net2593;
wire net4933;
wire net10676;
wire net2294;
wire net4104;
wire net4124;
wire net5741;
wire net1509;
wire net4535;
wire net1298;
wire net936;
wire net788;
wire net3654;
wire net8416;
wire net1955;
wire net6145;
wire net8910;
wire net1339;
wire net4338;
wire net938;
wire net940;
wire net3761;
wire net3813;
wire net7178;
wire net3405;
wire net3979;
wire net8790;
wire net1147;
wire net5633;
wire net9952;
wire net1093;
wire net941;
wire net1737;
wire net943;
wire net4220;
wire net1657;
wire net990;
wire net10765;
wire net7677;
wire net946;
wire net1980;
wire net3189;
wire net1907;
wire net6461;
wire net7896;
wire net1364;
wire net1191;
wire net1136;
wire net6214;
wire net8267;
wire net3093;
wire net948;
wire net614;
wire net5026;
wire net2414;
wire net6419;
wire net1969;
wire net8313;
wire net5403;
wire net1024;
wire net3226;
wire net4409;
wire net8041;
wire net953;
wire net3329;
wire net5784;
wire net954;
wire net2223;
wire net1183;
wire net959;
wire net248;
wire net6128;
wire net7901;
wire net4076;
wire net2609;
wire net5354;
wire net5814;
wire net170;
wire net1194;
wire net391;
wire net1407;
wire net11013;
wire net331;
wire net78;
wire net963;
wire net521;
wire net4931;
wire net5700;
wire net9913;
wire net1027;
wire net11155;
wire net8818;
wire net1816;
wire net1661;
wire net974;
wire net6288;
wire net5583;
wire net2004;
wire net979;
wire net980;
wire out16;
wire net1700;
wire net6723;
wire net4557;
wire net983;
wire net3282;
wire net8506;
wire net815;
wire net991;
wire net203;
wire net2267;
wire net1299;
wire net1928;
wire net6476;
wire net2856;
wire net1776;
wire net1000;
wire net3150;
wire net1003;
wire net466;
wire net2854;
wire net4139;
wire net789;
wire net1005;
wire net1008;
wire net3591;
wire net6654;
wire net2897;
wire net1427;
wire net8229;
wire net3604;
wire net8088;
wire net2662;
wire net1013;
wire net882;
wire net3343;
wire net11075;
wire net3208;
wire net10370;
wire net1629;
wire net416;
wire net4440;
wire net1023;
wire net2537;
wire net498;
wire net4856;
wire net1541;
wire net528;
wire net6203;
wire net1115;
wire net6766;
wire net10987;
wire net10205;
wire net2198;
wire net5411;
wire net1031;
wire net1694;
wire net2799;
wire net11024;
wire net4429;
wire net10982;
wire net1035;
wire net7883;
wire net4482;
wire net5263;
wire net284;
wire net5660;
wire net1510;
wire net29;
wire net4527;
wire net606;
wire net4646;
wire net7957;
wire net1036;
wire net3263;
wire net4394;
wire net1871;
wire net9302;
wire net694;
wire net2770;
wire net1042;
wire net4513;
wire net9744;
wire net7345;
wire net9510;
wire net3703;
wire net567;
wire net1044;
wire net630;
wire net3048;
wire net7793;
wire net5668;
wire net1152;
wire net2895;
wire net5524;
wire net4010;
wire net2316;
wire net1045;
wire net2297;
wire net7637;
wire net1711;
wire net1400;
wire net5167;
wire net4267;
wire net1269;
wire net250;
wire net4990;
wire net2531;
wire net2613;
wire net5519;
wire net1048;
wire net6465;
wire net2755;
wire net1422;
wire net1879;
wire net10432;
wire net8420;
wire net1020;
wire net2492;
wire net1056;
wire net10314;
wire net2501;
wire net4425;
wire net5262;
wire net6697;
wire net6813;
wire net4601;
wire net5538;
wire net2454;
wire net5305;
wire net10434;
wire net602;
wire net1744;
wire net1062;
wire net9229;
wire net3751;
wire net10250;
wire net2614;
wire net1066;
wire net1067;
wire net6671;
wire net1071;
wire net42;
wire net5064;
wire net1072;
wire net4971;
wire net8967;
wire net8211;
wire net2780;
wire net1642;
wire net3231;
wire net9819;
wire net1622;
wire net2055;
wire net10626;
wire net1630;
wire net7563;
wire net1073;
wire net1227;
wire net1076;
wire net1361;
wire net1150;
wire net9551;
wire net5038;
wire net2301;
wire net6455;
wire net11219;
wire net9730;
wire net6267;
wire net1868;
wire net1079;
wire net5272;
wire net2472;
wire net92;
wire net2809;
wire net3886;
wire net1500;
wire net3962;
wire net9643;
wire net6434;
wire net880;
wire net6764;
wire net5410;
wire net739;
wire net1081;
wire net386;
wire net5669;
wire net2757;
wire net1094;
wire net1323;
wire net7223;
wire net142;
wire net2011;
wire net5447;
wire net2612;
wire net389;
wire net7481;
wire net1098;
wire net9150;
wire net1406;
wire net273;
wire net1099;
wire net1493;
wire net1101;
wire net1103;
wire net10568;
wire net9814;
wire net7102;
wire net1105;
wire net3152;
wire net5284;
wire net2405;
wire net6684;
wire net8133;
wire net16;
wire net2206;
wire net2455;
wire net4515;
wire net1108;
wire net3835;
wire net9584;
wire net5229;
wire net1978;
wire net3768;
wire net3069;
wire net1634;
wire net1665;
wire net1039;
wire net9440;
wire net4026;
wire net3072;
wire net5963;
wire net1112;
wire net1119;
wire net314;
wire net1090;
wire net1120;
wire net1523;
wire net4023;
wire net1126;
wire net7192;
wire net3365;
wire net1818;
wire net1127;
wire net1712;
wire net10781;
wire net8440;
wire net1129;
wire net4336;
wire net5415;
wire net5455;
wire net1130;
wire net11138;
wire net1131;
wire net4742;
wire net5210;
wire net3065;
wire net684;
wire net1132;
wire out23;
wire net1589;
wire net7589;
wire net1133;
wire net8340;
wire net3292;
wire net7095;
wire net3054;
wire net2644;
wire net6872;
wire net6225;
wire net2564;
wire net5165;
wire net6980;
wire net619;
wire net1141;
wire net2133;
wire net2594;
wire net4915;
wire net2488;
wire net5394;
wire out15;
wire net1144;
wire net4439;
wire net8767;
wire net1149;
wire net1077;
wire net456;
wire net7137;
wire net10917;
wire net392;
wire net6234;
wire net10560;
wire net1230;
wire net9121;
wire net1652;
wire net1411;
wire net3602;
wire net2121;
wire net8599;
wire net1160;
wire net4060;
wire net2795;
wire net2976;
wire net2937;
wire net9707;
wire net2320;
wire net1161;
wire net6677;
wire net11084;
wire net2715;
wire net2512;
wire net1164;
wire net1303;
wire net7239;
wire net2112;
wire net3499;
wire net1996;
wire net9101;
wire net6324;
wire net62;
wire net1171;
wire net2434;
wire net2540;
wire net5069;
wire net9521;
wire net3075;
wire net1174;
wire net6228;
wire net5421;
wire net201;
wire net9556;
wire net9092;
wire net1906;
wire net3566;
wire net2944;
wire net1180;
wire net5464;
wire net7319;
wire net2920;
wire net2139;
wire net2359;
wire net4908;
wire net3430;
wire net615;
wire net5820;
wire net10952;
wire net460;
wire net6877;
wire net1184;
wire net2867;
wire net2239;
wire net8590;
wire net1799;
wire net1186;
wire net9626;
wire net821;
wire net9792;
wire net2449;
wire net9388;
wire net34;
wire net5867;
wire net9442;
wire net358;
wire net1516;
wire net4110;
wire net6761;
wire net8817;
wire net1281;
wire net3603;
wire net9662;
wire net8310;
wire net76;
wire net3887;
wire net1199;
wire net1268;
wire net1311;
wire net1201;
wire net1202;
wire net10166;
wire net4551;
wire net7702;
wire net4609;
wire net9776;
wire net3424;
wire net8662;
wire net6876;
wire net1206;
wire net3044;
wire net2090;
wire net558;
wire net4671;
wire net668;
wire net3422;
wire net1578;
wire net5838;
wire net1209;
wire net7328;
wire net9218;
wire net226;
wire net7638;
wire net1604;
wire net3138;
wire net1313;
wire net8698;
wire net1217;
wire net2403;
wire net4154;
wire net4313;
wire net120;
wire net2605;
wire net4493;
wire net1267;
wire net5645;
wire net2394;
wire net2099;
wire net1222;
wire net1491;
wire net1225;
wire net6591;
wire net1228;
wire net2369;
wire net2489;
wire net9921;
wire net2046;
wire net883;
wire net5483;
wire net964;
wire net5827;
wire net11101;
wire net1232;
wire net256;
wire net1238;
wire net6636;
wire net2803;
wire net3091;
wire net2376;
wire net8563;
wire net8056;
wire net1240;
wire net8228;
wire net888;
wire net747;
wire net3520;
wire net1244;
wire net9414;
wire net5271;
wire net1718;
wire net5166;
wire net5974;
wire net215;
wire net1245;
wire net3627;
wire net6431;
wire net7465;
wire net11019;
wire net3114;
wire net1248;
wire net2228;
wire net1251;
wire net4849;
wire net2794;
wire net3258;
wire net3104;
wire net1231;
wire net2868;
wire net140;
wire net1255;
wire net8674;
wire net2146;
wire net1162;
wire net3429;
wire net9049;
wire net1257;
wire net2991;
wire net4793;
wire net91;
wire net1990;
wire net67;
wire net401;
wire net5257;
wire net3970;
wire net654;
wire net1276;
wire net1278;
wire net8943;
wire net909;
wire net3960;
wire out21;
wire net4231;
wire net9125;
wire net5037;
wire net6927;
wire net1279;
wire net1598;
wire net6526;
wire net5758;
wire net798;
wire net1280;
wire net5724;
wire net8298;
wire net1307;
wire net7681;
wire net5378;
wire net2885;
wire net468;
wire net6398;
wire net421;
wire net1480;
wire net636;
wire net10227;
wire net3092;
wire net1282;
wire net4068;
wire net11225;
wire net6221;
wire net6692;
wire net1283;
wire net5194;
wire net5400;
wire net9077;
wire net1357;
wire net1286;
wire net1288;
wire net7597;
wire net5774;
wire net11005;
wire net1289;
wire net3551;
wire net1292;
wire net6576;
wire net10627;
wire net2699;
wire net1296;
wire net1550;
wire net1911;
wire net10539;
wire net9062;
wire net4215;
wire net1301;
wire net1302;
wire net7353;
wire net688;
wire net1553;
wire net1471;
wire net4748;
wire net7158;
wire net1306;
wire net1585;
wire net8679;
wire net8184;
wire net4958;
wire net5277;
wire net10516;
wire net1316;
wire net2360;
wire net6774;
wire net440;
wire net7492;
wire net4133;
wire net1831;
wire net1522;
wire net1322;
wire net4230;
wire net2802;
wire net2558;
wire net5630;
wire net1327;
wire net5156;
wire net1398;
wire net3107;
wire net3790;
wire net1619;
wire net9117;
wire net1341;
wire net2406;
wire net1342;
wire net1350;
wire net1300;
wire net2464;
wire net5629;
wire net6148;
wire net1260;
wire net1351;
wire net10875;
wire net4470;
wire net1355;
wire net5887;
wire net1483;
wire net8931;
wire net2958;
wire net4234;
wire net834;
wire net10262;
wire net5790;
wire net1360;
wire net3935;
wire net7463;
wire net2441;
wire net1627;
wire net1562;
wire net10040;
wire net3183;
wire net643;
wire net1319;
wire net7959;
wire net2169;
wire net1366;
wire net5057;
wire net2589;
wire net4462;
wire net952;
wire net3448;
wire net1580;
wire net6796;
wire net351;
wire net4452;
wire net8090;
wire net848;
wire net10723;
wire net7226;
wire net1375;
wire net9872;
wire net3464;
wire net3925;
wire net973;
wire net451;
wire net2734;
wire net7685;
wire net1378;
wire net1092;
wire net6882;
wire net8703;
wire net1380;
wire net7828;
wire net1381;
wire net4387;
wire net10426;
wire net6425;
wire net9614;
wire net1382;
wire net10025;
wire net1389;
wire net2880;
wire net1435;
wire net9829;
wire net2466;
wire net804;
wire net10680;
wire net3607;
wire net937;
wire net1385;
wire net1386;
wire net5539;
wire net1388;
wire net3045;
wire in15;
wire net711;
wire net1591;
wire net1784;
wire net7070;
wire net1391;
wire net2080;
wire net10203;
wire net2548;
wire net719;
wire net3572;
wire net1394;
wire net1395;
wire net2721;
wire net6905;
wire net1962;
wire net1399;
wire net8928;
wire net931;
wire net381;
wire net429;
wire net1402;
wire net7015;
wire net1403;
wire net2213;
wire net2982;
wire net484;
wire net2075;
wire net4768;
wire net1085;
wire net1404;
wire net828;
wire net2450;
wire net1413;
wire net321;
wire net4081;
wire net2883;
wire net7450;
wire net2775;
wire net6337;
wire net8775;
wire net405;
wire net10391;
wire net10069;
wire net7504;
wire net1424;
wire net2423;
wire net1431;
wire net6565;
wire net6264;
wire net1944;
wire net1637;
wire net1432;
wire net2929;
wire net1600;
wire net3386;
wire net1433;
wire net1607;
wire net2250;
wire net1157;
wire net8801;
wire net1438;
wire net1441;
wire net5553;
wire net11134;
wire net9168;
wire net1344;
wire net1453;
wire net7101;
wire net7276;
wire net6472;
wire net697;
wire net4565;
wire net2999;
wire net433;
wire net6864;
wire net1333;
wire net1457;
wire net899;
wire net3537;
wire net1091;
wire net5837;
wire net1454;
wire net10577;
wire net7506;
wire net5360;
wire net1455;
wire net2254;
wire net2641;
wire net1844;
wire net2065;
wire net7475;
wire net3050;
wire net1456;
wire net1458;
wire net2844;
wire net7295;
wire net576;
wire net3043;
wire net10195;
wire net1626;
wire net6971;
wire net2683;
wire net1143;
wire net6038;
wire net6682;
wire net1461;
wire net1579;
wire net3563;
wire net1353;
wire net6229;
wire net1469;
wire net1169;
wire net1084;
wire net7262;
wire net4622;
wire net5027;
wire net5778;
wire net6068;
wire net1470;
wire net3518;
wire net6637;
wire net929;
wire net1473;
wire net447;
wire net1189;
wire net1478;
wire net5009;
wire net7022;
wire net2175;
wire net1271;
wire net5779;
wire net10390;
wire net3154;
wire net1484;
wire net6186;
wire net6975;
wire net7650;
wire net803;
wire net4015;
wire net3144;
wire net3644;
wire net3255;
wire net3019;
wire net1494;
wire net4079;
wire net5062;
wire net1496;
wire net5688;
wire net2966;
wire net9037;
wire net1497;
wire net6114;
wire net7204;
wire net3013;
wire net3181;
wire net1950;
wire net1504;
wire net10191;
wire net8596;
wire net3524;
wire net1670;
wire net4393;
wire net829;
wire net10192;
wire net1506;
wire net6573;
wire net8278;
wire net8268;
wire net14;
wire net8384;
wire net5695;
wire net1512;
wire net10688;
wire net5289;
wire net669;
wire net1513;
wire net10463;
wire net1514;
wire net10003;
wire net3549;
wire net1648;
wire net316;
wire net8481;
wire net1618;
wire net2562;
wire net7338;
wire net1916;
wire net1760;
wire net7418;
wire net8716;
wire net8200;
wire net1524;
wire net11018;
wire net1833;
wire net709;
wire in14;
wire net9981;
wire net3984;
wire net6730;
wire net8866;
wire net2671;
wire net375;
wire net5647;
wire net1485;
wire net1531;
wire net6607;
wire net1533;
wire net10014;
wire net1536;
wire net3490;
wire net10103;
wire net1584;
wire net5549;
wire net1735;
wire net5614;
wire net122;
wire net1547;
wire net9264;
wire net2178;
wire net1798;
wire net5058;
wire net1548;
wire net3954;
wire net7011;
wire net6924;
wire net115;
wire net7457;
wire net1554;
wire net8108;
wire net6645;
wire net778;
wire net557;
wire net190;
wire net5599;
wire net1557;
wire net3479;
wire net1559;
wire net677;
wire net1570;
wire net1746;
wire net837;
wire net3793;
wire net4847;
wire net5776;
wire net7016;
wire net77;
wire net1843;
wire net956;
wire net796;
wire net6973;
wire net7159;
wire net4035;
wire net4374;
wire net1564;
wire net4072;
wire net2882;
wire net7635;
wire net2549;
wire net8748;
wire net1565;
wire net2116;
wire net3988;
wire net125;
wire net1926;
wire net1574;
wire net10774;
wire net1576;
wire net2919;
wire net8064;
wire net4413;
wire net1577;
wire net3283;
wire net1581;
wire net5264;
wire net4039;
wire net1587;
wire net8352;
wire net2087;
wire net1963;
wire net1920;
wire net6989;
wire net1594;
wire net3457;
wire net8204;
wire net7235;
wire net7241;
wire net1285;
wire net1078;
wire net242;
wire net2141;
wire net7082;
wire net9770;
wire net1606;
wire net1924;
wire net7046;
wire net1609;
wire net2523;
wire net308;
wire net2266;
wire net4901;
wire net1167;
wire net2669;
wire net7103;
wire net3805;
wire net2785;
wire net942;
wire net5727;
wire net1572;
wire net7555;
wire net1304;
wire net1620;
wire net257;
wire net1852;
wire net5555;
wire net3415;
wire net9986;
wire net1623;
wire net2355;
wire net1124;
wire net7185;
wire net1697;
wire net3108;
wire net1633;
wire net4148;
wire net8192;
wire net3106;
wire net5579;
wire net5371;
wire net8582;
wire net618;
wire net2690;
wire net1641;
wire net527;
wire net1644;
wire net1646;
wire net1651;
wire net1650;
wire net4710;
wire net2909;
wire net2028;
wire net5440;
wire net4181;
wire net3117;
wire net4620;
wire net1490;
wire net4589;
wire net205;
wire net4058;
wire net4185;
wire net2774;
wire net1479;
wire net6351;
wire net867;
wire net1904;
wire net7945;
wire net1669;
wire net623;
wire net4200;
wire net10653;
wire net10534;
wire net1671;
wire net8289;
wire net2686;
wire net2217;
wire net1672;
wire net3358;
wire net921;
wire net6483;
wire net712;
wire net1674;
wire net2824;
wire net3040;
wire net1682;
wire net108;
wire net3196;
wire net7296;
wire net7963;
wire net3241;
wire net9301;
wire net271;
wire net5242;
wire net5746;
wire net1685;
wire net3041;
wire net3933;
wire net1751;
wire net1703;
wire net1686;
wire net10429;
wire net10159;
wire net782;
wire net1690;
wire net52;
wire net1692;
wire net2092;
wire net6640;
wire net1698;
wire net439;
wire net5000;
wire net5950;
wire net605;
wire out3;
wire net2484;
wire net10331;
wire net3296;
wire net6965;
wire net1706;
wire net6039;
wire net7952;
wire net1709;
wire net692;
wire net6385;
wire net3713;
wire net7979;
wire net3716;
wire net4352;
wire net4398;
wire net1667;
wire net3717;
wire net3259;
wire net3719;
wire net1246;
wire net5799;
wire net3720;
wire net543;
wire net3722;
wire net1599;
wire net3772;
wire net9031;
wire net4657;
wire net1247;
wire net5494;
wire net982;
wire net7423;
wire net4796;
wire net3723;
wire net5843;
wire net3725;
wire net5002;
wire net3727;
wire net3728;
wire net6862;
wire net3730;
wire net10054;
wire net9172;
wire net3731;
wire net5967;
wire net3732;
wire net3734;
wire net10794;
wire net9042;
wire net3735;
wire net2432;
wire net4071;
wire net2127;
wire net3736;
wire net9254;
wire net3739;
wire net8315;
wire net4087;
wire net8813;
wire net5849;
wire net8031;
wire net1866;
wire net5656;
wire net3740;
wire net3741;
wire net9864;
wire net9070;
wire net9009;
wire net1758;
wire net3743;
wire net9827;
wire net3744;
wire net3222;
wire net260;
wire net3748;
wire net7774;
wire net6023;
wire net3749;
wire net4163;
wire net1356;
wire net3754;
wire net3756;
wire net6639;
wire net1616;
wire net7130;
wire net3757;
wire net3758;
wire net3715;
wire net7458;
wire net1187;
wire net3759;
wire net3763;
wire net3764;
wire net8499;
wire net8446;
wire net3766;
wire net10466;
wire net6661;
wire net3767;
wire net3774;
wire net10694;
wire net4178;
wire net3776;
wire net5208;
wire net7120;
wire net5782;
wire net1444;
wire net6655;
wire net3779;
wire net3918;
wire net2336;
wire net3780;
wire net3783;
wire net3786;
wire net8483;
wire net1242;
wire net3787;
wire net3928;
wire net3788;
wire net3789;
wire net3265;
wire net1211;
wire net4874;
wire net6048;
wire net8214;
wire net4014;
wire net6449;
wire net4736;
wire net7576;
wire net3301;
wire net3796;
wire net5173;
wire net4735;
wire net2328;
wire net7142;
wire net3798;
wire net3799;
wire net3800;
wire net3801;
wire net3807;
wire net9977;
wire net6492;
wire net3809;
wire net4665;
wire net1086;
wire net3810;
wire net7347;
wire net3812;
wire net5376;
wire net3814;
wire net6329;
wire net10766;
wire net3433;
wire net3817;
wire net7000;
wire net3818;
wire net3819;
wire net6335;
wire net3820;
wire net3821;
wire net10531;
wire net3822;
wire net8233;
wire net3826;
wire net5092;
wire net3827;
wire net10111;
wire net9762;
wire net4103;
wire net3828;
wire net7766;
wire net3829;
wire net3846;
wire net3830;
wire net6473;
wire net3833;
wire net2907;
wire net6026;
wire net3834;
wire net10659;
wire net3837;
wire net2986;
wire net6387;
wire net3653;
wire net3839;
wire net3840;
wire net3841;
wire net4782;
wire net5613;
wire net3842;
wire net716;
wire net3844;
wire net7817;
wire net3847;
wire net3824;
wire net4951;
wire net2713;
wire net3849;
wire net40;
wire net6172;
wire net3851;
wire net11121;
wire net3853;
wire net3854;
wire net9441;
wire net4408;
wire net3855;
wire net3857;
wire net3861;
wire net3862;
wire net3864;
wire net9531;
wire net3866;
wire net7778;
wire net4510;
wire net3867;
wire net3868;
wire net3869;
wire net9433;
wire net3870;
wire net5140;
wire net3871;
wire net4967;
wire net1195;
wire net6142;
wire net3872;
wire net3874;
wire net5704;
wire net4161;
wire net3437;
wire net3875;
wire net8548;
wire net2922;
wire net1783;
wire net3877;
wire net7940;
wire net3878;
wire net10501;
wire net3879;
wire net3880;
wire net5158;
wire net10057;
wire net7808;
wire net3598;
wire net3882;
wire net1053;
wire net3888;
wire net10682;
wire net3629;
wire net3889;
wire net3891;
wire net3893;
wire net8098;
wire net465;
wire net1860;
wire net3894;
wire net3895;
wire net9297;
wire net8664;
wire net2418;
wire net3902;
wire net7444;
wire net3555;
wire net3903;
wire net3904;
wire net11020;
wire net7987;
wire net3905;
wire net5080;
wire net3906;
wire net9808;
wire net4016;
wire net3907;
wire net5530;
wire net3909;
wire net4811;
wire net8375;
wire net7773;
wire net3910;
wire net3911;
wire net5649;
wire net3912;
wire net3916;
wire net4733;
wire net6124;
wire net5456;
wire net5496;
wire net6298;
wire net6578;
wire net9219;
wire net3917;
wire net7071;
wire net3919;
wire net3272;
wire net3922;
wire net5664;
wire net6731;
wire net3924;
wire net11153;
wire net1354;
wire net3926;
wire net3929;
wire net8804;
wire net3931;
wire net1216;
wire net1750;
wire net1753;
wire net3932;
wire net1532;
wire net6073;
wire net3934;
wire net3936;
wire net5578;
wire net8604;
wire net3937;
wire net9447;
wire net3664;
wire net3938;
wire net3940;
wire net900;
wire net3941;
wire net10112;
wire net1193;
wire net4764;
wire net3943;
wire net3946;
wire net3947;
wire net3948;
wire net3951;
wire net3952;
wire net3953;
wire net3956;
wire net3957;
wire net9477;
wire net3959;
wire net3963;
wire net6043;
wire net3966;
wire net5412;
wire net6787;
wire net3968;
wire net5007;
wire net3971;
wire net419;
wire net3974;
wire net9196;
wire net3975;
wire net4235;
wire net6046;
wire net3978;
wire net1515;
wire net4186;
wire net9345;
wire net5622;
wire net3981;
wire net10536;
wire net3982;
wire net1936;
wire net3985;
wire net3986;
wire net3991;
wire net3992;
wire net7170;
wire net11081;
wire net2282;
wire net3993;
wire net3994;
wire net6120;
wire net3996;
wire net3997;
wire net6358;
wire net3998;
wire net7947;
wire net3706;
wire net4089;
wire net3999;
wire net8089;
wire net2828;
wire net4003;
wire net2490;
wire net6403;
wire net4109;
wire net5126;
wire net4005;
wire net6630;
wire net10695;
wire net4007;
wire net4008;
wire net9754;
wire net8376;
wire net4012;
wire net46;
wire net4018;
wire net6543;
wire net4020;
wire net7435;
wire net4021;
wire net4926;
wire net4022;
wire net5900;
wire net1135;
wire net4024;
wire net11200;
wire net4580;
wire net6072;
wire net11071;
wire net8061;
wire net4027;
wire net6510;
wire net539;
wire net5386;
wire net7047;
wire net4028;
wire net4030;
wire net4031;
wire net4033;
wire net4036;
wire net4037;
wire net4820;
wire net6998;
wire net4038;
wire net4040;
wire net4042;
wire net666;
wire net4043;
wire net4276;
wire net4045;
wire net1917;
wire net5743;
wire net9354;
wire net5164;
wire net994;
wire net4046;
wire net4049;
wire net9549;
wire net8630;
wire net7611;
wire net4051;
wire net4052;
wire net6427;
wire net4053;
wire net4055;
wire net8562;
wire net4057;
wire net4059;
wire net10807;
wire net10788;
wire net8687;
wire net6422;
wire net658;
wire net5503;
wire net4061;
wire net4062;
wire net10777;
wire net5685;
wire net7065;
wire net4064;
wire net4084;
wire net8872;
wire net790;
wire net4065;
wire net6176;
wire net7839;
wire net6634;
wire net4066;
wire net565;
wire net4067;
wire net4069;
wire net8334;
wire net2310;
wire net4070;
wire net6541;
wire net4073;
wire net4680;
wire net6322;
wire net4077;
wire net7664;
wire net907;
wire net150;
wire net4078;
wire net4080;
wire net4082;
wire net9566;
wire net4083;
wire net10581;
wire net8162;
wire net2623;
wire net4090;
wire net5299;
wire net4091;
wire net10106;
wire net9072;
wire net4719;
wire net4093;
wire net5948;
wire net4095;
wire out24;
wire net4728;
wire net4101;
wire net8008;
wire net4434;
wire net5227;
wire net6448;
wire net5991;
wire net6763;
wire net5088;
wire net10674;
wire net4105;
wire net1423;
wire net4106;
wire net10654;
wire net4112;
wire net4114;
wire net7230;
wire net4117;
wire net3724;
wire net4119;
wire net4123;
wire net3425;
wire net5469;
wire net5321;
wire net6866;
wire net2358;
wire net4125;
wire net4126;
wire net4127;
wire net10113;
wire net5769;
wire net4129;
wire net4131;
wire net9562;
wire net4132;
wire net4136;
wire net3038;
wire net4140;
wire net7838;
wire net2465;
wire net4141;
wire net4142;
wire net82;
wire net4144;
wire net8533;
wire net1134;
wire net4145;
wire net4146;
wire net4147;
wire net1235;
wire net5116;
wire net2984;
wire net4150;
wire net8059;
wire net4152;
wire net7951;
wire net2786;
wire net5389;
wire net410;
wire net4155;
wire net449;
wire net7344;
wire net4160;
wire net4164;
wire net3087;
wire net4165;
wire net1142;
wire net4168;
wire net3156;
wire net4169;
wire net1417;
wire net2185;
wire net4171;
wire net5230;
wire net4173;
wire net4177;
wire net2511;
wire net4182;
wire net7831;
wire net6506;
wire net10172;
wire net148;
wire net4183;
wire net4187;
wire net5074;
wire net4189;
wire net6649;
wire net9271;
wire net5071;
wire net4192;
wire net3901;
wire net6993;
wire net4193;
wire net497;
wire net4194;
wire net8116;
wire net6255;
wire net7270;
wire net4197;
wire net2027;
wire net4198;
wire net9998;
wire net4199;
wire net10137;
wire net4265;
wire net8424;
wire net6310;
wire net4203;
wire net4205;
wire net4207;
wire net4208;
wire net1701;
wire net4209;
wire net3564;
wire net5302;
wire net5423;
wire net2768;
wire net4212;
wire net4217;
wire net4221;
wire net3328;
wire net4222;
wire net4648;
wire net235;
wire net5990;
wire net4223;
wire net8094;
wire net4224;
wire net917;
wire net4226;
wire net4227;
wire net10813;
wire net4228;
wire net4232;
wire net11000;
wire net4233;
wire net5207;
wire net3729;
wire net4237;
wire net4240;
wire net4241;
wire net2218;
wire net7189;
wire net11129;
wire net4245;
wire net6204;
wire net9656;
wire net4246;
wire net2965;
wire net5198;
wire net4247;
wire net6125;
wire net4248;
wire net6416;
wire net4249;
wire net4251;
wire net6488;
wire net4253;
wire net8657;
wire net4256;
wire net1628;
wire net4258;
wire net6785;
wire net9950;
wire net4259;
wire net5345;
wire net7104;
wire net4262;
wire net8000;
wire net1439;
wire net4263;
wire net3178;
wire net4269;
wire net1566;
wire net4264;
wire net4268;
wire net5434;
wire net4274;
wire net5135;
wire net3243;
wire net342;
wire net4275;
wire net2624;
wire net4278;
wire net54;
wire net4279;
wire net4281;
wire net11179;
wire net4631;
wire net4283;
wire net9308;
wire net9262;
wire net4284;
wire net4285;
wire net4286;
wire net4588;
wire net4612;
wire net3319;
wire net4288;
wire net2177;
wire net4289;
wire net4291;
wire net4292;
wire net4294;
wire net4295;
wire net4297;
wire net8135;
wire net4298;
wire net11022;
wire net4299;
wire net7079;
wire net4300;
wire net8065;
wire net2587;
wire net4302;
wire net2632;
wire net4826;
wire net1416;
wire net4305;
wire net2024;
wire net5944;
wire net7115;
wire net4311;
wire net6991;
wire net10799;
wire net7608;
wire net4314;
wire net8933;
wire net8019;
wire net4491;
wire net4318;
wire net4325;
wire net4625;
wire net4328;
wire net6252;
wire net4331;
wire net7384;
wire net10960;
wire net10251;
wire net519;
wire net4157;
wire net4332;
wire net4836;
wire net7256;
wire net4333;
wire net4334;
wire net4335;
wire net6361;
wire net8393;
wire net4339;
wire net7390;
wire net10243;
wire net4340;
wire net3335;
wire net4341;
wire net8141;
wire net5502;
wire net4342;
wire net8797;
wire net4188;
wire net4343;
wire net4970;
wire net4344;
wire net4345;
wire net2322;
wire net5401;
wire net2321;
wire net5049;
wire net10478;
wire net9698;
wire net4349;
wire net4350;
wire net5060;
wire net10876;
wire net4351;
wire net7329;
wire net8085;
wire net6504;
wire net4356;
wire net4357;
wire net4358;
wire net2717;
wire net4359;
wire net6894;
wire net5086;
wire net4360;
wire net10554;
wire net7722;
wire net6151;
wire net10462;
wire net4361;
wire net118;
wire net4364;
wire net1121;
wire net4367;
wire net4368;
wire net4369;
wire net4371;
wire net8451;
wire net517;
wire net4375;
wire net7495;
wire net7126;
wire net4376;
wire net6380;
wire net6849;
wire net4377;
wire net1082;
wire net6376;
wire in19;
wire net4379;
wire net4380;
wire net7190;
wire net4381;
wire net7639;
wire net1845;
wire net5429;
wire net4382;
wire net4383;
wire net10881;
wire net302;
wire net1740;
wire net4385;
wire net10217;
wire net4000;
wire net4386;
wire net1762;
wire net1679;
wire net4261;
wire net4388;
wire net7815;
wire net5114;
wire net6629;
wire net4392;
wire net4395;
wire net4396;
wire net10512;
wire net4853;
wire net4397;
wire net5100;
wire net5255;
wire net10562;
wire net8171;
wire net4399;
wire net4403;
wire net10628;
wire net3897;
wire net6299;
wire net2945;
wire in11;
wire net4405;
wire net4410;
wire net10966;
wire net4412;
wire net6539;
wire net4416;
wire net4417;
wire net4418;
wire net4419;
wire net9838;
wire net8285;
wire net6481;
wire net8846;
wire net4421;
wire net2314;
wire net6268;
wire net4423;
wire net4426;
wire net4427;
wire net6436;
wire net4428;
wire net7111;
wire net188;
wire net5529;
wire net4433;
wire net9370;
wire net4436;
wire net10199;
wire net4667;
wire net339;
wire net6821;
wire net4438;
wire net4957;
wire net4442;
wire net369;
wire net2445;
wire net4445;
wire net6758;
wire net4446;
wire net5597;
wire net434;
wire net4448;
wire net4450;
wire net7854;
wire net5388;
wire net6585;
wire net4458;
wire net3482;
wire net4461;
wire net2303;
wire net5589;
wire net1655;
wire net424;
wire net4463;
wire net4464;
wire net7837;
wire net4466;
wire net4467;
wire net4469;
wire net1801;
wire net4471;
wire net10642;
wire net10605;
wire net4293;
wire net2136;
wire net5912;
wire net1254;
wire net4474;
wire net4476;
wire net4477;
wire net1691;
wire net4478;
wire net4479;
wire net5021;
wire net4481;
wire net5498;
wire net4484;
wire net7430;
wire net4485;
wire net4486;
wire net4490;
wire net5377;
wire net8237;
wire net4492;
wire net6179;
wire net4494;
wire net4496;
wire net173;
wire net4501;
wire net4503;
wire net4637;
wire net3594;
wire net4504;
wire net7382;
wire net4505;
wire net10346;
wire net675;
wire net4506;
wire net5381;
wire net4508;
wire net2551;
wire net5625;
wire net622;
wire net4509;
wire net2947;
wire net4511;
wire net6366;
wire net5926;
wire net4516;
wire net7599;
wire net4522;
wire net4523;
wire net4524;
wire net4525;
wire net8173;
wire net8115;
wire net4526;
wire net2153;
wire net4530;
wire net2306;
wire net4531;
wire net4534;
wire net11167;
wire net268;
wire net1534;
wire net5428;
wire net4536;
wire net5347;
wire net4539;
wire net5573;
wire net1487;
wire net4540;
wire net4541;
wire net4543;
wire net5420;
wire net469;
wire net4546;
wire net10702;
wire net6560;
wire net4722;
wire net7023;
wire net7332;
wire net4547;
wire net4549;
wire net4550;
wire net4552;
wire net4554;
wire net435;
wire net4555;
wire net5711;
wire net7081;
wire net9599;
wire net4556;
wire net4558;
wire net10077;
wire net508;
wire net4559;
wire net4562;
wire net187;
wire net6668;
wire net4567;
wire net7330;
wire net4569;
wire net6642;
wire net2835;
wire net3206;
wire net4571;
wire net4287;
wire net4572;
wire net4590;
wire net4574;
wire net4575;
wire net10939;
wire net7741;
wire net3373;
wire net4576;
wire net4578;
wire net2095;
wire net6916;
wire net1358;
wire net7321;
wire net4581;
wire net5319;
wire net4583;
wire net6245;
wire net9944;
wire net4585;
wire net3823;
wire net4659;
wire net1590;
wire net4587;
wire net3580;
wire net4592;
wire net5728;
wire net1476;
wire net4593;
wire net4594;
wire net4596;
wire net7735;
wire net6534;
wire net4597;
wire net4598;
wire net7356;
wire net4599;
wire net3976;
wire net4600;
wire net4602;
wire net7048;
wire net4604;
wire net11052;
wire net5322;
wire net6669;
wire net9886;
wire net2676;
wire net4606;
wire net404;
wire out1;
wire net6958;
wire net30;
wire net4611;
wire net4731;
wire net1890;
wire net4613;
wire net6370;
wire net3781;
wire net4614;
wire net4615;
wire net3709;
wire net4616;
wire net4617;
wire net6732;
wire net10542;
wire net4621;
wire net4626;
wire in0;
wire net6919;
wire net3151;
wire net4627;
wire net6001;
wire net2926;
wire net3777;
wire net6932;
wire net3671;
wire net4628;
wire net1363;
wire net4629;
wire net3645;
wire net4630;
wire net4632;
wire net6084;
wire net4634;
wire net4635;
wire net2417;
wire net4050;
wire net4638;
wire net8045;
wire net4838;
wire net4640;
wire net6930;
wire net4641;
wire net4643;
wire net5043;
wire net1808;
wire net6949;
wire net8586;
wire net6572;
wire net4651;
wire net4654;
wire net4655;
wire net9372;
wire net7964;
wire net4656;
wire net5752;
wire net4660;
wire net8182;
wire net4752;
wire net4661;
wire net7419;
wire net4662;
wire net8181;
wire net4663;
wire net4664;
wire net4669;
wire net6152;
wire net4670;
wire net8072;
wire net222;
wire net4672;
wire net4674;
wire net2797;
wire net4675;
wire net4676;
wire net1915;
wire net4677;
wire net4678;
wire net4679;
wire net1274;
wire net4682;
wire net2288;
wire net4686;
wire net4687;
wire net8676;
wire net4688;
wire net4690;
wire net4691;
wire net4755;
wire net8709;
wire net2990;
wire net4693;
wire net4694;
wire net9348;
wire net3700;
wire net4644;
wire net4695;
wire net9468;
wire net4697;
wire net4698;
wire net9340;
wire net4699;
wire net4701;
wire net7827;
wire net4702;
wire net4703;
wire net7273;
wire net6987;
wire net4705;
wire net992;
wire net4707;
wire net8500;
wire net4711;
wire net4366;
wire net5355;
wire net4712;
wire net4713;
wire net6320;
wire net4714;
wire net1088;
wire net218;
wire net4715;
wire net4257;
wire net4716;
wire net4717;
wire net3264;
wire net5742;
wire net4720;
wire net8807;
wire net2751;
wire net4999;
wire net4721;
wire net7720;
wire net4048;
wire net6839;
wire net5161;
wire net4723;
wire net4724;
wire net4725;
wire net4726;
wire net4727;
wire net7676;
wire net4729;
wire net4730;
wire net3990;
wire net6978;
wire net4732;
wire net4734;
wire net7237;
wire net4739;
wire net4740;
wire net4743;
wire net1933;
wire net2850;
wire net4102;
wire net4744;
wire net4746;
wire net4882;
wire net4166;
wire net4749;
wire net4751;
wire net2998;
wire net4753;
wire net4758;
wire net6067;
wire net4835;
wire net4760;
wire net2606;
wire net4761;
wire net4355;
wire net6393;
wire net4762;
wire net9964;
wire net4765;
wire net10805;
wire net9198;
wire net5598;
wire net4767;
wire net1117;
wire net4769;
wire net743;
wire net4770;
wire net6936;
wire net5190;
wire net4771;
wire net4772;
wire net4404;
wire net4432;
wire net6470;
wire net4009;
wire net4776;
wire net4777;
wire net10029;
wire net7995;
wire net7094;
wire net7718;
wire net4778;
wire net4271;
wire net6410;
wire net1106;
wire net4780;
wire net9627;
wire net4783;
wire net4784;
wire net4785;
wire net4430;
wire net4786;
wire net4788;
wire net4791;
wire net4792;
wire net2366;
wire net1543;
wire net4795;
wire net4797;
wire net289;
wire net4800;
wire net2808;
wire net4801;
wire net4805;
wire net4324;
wire net7028;
wire net4806;
wire net4807;
wire net2771;
wire net6437;
wire net740;
wire net4809;
wire net6482;
wire net10354;
wire net470;
wire net4810;
wire net4814;
wire net4816;
wire net4822;
wire net5564;
wire net4823;
wire net10849;
wire net4824;
wire net4519;
wire net4825;
wire net4827;
wire net4829;
wire net6016;
wire net4830;
wire net9223;
wire net6438;
wire net4831;
wire net2367;
wire net4834;
wire net6417;
wire net4837;
wire net10115;
wire net4845;
wire net5287;
wire net3161;
wire net5986;
wire net6432;
wire net3690;
wire net4214;
wire net4848;
wire net4850;
wire net4851;
wire net4548;
wire net5384;
wire net8847;
wire net4857;
wire net4858;
wire net4860;
wire net4861;
wire net4862;
wire net1517;
wire net4864;
wire net4865;
wire net4867;
wire net509;
wire net4870;
wire net4871;
wire net8415;
wire net4872;
wire net1521;
wire net5129;
wire net9540;
wire net1932;
wire net4817;
wire net4875;
wire net5182;
wire net6699;
wire net4876;
wire net10157;
wire net4877;
wire net4879;
wire net4880;
wire net9920;
wire net4883;
wire net720;
wire net4885;
wire net10708;
wire net4886;
wire net4887;
wire net9532;
wire net4888;
wire net7461;
wire net4889;
wire net7941;
wire net4891;
wire net8333;
wire net4892;
wire net9201;
wire net5730;
wire net6059;
wire net8431;
wire net4894;
wire net4895;
wire net4897;
wire net4092;
wire net4898;
wire net6345;
wire net4900;
wire net2433;
wire net4903;
wire net3205;
wire net4905;
wire net4906;
wire net5635;
wire net4909;
wire net10890;
wire net6191;
wire net1675;
wire net5118;
wire net5154;
wire net6915;
wire net4912;
wire net7060;
wire net4914;
wire net7388;
wire net4916;
wire net184;
wire net4918;
wire net6687;
wire net4919;
wire net7888;
wire net4277;
wire net5485;
wire net9939;
wire net9359;
wire net7512;
wire net4920;
wire net5176;
wire net4921;
wire net9242;
wire net4923;
wire net4925;
wire net4928;
wire net8160;
wire net5847;
wire net10977;
wire net6242;
wire net4929;
wire net2194;
wire net4932;
wire net5937;
wire net2341;
wire net4934;
wire net6550;
wire net7578;
wire net4935;
wire net4518;
wire net4936;
wire net4938;
wire net4940;
wire net8324;
wire net4941;
wire net2615;
wire net6917;
wire net4942;
wire net4943;
wire net5581;
wire net7210;
wire net4946;
wire net2961;
wire net745;
wire net4149;
wire net6738;
wire net4947;
wire net4950;
wire net4952;
wire net5111;
wire net4953;
wire net4954;
wire net299;
wire net4956;
wire net6887;
wire net4963;
wire net10790;
wire net10450;
wire net4965;
wire net9849;
wire net6681;
wire net7099;
wire net10093;
wire net7312;
wire net4794;
wire net5444;
wire net1325;
wire net4966;
wire net353;
wire net4968;
wire net5995;
wire net4969;
wire net4974;
wire net4977;
wire net683;
wire net7247;
wire net4980;
wire net5342;
wire net4981;
wire net2281;
wire net4982;
wire net6658;
wire net6674;
wire net4983;
wire net4985;
wire net875;
wire net4986;
wire net4989;
wire net6933;
wire net5282;
wire net6486;
wire net11139;
wire net4992;
wire net8936;
wire net4994;
wire net647;
wire net7043;
wire net4995;
wire net4997;
wire net6323;
wire net8163;
wire net6300;
wire net4115;
wire net5001;
wire net7886;
wire net5606;
wire net3018;
wire net5003;
wire net6426;
wire net2744;
wire net5006;
wire net9319;
wire net5008;
wire net5011;
wire net4013;
wire net5012;
wire net5014;
wire net4242;
wire net5015;
wire net10352;
wire net4902;
wire net5018;
wire net8566;
wire net5239;
wire net420;
wire net6304;
wire net7293;
wire net41;
wire net5020;
wire net6804;
wire net5023;
wire net3357;
wire net3674;
wire net5028;
wire net10038;
wire net2179;
wire net5029;
wire net9736;
wire net9706;
wire net5032;
wire net5033;
wire net5034;
wire net1539;
wire net5035;
wire net5039;
wire net5041;
wire net303;
wire net6180;
wire net5045;
wire net5046;
wire net5047;
wire net5050;
wire net5051;
wire net10940;
wire net5056;
wire net4561;
wire net5063;
wire net7263;
wire net6409;
wire net8351;
wire net6540;
wire net3930;
wire net3792;
wire net7433;
wire net5226;
wire net6981;
wire net5073;
wire net5076;
wire net10502;
wire net5078;
wire net5807;
wire net6163;
wire net5079;
wire net5082;
wire net5083;
wire net7736;
wire net5793;
wire net5085;
wire net5089;
wire net9895;
wire net5094;
wire net6646;
wire net5096;
wire net7460;
wire net950;
wire net5101;
wire net5545;
wire net2598;
wire net4201;
wire net5104;
wire net5107;
wire net5109;
wire net8622;
wire net8581;
wire net5113;
wire net5234;
wire net7432;
wire net7747;
wire net548;
wire net5115;
wire net4029;
wire net5233;
wire net5120;
wire net1810;
wire net5121;
wire net5122;
wire net3287;
wire net5124;
wire net5125;
wire net7689;
wire net5127;
wire net5128;
wire net10013;
wire net6132;
wire net7279;
wire net580;
wire net5130;
wire net9837;
wire net5133;
wire net5134;
wire net10133;
wire net5136;
wire net5137;
wire net6913;
wire net1605;
wire net5138;
wire net3677;
wire net5139;
wire net1612;
wire net5141;
wire net39;
wire net5142;
wire net9498;
wire net5103;
wire net5143;
wire net5144;
wire net5145;
wire net7073;
wire net4195;
wire net5146;
wire net5149;
wire net6961;
wire net9329;
wire net820;
wire net5150;
wire net5151;
wire net5155;
wire net5160;
wire net5162;
wire net9817;
wire net2273;
wire net5163;
wire net5296;
wire net6698;
wire net5168;
wire net9539;
wire net5169;
wire net7844;
wire net814;
wire net5707;
wire net11224;
wire net5170;
wire net5171;
wire net5174;
wire net5175;
wire net6844;
wire net6081;
wire net1111;
wire net5179;
wire net10139;
wire net5181;
wire net5185;
wire net5188;
wire net8154;
wire net5189;
wire net5196;
wire net8401;
wire net5197;
wire net8955;
wire net8670;
wire net5201;
wire net6759;
wire net5203;
wire net5204;
wire net2130;
wire net5205;
wire net5206;
wire net1166;
wire net5209;
wire net2910;
wire net6890;
wire net5212;
wire net7976;
wire net6292;
wire net5213;
wire net5219;
wire net5223;
wire net9945;
wire net6112;
wire net206;
wire net2812;
wire net363;
wire net5228;
wire net2483;
wire net6875;
wire net3136;
wire net5232;
wire net5907;
wire net7206;
wire net2467;
wire net5237;
wire net5240;
wire net6362;
wire net4959;
wire net6119;
wire net1779;
wire net5241;
wire net253;
wire net5244;
wire net5246;
wire net5249;
wire net9189;
wire net5251;
wire net1966;
wire net5252;
wire net7037;
wire net5254;
wire net4424;
wire net5256;
wire net5259;
wire net3353;
wire net4308;
wire net5260;
wire net7398;
wire net5266;
wire net11218;
wire net10298;
wire net5270;
wire net5273;
wire net7288;
wire net6106;
wire net5275;
wire net6333;
wire net4595;
wire net5276;
wire net5280;
wire net8294;
wire net5281;
wire net5286;
wire net2837;
wire net5994;
wire net5290;
wire net1445;
wire net6386;
wire net1038;
wire net5291;
wire net6525;
wire net6164;
wire net5297;
wire net5298;
wire net8515;
wire net4473;
wire net5068;
wire net5300;
wire net5301;
wire net10949;
wire net10213;
wire net5304;
wire net5830;
wire net5307;
wire net4878;
wire net5310;
wire net5311;
wire net2300;
wire net3794;
wire net7265;
wire net9400;
wire net5314;
wire net6536;
wire net5317;
wire net3123;
wire net5320;
wire net1979;
wire net6193;
wire net5323;
wire net3825;
wire net5324;
wire net6901;
wire net5325;
wire net5327;
wire net9094;
wire net3025;
wire net5813;
wire net5328;
wire net5331;
wire net9996;
wire net5333;
wire net5835;
wire net5334;
wire net9719;
wire net355;
wire net5336;
wire net5337;
wire net8999;
wire net8879;
wire net5338;
wire net5339;
wire net1815;
wire net5340;
wire net5627;
wire net5224;
wire net7195;
wire net5557;
wire net5773;
wire net5352;
wire net10616;
wire net4502;
wire net5353;
wire net5356;
wire net2196;
wire net6211;
wire net5357;
wire net10427;
wire net4100;
wire net5717;
wire net6232;
wire net9572;
wire net5359;
wire net5615;
wire net5361;
wire net5364;
wire net10776;
wire net8435;
wire net531;
wire net1764;
wire net5365;
wire net6631;
wire net5366;
wire net5370;
wire net7203;
wire net5374;
wire net5383;
wire net5385;
wire net5390;
wire net5391;
wire net6659;
wire net5393;
wire net5395;
wire net5398;
wire net4704;
wire net5402;
wire net5404;
wire net1535;
wire net5405;
wire net5408;
wire net5413;
wire net5416;
wire net10706;
wire net5417;
wire net5418;
wire net1015;
wire net5419;
wire net26;
wire net5424;
wire net10402;
wire net5425;
wire net5426;
wire net5433;
wire net681;
wire net5435;
wire net5437;
wire net5439;
wire net10484;
wire net5775;
wire net5441;
wire net5442;
wire net10284;
wire net5445;
wire net9527;
wire net5448;
wire net5450;
wire net2925;
wire net5451;
wire net4976;
wire net5452;
wire net7283;
wire net5453;
wire net6626;
wire net104;
wire net5454;
wire net4472;
wire net5459;
wire net6216;
wire net6463;
wire net5461;
wire net5072;
wire net5462;
wire net5466;
wire net5467;
wire net5468;
wire net8491;
wire net7445;
wire net319;
wire net5535;
wire net5470;
wire net5471;
wire net6212;
wire net5472;
wire net5475;
wire net5476;
wire net5477;
wire net7316;
wire net5478;
wire net6867;
wire net6295;
wire net1049;
wire net5479;
wire net5486;
wire net5487;
wire net3020;
wire net850;
wire net1505;
wire net5489;
wire net5490;
wire net5491;
wire net9169;
wire net6140;
wire net5495;
wire out25;
wire net7649;
wire net5677;
wire net5500;
wire net5501;
wire net6617;
wire net5505;
wire net10668;
wire net5506;
wire net9867;
wire net1156;
wire net5509;
wire net9728;
wire net5618;
wire net6800;
wire net10004;
wire net5510;
wire net5511;
wire net10974;
wire net5513;
wire net1972;
wire net5514;
wire net9230;
wire net9179;
wire net5920;
wire net5515;
wire net5516;
wire net5517;
wire net1719;
wire net5522;
wire net2462;
wire net2059;
wire net1873;
wire net5523;
wire net5526;
wire net5527;
wire net5528;
wire net7464;
wire net5531;
wire net3896;
wire net7289;
wire net5532;
wire net6032;
wire net6407;
wire net2181;
wire net5534;
wire net5537;
wire net352;
wire net5540;
wire net4624;
wire net5541;
wire net5542;
wire net5543;
wire net5544;
wire net5547;
wire net5550;
wire net5551;
wire net3942;
wire net5552;
wire net5562;
wire net1312;
wire net5565;
wire net5566;
wire net5567;
wire net5809;
wire net7336;
wire net5942;
wire net7438;
wire net5571;
wire net11030;
wire net111;
wire net5574;
wire net947;
wire net5575;
wire net5157;
wire net5295;
wire net5580;
wire net4210;
wire net5584;
wire net10477;
wire net5585;
wire net4779;
wire net6071;
wire net5587;
wire net5591;
wire net6742;
wire net5592;
wire net5593;
wire net9897;
wire net5595;
wire net1309;
wire net5596;
wire net10021;
wire net7835;
wire net1869;
wire net5600;
wire net5106;
wire net5504;
wire net5601;
wire net6230;
wire net5604;
wire net5605;
wire net7090;
wire net9476;
wire net5608;
wire net3506;
wire net562;
wire net267;
wire net1324;
wire net5611;
wire net4435;
wire net5616;
wire net7620;
wire net5619;
wire net3456;
wire net5620;
wire net5059;
wire net5623;
wire net5631;
wire net5636;
wire net11037;
wire net5640;
wire net2168;
wire net1699;
wire net5641;
wire net7829;
wire net2843;
wire net119;
wire net5642;
wire net568;
wire net5643;
wire net9163;
wire net918;
wire net5644;
wire net5646;
wire net1824;
wire net3261;
wire net5650;
wire net8443;
wire net5651;
wire net5652;
wire net6884;
wire net5653;
wire net5654;
wire net5655;
wire net5657;
wire net6440;
wire net5658;
wire net8559;
wire net2166;
wire net5659;
wire net5662;
wire net10888;
wire net6037;
wire net4365;
wire net7001;
wire net4642;
wire net5663;
wire net5665;
wire net7455;
wire net5666;
wire net5671;
wire net7532;
wire net5052;
wire net5672;
wire net32;
wire net5676;
wire net769;
wire net5679;
wire net10366;
wire net3497;
wire net3404;
wire net5684;
wire net5687;
wire net5770;
wire net5691;
wire net6623;
wire net3659;
wire net5693;
wire net5694;
wire net8848;
wire net4913;
wire net5698;
wire net6213;
wire net5804;
wire net5215;
wire net6653;
wire net5703;
wire net1872;
wire net5705;
wire net9559;
wire net2373;
wire net7174;
wire net7807;
wire net865;
wire net5706;
wire net5708;
wire net2443;
wire net5710;
wire net6819;
wire net266;
wire net5713;
wire net5714;
wire net4480;
wire net4991;
wire net5715;
wire net5716;
wire net8250;
wire net3804;
wire net6169;
wire net5718;
wire net5720;
wire net232;
wire net5721;
wire net5722;
wire net5723;
wire net5725;
wire net5726;
wire net6183;
wire net5729;
wire net9307;
wire net6842;
wire net5731;
wire net5632;
wire net5903;
wire net1128;
wire net4544;
wire net6564;
wire net5732;
wire net7348;
wire net5734;
wire net9135;
wire net5736;
wire net5737;
wire net5738;
wire net5740;
wire net8540;
wire net4623;
wire net5744;
wire net5747;
wire net6686;
wire net9334;
wire net7057;
wire net3313;
wire net5750;
wire net5751;
wire net5754;
wire net3256;
wire net5755;
wire net5757;
wire net590;
wire net5760;
wire net5761;
wire net8373;
wire net7557;
wire net5316;
wire net5762;
wire net6834;
wire net11149;
wire net9846;
wire net5763;
wire net2607;
wire net7272;
wire net3483;
wire net2635;
wire net1995;
wire net5766;
wire net6253;
wire net5772;
wire net5777;
wire net8800;
wire net5781;
wire net7323;
wire net5783;
wire net6845;
wire net7187;
wire net5785;
wire net7885;
wire net2013;
wire net5786;
wire net4420;
wire net5787;
wire net5788;
wire net7819;
wire net5791;
wire net5796;
wire net5797;
wire net2898;
wire net5798;
wire net5915;
wire net5802;
wire net7739;
wire net5054;
wire net6790;
wire net1154;
wire net5803;
wire net5810;
wire net2860;
wire net5811;
wire net708;
wire net2739;
wire net5739;
wire net6413;
wire net10163;
wire net5812;
wire net5817;
wire net6049;
wire net5818;
wire net5819;
wire net9794;
wire net7284;
wire net2319;
wire net5821;
wire net7025;
wire net1474;
wire net5822;
wire net8561;
wire net2748;
wire net5824;
wire net5825;
wire net5826;
wire net5828;
wire net2286;
wire net5831;
wire net2862;
wire net5004;
wire net5832;
wire net5836;
wire net6822;
wire net5840;
wire net156;
wire net5842;
wire net1662;
wire net6516;
wire net5844;
wire net5805;
wire net6977;
wire net5846;
wire net3477;
wire net5850;
wire net2420;
wire net5851;
wire net764;
wire net5852;
wire net7400;
wire net10481;
wire net3223;
wire net5854;
wire net5855;
wire net4706;
wire net5856;
wire net7117;
wire net5857;
wire net5859;
wire net10737;
wire net5860;
wire net6155;
wire net5861;
wire net5274;
wire net5862;
wire net5865;
wire net5870;
wire net5871;
wire net5872;
wire net5873;
wire net4322;
wire net5875;
wire net6695;
wire net124;
wire net4890;
wire net5880;
wire net1787;
wire net5888;
wire net8053;
wire net5153;
wire net7024;
wire net9811;
wire net1953;
wire net7454;
wire net10584;
wire net5894;
wire net6812;
wire net5895;
wire net1880;
wire net5896;
wire net5897;
wire net1058;
wire net5898;
wire net8476;
wire net5853;
wire net5899;
wire net1377;
wire net5901;
wire net5902;
wire net3765;
wire net5904;
wire net8522;
wire net5905;
wire net5909;
wire net4873;
wire net5910;
wire net400;
wire net5911;
wire net5916;
wire net1847;
wire net5917;
wire net5918;
wire net5919;
wire net5921;
wire net5922;
wire net8697;
wire net7118;
wire net5923;
wire net5927;
wire net10964;
wire net10657;
wire net6279;
wire net5929;
wire net2017;
wire net5931;
wire net5932;
wire net9834;
wire net5934;
wire net3708;
wire net5935;
wire net2901;
wire net6693;
wire net5938;
wire net9697;
wire net5939;
wire net5414;
wire net305;
wire net5940;
wire net11043;
wire net5945;
wire net7093;
wire net5949;
wire net7602;
wire net5261;
wire net5951;
wire net7389;
wire net9078;
wire net840;
wire net5954;
wire net5753;
wire net5955;
wire net6371;
wire net5956;
wire net1649;
wire net1464;
wire net5957;
wire net5958;
wire net7978;
wire net2590;
wire net5959;
wire net8883;
wire net5960;
wire net9140;
wire net3540;
wire net6471;
wire net10397;
wire net5962;
wire net1123;
wire net5964;
wire net6928;
wire net10110;
wire net1919;
wire net5969;
wire net9120;
wire net6865;
wire net5970;
wire out13;
wire net6189;
wire net9542;
wire net5971;
wire net5972;
wire net5973;
wire net2582;
wire net5975;
wire net2957;
wire net3816;
wire net5978;
wire net5979;
wire net2912;
wire net5981;
wire net6988;
wire net5982;
wire net754;
wire net5983;
wire net5985;
wire net5988;
wire net5992;
wire net9902;
wire net9815;
wire net2183;
wire net6556;
wire net5996;
wire net3213;
wire net6996;
wire net5998;
wire net6000;
wire net6005;
wire net6007;
wire net7421;
wire net2044;
wire net1752;
wire net1949;
wire net6008;
wire net6009;
wire net2470;
wire net6010;
wire net10449;
wire net6011;
wire net2851;
wire net6012;
wire net6013;
wire net10655;
wire net6014;
wire net1229;
wire net6015;
wire net6018;
wire net2905;
wire net1392;
wire net6020;
wire net6021;
wire net8517;
wire net1825;
wire net6022;
wire net6029;
wire net6030;
wire net6031;
wire net10045;
wire net6290;
wire net5269;
wire net6033;
wire net6034;
wire net8402;
wire net6040;
wire net6041;
wire net9670;
wire net2496;
wire net2052;
wire net6042;
wire net6045;
wire net6047;
wire net6050;
wire net3334;
wire net6051;
wire net6052;
wire net6053;
wire net2611;
wire net4158;
wire net6054;
wire net1061;
wire net6055;
wire net6056;
wire net9458;
wire net6060;
wire net4488;
wire net6061;
wire net11097;
wire net4603;
wire net6457;
wire net6512;
wire net5380;
wire net7123;
wire net5329;
wire net6062;
wire net6065;
wire net6066;
wire net6074;
wire net6075;
wire net228;
wire net5178;
wire net6076;
wire net10062;
wire net6078;
wire net6080;
wire net6082;
wire net6083;
wire net11089;
wire net6085;
wire net6086;
wire net6143;
wire net2619;
wire net2190;
wire net6087;
wire net6090;
wire net3636;
wire net6091;
wire net4056;
wire net6093;
wire net7175;
wire net431;
wire net6098;
wire net3271;
wire net5231;
wire net6100;
wire net7826;
wire net6101;
wire net1294;
wire net6102;
wire net5409;
wire net6628;
wire net8302;
wire net1527;
wire net6158;
wire net6103;
wire net3051;
wire net6104;
wire net1041;
wire net5250;
wire net6105;
wire net7386;
wire net6108;
wire net6109;
wire net4804;
wire net6110;
wire net1263;
wire net1397;
wire net6111;
wire net6113;
wire net6399;
wire net6117;
wire net1349;
wire net6118;
wire net1352;
wire net6121;
wire net6126;
wire net6127;
wire net6129;
wire net1273;
wire net6130;
wire net1561;
wire net6133;
wire net6134;
wire net6135;
wire net4537;
wire net7213;
wire net6136;
wire net6137;
wire net6138;
wire net6139;
wire net6141;
wire net8176;
wire net6144;
wire net6146;
wire net1070;
wire net6888;
wire net10090;
wire net6154;
wire net7097;
wire net8309;
wire net6162;
wire net6902;
wire net6165;
wire net6167;
wire net7191;
wire net11060;
wire net7981;
wire net6289;
wire net6168;
wire net6171;
wire net7299;
wire net7893;
wire net6174;
wire net7903;
wire net7443;
wire net6175;
wire net8258;
wire net6177;
wire net10537;
wire net5110;
wire net6181;
wire net6173;
wire net6182;
wire net10233;
wire net6184;
wire net6185;
wire net10035;
wire net6187;
wire net5474;
wire net1902;
wire net1540;
wire net6190;
wire net2342;
wire net6195;
wire net6196;
wire net9206;
wire net6602;
wire net1715;
wire net6199;
wire net6200;
wire net10457;
wire net6201;
wire net6206;
wire net6208;
wire net9047;
wire net6004;
wire net6209;
wire net7757;
wire net4854;
wire net6210;
wire net6215;
wire net2109;
wire net6217;
wire net3514;
wire net6219;
wire net6220;
wire net11136;
wire net6222;
wire net3412;
wire net341;
wire net6223;
wire net6224;
wire net6227;
wire net4134;
wire net6231;
wire net6233;
wire net5016;
wire net6235;
wire net2546;
wire net6259;
wire net6236;
wire net9590;
wire net1728;
wire net6811;
wire net6238;
wire net7682;
wire net6239;
wire net6241;
wire net6243;
wire net6244;
wire net9123;
wire net1537;
wire net5667;
wire net5570;
wire net6246;
wire net7003;
wire net2035;
wire net1529;
wire net6247;
wire net6250;
wire net2158;
wire net6392;
wire net8147;
wire net6254;
wire net6257;
wire net6258;
wire net9888;
wire net5686;
wire net4911;
wire net6260;
wire net6261;
wire net9954;
wire net6262;
wire net8647;
wire net8601;
wire net1345;
wire net6263;
wire net4459;
wire net136;
wire net6265;
wire net4718;
wire net6266;
wire net8307;
wire net6269;
wire net6270;
wire net6271;
wire net6273;
wire net6274;
wire net6276;
wire net9048;
wire net6282;
wire net7846;
wire net6283;
wire net6571;
wire net6284;
wire net6285;
wire net6286;
wire net6899;
wire net6287;
wire net6291;
wire net8783;
wire net1647;
wire net6293;
wire net1807;
wire net6294;
wire net2395;
wire net1891;
wire net6301;
wire net6305;
wire net3012;
wire net6306;
wire net2124;
wire net6918;
wire net6308;
wire net1957;
wire net1096;
wire net2225;
wire net4088;
wire net6309;
wire net2762;
wire net6313;
wire net6314;
wire net9716;
wire net6406;
wire net8349;
wire net6096;
wire net6315;
wire net6317;
wire net6318;
wire net8291;
wire net6319;
wire net6321;
wire net9321;
wire net6325;
wire net2711;
wire net6326;
wire net6327;
wire net8037;
wire net595;
wire net6328;
wire net7125;
wire net6330;
wire net10128;
wire net5081;
wire net6331;
wire net6334;
wire net8180;
wire net6336;
wire net9243;
wire net6338;
wire net4307;
wire net6339;
wire net6341;
wire net8078;
wire net6468;
wire net6342;
wire net6343;
wire net6346;
wire net3583;
wire net2553;
wire net1107;
wire net6347;
wire net6348;
wire net6349;
wire net6352;
wire net6355;
wire net6359;
wire net10443;
wire net6374;
wire net6505;
wire net6364;
wire net7154;
wire net6365;
wire net9413;
wire net427;
wire net6367;
wire net8036;
wire net6369;
wire net11180;
wire net8792;
wire net6372;
wire net6375;
wire net6377;
wire net6378;
wire net2051;
wire net6379;
wire net9460;
wire net6382;
wire net6383;
wire net10495;
wire net6384;
wire net6388;
wire net6389;
wire net169;
wire net6391;
wire net10058;
wire net6394;
wire net3131;
wire net6396;
wire net6739;
wire net8224;
wire net6397;
wire net6401;
wire net6402;
wire net6405;
wire net8962;
wire net6408;
wire net6491;
wire net6411;
wire net6753;
wire net6412;
wire net8886;
wire net1004;
wire net6415;
wire net6784;
wire net11029;
wire net1047;
wire net6418;
wire net11096;
wire net9655;
wire net6420;
wire net7667;
wire net2685;
wire net6903;
wire net6424;
wire net6428;
wire net7002;
wire net687;
wire net1412;
wire net7179;
wire net3742;
wire net6430;
wire net4121;
wire net6433;
wire net3472;
wire net6439;
wire net4270;
wire net6443;
wire net6444;
wire net6445;
wire net9681;
wire net6446;
wire net8246;
wire net5878;
wire net6447;
wire net3750;
wire net4391;
wire net6452;
wire net6453;
wire net6454;
wire net7039;
wire net6456;
wire net6459;
wire net6460;
wire net3385;
wire net6469;
wire net6475;
wire net1898;
wire net6477;
wire net6478;
wire net6479;
wire net1546;
wire net6480;
wire net7717;
wire net7161;
wire net4639;
wire net6487;
wire net6489;
wire net6493;
wire net1140;
wire net6494;
wire net6497;
wire net9471;
wire net6499;
wire net6501;
wire net5431;
wire net6503;
wire net5863;
wire net6535;
wire net6603;
wire net6507;
wire net6508;
wire net5733;
wire net7480;
wire net7542;
wire net6511;
wire net10589;
wire net10083;
wire net6513;
wire net6514;
wire net9543;
wire net6515;
wire net6562;
wire net6518;
wire net11207;
wire net2963;
wire net6519;
wire net243;
wire net6520;
wire net1390;
wire net6523;
wire net6524;
wire net7709;
wire net4741;
wire net6823;
wire net6527;
wire net6529;
wire net8122;
wire net6077;
wire net6533;
wire net10068;
wire net6538;
wire net6544;
wire net6547;
wire net6552;
wire net2348;
wire net6553;
wire net6554;
wire net6685;
wire net7393;
wire net6557;
wire net5634;
wire net6558;
wire net10010;
wire net2820;
wire net6559;
wire net6561;
wire net6563;
wire net6567;
wire net9102;
wire net1583;
wire net5546;
wire net6568;
wire net10471;
wire net6570;
wire net1102;
wire net6575;
wire net4019;
wire net6577;
wire net1138;
wire net6581;
wire net10459;
wire net10325;
wire net3324;
wire net6582;
wire net9067;
wire net6583;
wire net781;
wire net6599;
wire net6586;
wire net6587;
wire net9702;
wire net6588;
wire net6589;
wire net6202;
wire net6590;
wire net6592;
wire net7534;
wire net6593;
wire net586;
wire net4514;
wire net7391;
wire net5438;
wire net6597;
wire net6605;
wire net6608;
wire net8079;
wire net6609;
wire net6632;
wire net3359;
wire net6610;
wire net10993;
wire net6611;
wire net8248;
wire net471;
wire net6613;
wire net6614;
wire net3614;
wire net4538;
wire net6615;
wire net6616;
wire net6620;
wire net4312;
wire net6621;
wire net6624;
wire net6627;
wire net9558;
wire net6633;
wire net6643;
wire net6648;
wire net6650;
wire net9874;
wire net6656;
wire net8490;
wire net6662;
wire net277;
wire net6665;
wire net5869;
wire net6670;
wire net6672;
wire net6675;
wire net6678;
wire net5848;
wire net6679;
wire net6683;
wire net2350;
wire net6688;
wire net4681;
wire net6690;
wire net6694;
wire net6696;
wire net6704;
wire net1337;
wire net827;
wire net6709;
wire net11117;
wire net7734;
wire net5484;
wire net4984;
wire net6969;
wire net6710;
wire net8892;
wire net3675;
wire net5065;
wire net6711;
wire net3746;
wire net6713;
wire net10392;
wire net6716;
wire net6719;
wire net2410;
wire net6340;
wire net6722;
wire net6726;
wire net7252;
wire net6728;
wire net5521;
wire net6729;
wire net8757;
wire net6734;
wire net4582;
wire net5187;
wire net6736;
wire net547;
wire net6741;
wire net6746;
wire net6747;
wire net9501;
wire net1198;
wire net6748;
wire net6749;
wire net6750;
wire net3253;
wire net6751;
wire net6752;
wire net3190;
wire net1328;
wire net6754;
wire net10188;
wire net9763;
wire net5220;
wire net6755;
wire net6929;
wire net6756;
wire net10643;
wire net6757;
wire net6762;
wire net11226;
wire net10697;
wire net7334;
wire net5318;
wire net6765;
wire net5968;
wire net6768;
wire net2340;
wire net6769;
wire net7232;
wire net6771;
wire net10373;
wire net6772;
wire net2382;
wire net109;
wire net7437;
wire net6773;
wire net1362;
wire net7146;
wire net6775;
wire net6777;
wire net6778;
wire net987;
wire net7236;
wire net6779;
wire net7050;
wire net6780;
wire net5997;
wire net6781;
wire net6794;
wire net6783;
wire net9664;
wire net165;
wire net4573;
wire net6788;
wire net6789;
wire net7062;
wire net6795;
wire net6207;
wire net6798;
wire net6801;
wire net3079;
wire net6802;
wire net7150;
wire net6803;
wire net6805;
wire net6807;
wire net6808;
wire net1659;
wire net6809;
wire net6814;
wire net6815;
wire net8700;
wire net6099;
wire net6817;
wire net6820;
wire net6825;
wire net4353;
wire net6827;
wire net11182;
wire net1782;
wire net6828;
wire net8794;
wire net6829;
wire net1988;
wire net6830;
wire net8583;
wire net6831;
wire net9563;
wire net6833;
wire net6835;
wire net6836;
wire net6837;
wire net806;
wire net6840;
wire net2207;
wire net5795;
wire net6841;
wire net6846;
wire net6847;
wire net6848;
wire net6851;
wire net9024;
wire net6854;
wire net11193;
wire net5569;
wire net6855;
wire net6857;
wire net8944;
wire net6859;
wire net151;
wire net6860;
wire net1905;
wire net6863;
wire net540;
wire net6869;
wire net6870;
wire net8052;
wire net1275;
wire net2315;
wire net6871;
wire net6873;
wire net5330;
wire net6874;
wire net1582;
wire net6878;
wire net6880;
wire net9593;
wire net6883;
wire net6886;
wire net6889;
wire net6891;
wire net9832;
wire net325;
wire net56;
wire net6893;
wire net6896;
wire net1794;
wire net6898;
wire net5771;
wire net6900;
wire net2148;
wire net4346;
wire net7375;
wire net6904;
wire net6906;
wire net6910;
wire net705;
wire net6912;
wire net6920;
wire net6925;
wire net10349;
wire net9718;
wire net6926;
wire net6931;
wire net5594;
wire net6935;
wire net4406;
wire net6937;
wire net6938;
wire net6939;
wire net4004;
wire net6942;
wire net1151;
wire net6943;
wire net6944;
wire net4175;
wire net6945;
wire net6947;
wire net399;
wire net6950;
wire net6952;
wire net6953;
wire net2993;
wire net6955;
wire net3863;
wire net6959;
wire net4407;
wire net6962;
wire net6963;
wire net4649;
wire net6964;
wire net2977;
wire net6966;
wire net786;
wire net7114;
wire net6967;
wire net3135;
wire net6970;
wire net2664;
wire net6972;
wire net6974;
wire net6983;
wire net10406;
wire net2682;
wire net6984;
wire net7121;
wire net6027;
wire net6985;
wire net413;
wire net6992;
wire net9842;
wire net7446;
wire net6995;
wire net7580;
wire net3987;
wire net6999;
wire net11055;
wire net7004;
wire net8137;
wire net805;
wire net7005;
wire net1239;
wire net7007;
wire net6024;
wire net5211;
wire net7008;
wire net7010;
wire net7012;
wire net7013;
wire net7014;
wire net7017;
wire net7019;
wire net7697;
wire net7228;
wire net10528;
wire net7020;
wire net7027;
wire net7030;
wire net7032;
wire net7033;
wire net7035;
wire net7036;
wire net7038;
wire net2186;
wire net7096;
wire net7040;
wire net9560;
wire net5868;
wire net7041;
wire net7992;
wire net7045;
wire net7049;
wire net7052;
wire net7055;
wire net23;
wire net7056;
wire net7058;
wire net7063;
wire net3501;
wire net3656;
wire net1805;
wire net7064;
wire net9910;
wire net1334;
wire net7066;
wire net7068;
wire net7077;
wire net7083;
wire net4563;
wire net7086;
wire net10273;
wire net304;
wire net7087;
wire net1370;
wire net7088;
wire net5005;
wire net7089;
wire net7091;
wire net7842;
wire net7098;
wire net7325;
wire net3806;
wire net7100;
wire net7105;
wire net7106;
wire net5102;
wire net7108;
wire net9914;
wire net7110;
wire net8565;
wire net7112;
wire net3553;
wire net7113;
wire net7116;
wire net7119;
wire net7128;
wire net7129;
wire net7133;
wire net7783;
wire net2727;
wire net7134;
wire net10803;
wire net10441;
wire net7135;
wire net7136;
wire net7138;
wire net10521;
wire net7140;
wire net7141;
wire net7143;
wire net5689;
wire net7144;
wire net7148;
wire net9487;
wire net7149;
wire net7673;
wire net6718;
wire net7152;
wire net9971;
wire net4843;
wire net7157;
wire net1624;
wire net7160;
wire net1320;
wire net7163;
wire net7851;
wire net7164;
wire net7165;
wire net1290;
wire net7167;
wire net5701;
wire net7168;
wire net7169;
wire net7496;
wire net6192;
wire net7171;
wire net1436;
wire net7172;
wire net9216;
wire net7173;
wire net7180;
wire net8535;
wire net7181;
wire net4320;
wire net7186;
wire net322;
wire net7188;
wire net7197;
wire net1176;
wire net7198;
wire net575;
wire net7199;
wire net1109;
wire net7200;
wire net307;
wire net7201;
wire net3733;
wire net7205;
wire net7207;
wire net7208;
wire net7209;
wire net7211;
wire net1708;
wire net7212;
wire net7076;
wire net7214;
wire net7215;
wire net9428;
wire net7217;
wire net7222;
wire net10975;
wire net9456;
wire net9109;
wire net7224;
wire net7225;
wire net9835;
wire net7067;
wire net7227;
wire net7229;
wire net9915;
wire net5941;
wire net7233;
wire net9395;
wire net3022;
wire net7234;
wire net8270;
wire net4310;
wire net7238;
wire net7240;
wire net7882;
wire net7243;
wire net5293;
wire net7248;
wire net7251;
wire net11066;
wire net7253;
wire net5892;
wire net1812;
wire net7254;
wire net6622;
wire net7255;
wire net5885;
wire net7258;
wire net7264;
wire net7780;
wire net4465;
wire net7266;
wire net7274;
wire net1875;
wire net7275;
wire net6635;
wire net7277;
wire net7280;
wire net7287;
wire net4456;
wire net7291;
wire net9999;
wire net7292;
wire net7297;
wire net7298;
wire net7301;
wire net1877;
wire net7304;
wire net7305;
wire net9008;
wire net7307;
wire net7308;
wire net3865;
wire net7313;
wire net7317;
wire net9564;
wire net7318;
wire net1680;
wire net7322;
wire net10744;
wire net7333;
wire net10740;
wire net7337;
wire net9232;
wire net7339;
wire net7340;
wire net7341;
wire net7342;
wire net7343;
wire net7350;
wire net8364;
wire net6521;
wire net7351;
wire net7352;
wire net1430;
wire net7357;
wire net7360;
wire net7362;
wire net7434;
wire net8473;
wire net7365;
wire net7366;
wire net7367;
wire net7574;
wire net3351;
wire net7369;
wire net11074;
wire net7371;
wire net5765;
wire net7373;
wire net9495;
wire net7376;
wire net8659;
wire net7377;
wire net7380;
wire net5343;
wire net7383;
wire net1019;
wire net7392;
wire net9546;
wire net7394;
wire net10170;
wire net61;
wire net7395;
wire net7397;
wire net7399;
wire net7401;
wire net9552;
wire net7403;
wire net1781;
wire net7404;
wire net7405;
wire net9472;
wire net7407;
wire net3778;
wire net6161;
wire net4468;
wire net3815;
wire net6116;
wire net7409;
wire net11171;
wire net10569;
wire net7411;
wire net7412;
wire net3515;
wire net4566;
wire net7413;
wire net10557;
wire net7420;
wire net6810;
wire net7422;
wire net2063;
wire net3883;
wire net6450;
wire net7424;
wire net4047;
wire net7426;
wire net4244;
wire net7436;
wire net6495;
wire net7153;
wire net7439;
wire net7442;
wire net7447;
wire net5463;
wire net7448;
wire net7449;
wire net7451;
wire net2900;
wire net7452;
wire net7856;
wire net7453;
wire net10978;
wire net7456;
wire net7459;
wire net4025;
wire net7468;
wire net10608;
wire net7471;
wire net3281;
wire net7472;
wire net7473;
wire net10832;
wire net5285;
wire net7474;
wire net7477;
wire net2173;
wire net7478;
wire net3606;
wire net7479;
wire net7482;
wire net3368;
wire net7485;
wire net7486;
INV_X32 c26(
.A(in20),
.ZN(net0)
);

INV_X4 c27(
.A(in17),
.ZN(net1)
);

XOR2_X2 c28(
.A(net0),
.B(in11),
.Z(net2)
);

INV_X1 c29(
.A(in10),
.ZN(net3)
);

XNOR2_X1 c30(
.A(net3),
.B(in2),
.ZN(net4)
);

INV_X2 c31(
.A(in8),
.ZN(net5)
);

INV_X8 c32(
.A(in17),
.ZN(net6)
);

INV_X16 c33(
.A(in2),
.ZN(net7)
);

OR3_X2 c34(
.A1(in21),
.A2(in9),
.A3(net0),
.ZN(net8)
);

INV_X32 c35(
.A(net8),
.ZN(net9)
);

OR2_X4 c36(
.A1(in22),
.A2(net2),
.ZN(net10)
);

INV_X4 c37(
.A(in3),
.ZN(net11)
);

OAI21_X2 c38(
.A(net9),
.B1(in6),
.B2(net40),
.ZN(net12)
);

OR2_X1 c39(
.A1(net5),
.A2(net3),
.ZN(net13)
);

XNOR2_X2 c40(
.A(net39),
.B(net2),
.ZN(net14)
);

OAI21_X1 c41(
.A(net7),
.B1(in0),
.B2(in12),
.ZN(net15)
);

INV_X1 c42(
.A(net10),
.ZN(net16)
);

INV_X2 c43(
.A(in15),
.ZN(net17)
);

INV_X8 c44(
.A(net39),
.ZN(net18)
);

INV_X16 c45(
.A(in6),
.ZN(net19)
);

INV_X32 c46(
.A(net17),
.ZN(net20)
);

AND2_X4 c47(
.A1(net18),
.A2(net39),
.ZN(net21)
);

INV_X4 c48(
.A(net14),
.ZN(net22)
);

INV_X1 c49(
.A(net22),
.ZN(net23)
);

INV_X2 c50(
.A(net3),
.ZN(net24)
);

INV_X8 c51(
.A(net8),
.ZN(net25)
);

AND2_X1 c52(
.A1(in0),
.A2(net2),
.ZN(net26)
);

INV_X16 c53(
.A(net23),
.ZN(net27)
);

INV_X32 c54(
.A(net1),
.ZN(net28)
);

AOI21_X2 c55(
.A(net23),
.B1(net27),
.B2(net18),
.ZN(net29)
);

INV_X4 c56(
.A(net28),
.ZN(net30)
);

INV_X1 c57(
.A(net20),
.ZN(net31)
);

AOI21_X1 c58(
.A(net13),
.B1(net1),
.B2(net31),
.ZN(net32)
);

NAND2_X1 c59(
.A1(net30),
.A2(net29),
.ZN(net33)
);

AOI21_X4 c60(
.A(net26),
.B1(net30),
.B2(net33),
.ZN(net34)
);

INV_X2 c61(
.A(net12),
.ZN(net35)
);

NAND2_X2 c62(
.A1(in22),
.A2(net31),
.ZN(net36)
);

NAND2_X4 c63(
.A1(net31),
.A2(net34),
.ZN(net37)
);

INV_X8 c64(
.A(in11),
.ZN(net38)
);

INV_X16 c65(
.A(in1),
.ZN(net39)
);

INV_X32 c66(
.A(in16),
.ZN(net40)
);

AND3_X1 c67(
.A1(net34),
.A2(in5),
.A3(net31),
.ZN(net41)
);

NAND3_X1 c68(
.A1(net2),
.A2(net31),
.A3(net3),
.ZN(net42)
);

INV_X4 c69(
.A(net42),
.ZN(net43)
);

NOR3_X4 c70(
.A1(net16),
.A2(net42),
.A3(net32),
.ZN(net44)
);

INV_X1 c71(
.A(net27),
.ZN(net45)
);

AND2_X2 c72(
.A1(in3),
.A2(net43),
.ZN(net46)
);

NOR3_X2 c73(
.A1(net32),
.A2(in18),
.A3(net45),
.ZN(net47)
);

XOR2_X1 c74(
.A(net40),
.B(net42),
.Z(net48)
);

NOR2_X1 c75(
.A1(net44),
.A2(in20),
.ZN(net49)
);

AND3_X4 c76(
.A1(net38),
.A2(net20),
.A3(net4),
.ZN(net50)
);

NAND3_X2 c77(
.A1(net15),
.A2(net38),
.A3(net12),
.ZN(net51)
);

OR3_X1 c78(
.A1(net4),
.A2(net10),
.A3(net11),
.ZN(net52)
);

MUX2_X1 c79(
.A(net11),
.B(net30),
.S(net49),
.Z(net53)
);

OAI21_X4 c80(
.A(net28),
.B1(net53),
.B2(net39),
.ZN(net54)
);

MUX2_X2 c81(
.A(net54),
.B(net44),
.S(in16),
.Z(net55)
);

NAND3_X4 c82(
.A1(net25),
.A2(net54),
.A3(net39),
.ZN(net56)
);

OR2_X2 c83(
.A1(net43),
.A2(net30),
.ZN(net57)
);

INV_X2 c84(
.A(net9658),
.ZN(net58)
);

INV_X8 c85(
.A(net30),
.ZN(net59)
);

OR3_X4 c86(
.A1(net24),
.A2(net106),
.A3(in13),
.ZN(net60)
);

INV_X16 c87(
.A(net47),
.ZN(net61)
);

NOR2_X4 c88(
.A1(net49),
.A2(net105),
.ZN(net62)
);

INV_X32 c89(
.A(net10399),
.ZN(net63)
);

INV_X4 c90(
.A(in14),
.ZN(net64)
);

INV_X1 c91(
.A(net40),
.ZN(net65)
);

INV_X2 c92(
.A(in13),
.ZN(net66)
);

INV_X8 c93(
.A(net36),
.ZN(net67)
);

INV_X16 c94(
.A(net43),
.ZN(net68)
);

INV_X32 c95(
.A(net9658),
.ZN(net69)
);

CLKGATETST_X1 c96(
.E(net58),
.SE(net106),
.CK(clk),
.GCK(net70)
);

INV_X4 c97(
.A(net105),
.ZN(net71)
);

INV_X1 c98(
.A(net36),
.ZN(net72)
);

INV_X2 c99(
.A(net104),
.ZN(net73)
);

INV_X8 c100(
.A(net71),
.ZN(net74)
);

NOR2_X2 c101(
.A1(in8),
.A2(net24),
.ZN(net75)
);

XOR2_X2 c102(
.A(net24),
.B(net40),
.Z(net76)
);

XNOR2_X1 c103(
.A(net69),
.B(net73),
.ZN(net77)
);

INV_X16 c104(
.A(net64),
.ZN(net78)
);

INV_X32 c105(
.A(net62),
.ZN(net79)
);

OR2_X4 c106(
.A1(net72),
.A2(net73),
.ZN(net80)
);

INV_X4 c107(
.A(net70),
.ZN(net81)
);

INV_X1 c108(
.A(net65),
.ZN(net82)
);

OR2_X1 c109(
.A1(net80),
.A2(net68),
.ZN(net83)
);

INV_X2 c110(
.A(net61),
.ZN(net84)
);

INV_X8 c111(
.A(net75),
.ZN(net85)
);

XNOR2_X2 c112(
.A(net72),
.B(net82),
.ZN(net86)
);

INV_X16 c113(
.A(net55),
.ZN(net87)
);

INV_X32 c114(
.A(in10),
.ZN(net88)
);

INV_X4 c115(
.A(net88),
.ZN(net89)
);

INV_X1 c116(
.A(net64),
.ZN(net90)
);

AND2_X4 c117(
.A1(net84),
.A2(net104),
.ZN(net91)
);

INV_X2 c118(
.A(net71),
.ZN(net92)
);

INV_X8 c119(
.A(net83),
.ZN(net93)
);

INV_X16 c120(
.A(net86),
.ZN(net94)
);

AND2_X1 c121(
.A1(net61),
.A2(net40),
.ZN(net95)
);

INV_X32 c122(
.A(net63),
.ZN(net96)
);

INV_X4 c123(
.A(net90),
.ZN(net97)
);

CLKGATETST_X2 c124(
.E(net81),
.SE(net37),
.CK(clk),
.GCK(net98)
);

NAND2_X1 c125(
.A1(net22),
.A2(net98),
.ZN(net99)
);

INV_X1 c126(
.A(in1),
.ZN(net100)
);

NAND2_X2 c127(
.A1(net69),
.A2(net55),
.ZN(net101)
);

DFFRS_X1 c128(
.D(net96),
.RN(net101),
.SN(net90),
.CK(clk),
.Q(net103),
.QN(net102)
);

INV_X2 c129(
.A(net13),
.ZN(net104)
);

INV_X8 c130(
.A(in14),
.ZN(net105)
);

INV_X16 c131(
.A(net55),
.ZN(net106)
);

INV_X32 c132(
.A(in18),
.ZN(net107)
);

INV_X4 c133(
.A(net79),
.ZN(net108)
);

CLKGATETST_X4 c134(
.E(net82),
.SE(net84),
.CK(clk),
.GCK(net109)
);

INV_X1 c135(
.A(net48),
.ZN(net110)
);

INV_X2 c136(
.A(net93),
.ZN(net111)
);

INV_X8 c137(
.A(net111),
.ZN(net112)
);

CLKGATETST_X8 c138(
.E(net84),
.SE(net87),
.CK(clk),
.GCK(net113)
);

NAND2_X4 c139(
.A1(net83),
.A2(net90),
.ZN(net114)
);

AND3_X2 c140(
.A1(net111),
.A2(net97),
.A3(net82),
.ZN(net115)
);

DFFR_X1 c141(
.D(net115),
.RN(net90),
.CK(clk),
.Q(net117),
.QN(net116)
);

DFFR_X2 c142(
.D(net112),
.RN(net109),
.CK(clk),
.Q(net119),
.QN(net118)
);

AND2_X2 c143(
.A1(net89),
.A2(net93),
.ZN(net120)
);

XOR2_X1 c144(
.A(net65),
.B(net108),
.Z(net121)
);

NOR2_X1 c145(
.A1(net118),
.A2(net10398),
.ZN(net122)
);

OR2_X2 c146(
.A1(net105),
.A2(net63),
.ZN(net123)
);

DFFRS_X2 c147(
.D(net101),
.RN(net55),
.SN(net74),
.CK(clk),
.Q(net125),
.QN(net124)
);

DFFS_X1 c148(
.D(net74),
.SN(net37),
.CK(clk),
.Q(net127),
.QN(net126)
);

DFFS_X2 c149(
.D(net87),
.SN(net122),
.CK(clk),
.Q(net129),
.QN(net128)
);

NOR2_X4 c150(
.A1(net127),
.A2(net58),
.ZN(net130)
);

NOR2_X2 c151(
.A1(net123),
.A2(net100),
.ZN(net131)
);

CLKGATETST_X1 c152(
.E(net80),
.SE(net115),
.CK(clk),
.GCK(net132)
);

XOR2_X2 c153(
.A(in18),
.B(net120),
.Z(net133)
);

NOR3_X1 c154(
.A1(net131),
.A2(net116),
.A3(net123),
.ZN(net134)
);

XNOR2_X1 c155(
.A(net97),
.B(net92),
.ZN(net135)
);

OR3_X2 c156(
.A1(net79),
.A2(net130),
.A3(net134),
.ZN(net136)
);

CLKGATETST_X2 c157(
.E(net121),
.SE(net126),
.CK(clk),
.GCK(net137)
);

OAI21_X2 c158(
.A(net109),
.B1(net124),
.B2(net137),
.ZN(net138)
);

SDFFRS_X1 c159(
.D(net134),
.RN(net136),
.SE(net135),
.SI(net120),
.SN(net87),
.CK(clk),
.Q(net140),
.QN(net139)
);

OAI21_X1 c160(
.A(net137),
.B1(net129),
.B2(net138),
.ZN(net141)
);

AOI21_X2 c161(
.A(net88),
.B1(net131),
.B2(net120),
.ZN(net142)
);

SDFFRS_X2 c162(
.D(net130),
.RN(net81),
.SE(net121),
.SI(net123),
.SN(net120),
.CK(clk),
.Q(net144),
.QN(net143)
);

AOI21_X1 c163(
.A(net125),
.B1(net5),
.B2(net72),
.ZN(net145)
);

AOI21_X4 c164(
.A(net135),
.B1(net102),
.B2(net137),
.ZN(net146)
);

OAI221_X4 c165(
.A(net103),
.B1(net145),
.B2(net141),
.C1(net132),
.C2(net120),
.ZN(net147)
);

INV_X16 c166(
.A(net76),
.ZN(net148)
);

INV_X32 c167(
.A(net48),
.ZN(net149)
);

OR2_X4 c168(
.A1(net149),
.A2(net94),
.ZN(net150)
);

INV_X4 c169(
.A(net9619),
.ZN(net151)
);

INV_X1 c170(
.A(in4),
.ZN(net152)
);

INV_X2 c171(
.A(net140),
.ZN(net153)
);

INV_X8 c172(
.A(net34),
.ZN(net154)
);

INV_X16 c173(
.A(net150),
.ZN(net155)
);

OR2_X1 c174(
.A1(net152),
.A2(net53),
.ZN(net156)
);

INV_X32 c175(
.A(net143),
.ZN(net157)
);

INV_X4 c176(
.A(net59),
.ZN(net158)
);

INV_X1 c177(
.A(net113),
.ZN(net159)
);

INV_X2 c178(
.A(net155),
.ZN(net160)
);

INV_X8 c179(
.A(net78),
.ZN(net161)
);

INV_X16 c180(
.A(net120),
.ZN(net162)
);

INV_X32 c181(
.A(net140),
.ZN(net163)
);

INV_X4 c182(
.A(net9619),
.ZN(net164)
);

INV_X1 c183(
.A(net163),
.ZN(net165)
);

XNOR2_X2 c184(
.A(net119),
.B(net113),
.ZN(net166)
);

AND3_X1 c185(
.A1(net119),
.A2(net113),
.A3(net85),
.ZN(net167)
);

INV_X2 c186(
.A(net146),
.ZN(net168)
);

INV_X8 c187(
.A(net53),
.ZN(net169)
);

AND2_X4 c188(
.A1(net166),
.A2(net132),
.ZN(net170)
);

INV_X16 c189(
.A(net148),
.ZN(net171)
);

INV_X32 c190(
.A(net164),
.ZN(net172)
);

INV_X4 c191(
.A(net99),
.ZN(net173)
);

AND2_X1 c192(
.A1(net145),
.A2(net170),
.ZN(net174)
);

INV_X1 c193(
.A(net172),
.ZN(net175)
);

INV_X2 c194(
.A(net171),
.ZN(net176)
);

INV_X8 c195(
.A(net9738),
.ZN(net177)
);

INV_X16 c196(
.A(net175),
.ZN(net178)
);

NAND2_X1 c197(
.A1(net169),
.A2(net53),
.ZN(net179)
);

NAND2_X2 c198(
.A1(net169),
.A2(net157),
.ZN(net180)
);

INV_X32 c199(
.A(in4),
.ZN(net181)
);

INV_X4 c200(
.A(net113),
.ZN(net182)
);

INV_X1 c201(
.A(net178),
.ZN(net183)
);

INV_X2 c202(
.A(in21),
.ZN(net184)
);

NAND2_X4 c203(
.A1(net76),
.A2(net167),
.ZN(net185)
);

NAND3_X1 c204(
.A1(net180),
.A2(net149),
.A3(net99),
.ZN(net186)
);

INV_X8 c205(
.A(net163),
.ZN(net187)
);

NOR3_X4 c206(
.A1(net144),
.A2(net48),
.A3(net177),
.ZN(net188)
);

AND2_X2 c207(
.A1(net184),
.A2(net159),
.ZN(net189)
);

XOR2_X1 c208(
.A(net177),
.B(net123),
.Z(net190)
);

NOR2_X1 c209(
.A1(net167),
.A2(net85),
.ZN(net191)
);

INV_X16 c210(
.A(net53),
.ZN(net192)
);

INV_X32 c211(
.A(net10717),
.ZN(net193)
);

INV_X4 c212(
.A(net174),
.ZN(net194)
);

OR2_X2 c213(
.A1(net191),
.A2(net158),
.ZN(net195)
);

NOR2_X4 c214(
.A1(net181),
.A2(net172),
.ZN(net196)
);

NOR2_X2 c215(
.A1(net146),
.A2(net151),
.ZN(net197)
);

INV_X1 c216(
.A(net195),
.ZN(net198)
);

INV_X2 c217(
.A(net195),
.ZN(net199)
);

NOR3_X2 c218(
.A1(net194),
.A2(net174),
.A3(net184),
.ZN(net200)
);

XOR2_X2 c219(
.A(net187),
.B(net169),
.Z(net201)
);

XNOR2_X1 c220(
.A(net201),
.B(net120),
.ZN(net202)
);

INV_X8 c221(
.A(net155),
.ZN(net203)
);

INV_X16 c222(
.A(net10684),
.ZN(net204)
);

AND3_X4 c223(
.A1(net199),
.A2(net172),
.A3(net185),
.ZN(net205)
);

INV_X32 c224(
.A(net99),
.ZN(net206)
);

CLKGATETST_X4 c225(
.E(net171),
.SE(net202),
.CK(clk),
.GCK(net207)
);

OR2_X4 c226(
.A1(net205),
.A2(net169),
.ZN(net208)
);

OR2_X1 c227(
.A1(net158),
.A2(net207),
.ZN(net209)
);

NAND3_X2 c228(
.A1(net78),
.A2(net197),
.A3(net202),
.ZN(net210)
);

INV_X4 c229(
.A(net200),
.ZN(net211)
);

OR3_X1 c230(
.A1(net176),
.A2(net118),
.A3(net10484),
.ZN(net212)
);

XNOR2_X2 c231(
.A(net179),
.B(net174),
.ZN(net213)
);

MUX2_X1 c232(
.A(net92),
.B(net110),
.S(net166),
.Z(net214)
);

OAI21_X4 c233(
.A(net203),
.B1(net191),
.B2(net139),
.ZN(net215)
);

AND2_X4 c234(
.A1(net204),
.A2(net176),
.ZN(net216)
);

AND2_X1 c235(
.A1(net182),
.A2(net10484),
.ZN(net217)
);

INV_X1 c236(
.A(net170),
.ZN(net218)
);

INV_X2 c237(
.A(net206),
.ZN(net219)
);

NAND2_X1 c238(
.A1(net209),
.A2(net156),
.ZN(net220)
);

OAI222_X2 c239(
.A1(net165),
.A2(net220),
.B1(net212),
.B2(net87),
.C1(net185),
.C2(net151),
.ZN(net221)
);

SDFF_X1 c240(
.D(net212),
.SE(net198),
.SI(net203),
.CK(clk),
.Q(net223),
.QN(net222)
);

NAND2_X2 c241(
.A1(net194),
.A2(net11141),
.ZN(net224)
);

MUX2_X2 c242(
.A(net201),
.B(net212),
.S(net11140),
.Z(net225)
);

NAND3_X4 c243(
.A1(net200),
.A2(net10484),
.A3(net11141),
.ZN(net226)
);

INV_X8 c244(
.A(net10307),
.ZN(net227)
);

OR3_X4 c245(
.A1(net227),
.A2(net205),
.A3(net10484),
.ZN(net228)
);

SDFF_X2 c246(
.D(net227),
.SE(net226),
.SI(net11141),
.CK(clk),
.Q(net230),
.QN(net229)
);

AND3_X2 c247(
.A1(net154),
.A2(net226),
.A3(net11140),
.ZN(net231)
);

NOR3_X1 c248(
.A1(net168),
.A2(net227),
.A3(net182),
.ZN(net232)
);

INV_X16 c249(
.A(net153),
.ZN(net233)
);

INV_X32 c250(
.A(net67),
.ZN(net234)
);

INV_X4 c251(
.A(net244),
.ZN(net235)
);

INV_X1 c252(
.A(net178),
.ZN(net236)
);

INV_X2 c253(
.A(net232),
.ZN(net237)
);

INV_X8 c254(
.A(net96),
.ZN(net238)
);

NAND2_X4 c255(
.A1(net233),
.A2(net166),
.ZN(net239)
);

INV_X16 c256(
.A(net11012),
.ZN(net240)
);

INV_X32 c257(
.A(net9593),
.ZN(net241)
);

INV_X4 c258(
.A(net16),
.ZN(net242)
);

INV_X1 c259(
.A(net73),
.ZN(net243)
);

INV_X2 c260(
.A(net94),
.ZN(net244)
);

INV_X8 c261(
.A(net188),
.ZN(net245)
);

INV_X16 c262(
.A(net25),
.ZN(net246)
);

INV_X32 c263(
.A(net73),
.ZN(net247)
);

INV_X4 c264(
.A(net5),
.ZN(net248)
);

INV_X1 c265(
.A(net217),
.ZN(net249)
);

INV_X2 c266(
.A(net242),
.ZN(net250)
);

INV_X8 c267(
.A(net240),
.ZN(net251)
);

AND2_X2 c268(
.A1(net173),
.A2(net235),
.ZN(net252)
);

XOR2_X1 c269(
.A(net157),
.B(net188),
.Z(net253)
);

NOR2_X1 c270(
.A1(net94),
.A2(net197),
.ZN(net254)
);

INV_X16 c271(
.A(net187),
.ZN(net255)
);

INV_X32 c272(
.A(net232),
.ZN(net256)
);

INV_X4 c273(
.A(net253),
.ZN(net257)
);

OR2_X2 c274(
.A1(net257),
.A2(net236),
.ZN(net258)
);

INV_X1 c275(
.A(net218),
.ZN(net259)
);

INV_X2 c276(
.A(net257),
.ZN(net260)
);

INV_X8 c277(
.A(net253),
.ZN(net261)
);

INV_X16 c278(
.A(net9592),
.ZN(net262)
);

OR3_X2 c279(
.A1(net254),
.A2(net249),
.A3(net262),
.ZN(net263)
);

OAI21_X2 c280(
.A(net258),
.B1(net234),
.B2(net261),
.ZN(net264)
);

NOR2_X4 c281(
.A1(net255),
.A2(net218),
.ZN(net265)
);

INV_X32 c282(
.A(net244),
.ZN(net266)
);

OAI21_X1 c283(
.A(net263),
.B1(net237),
.B2(net224),
.ZN(net267)
);

NOR2_X2 c284(
.A1(net266),
.A2(net243),
.ZN(net268)
);

XOR2_X2 c285(
.A(net197),
.B(net166),
.Z(net269)
);

XNOR2_X1 c286(
.A(net245),
.B(net173),
.ZN(net270)
);

INV_X4 c287(
.A(net238),
.ZN(net271)
);

INV_X1 c288(
.A(net236),
.ZN(net272)
);

INV_X2 c289(
.A(net9956),
.ZN(net273)
);

INV_X8 c290(
.A(net10926),
.ZN(net274)
);

INV_X16 c291(
.A(net10636),
.ZN(net275)
);

INV_X32 c292(
.A(net10782),
.ZN(net276)
);

AOI21_X2 c293(
.A(net249),
.B1(net265),
.B2(net179),
.ZN(net277)
);

OR2_X4 c294(
.A1(net256),
.A2(net141),
.ZN(net278)
);

INV_X4 c295(
.A(net166),
.ZN(net279)
);

DFFRS_X1 c296(
.D(net275),
.RN(net270),
.SN(net277),
.CK(clk),
.Q(net281),
.QN(net280)
);

OAI221_X2 c297(
.A(net272),
.B1(net217),
.B2(net178),
.C1(net251),
.C2(net276),
.ZN(net282)
);

INV_X1 c298(
.A(net279),
.ZN(net283)
);

INV_X2 c299(
.A(net282),
.ZN(net284)
);

AOI21_X1 c300(
.A(net153),
.B1(net264),
.B2(net240),
.ZN(net285)
);

OR2_X1 c301(
.A1(net271),
.A2(net235),
.ZN(net286)
);

DFFRS_X2 c302(
.D(net235),
.RN(net286),
.SN(net272),
.CK(clk),
.Q(net288),
.QN(net287)
);

XNOR2_X2 c303(
.A(net260),
.B(net270),
.ZN(net289)
);

AND2_X4 c304(
.A1(net241),
.A2(net280),
.ZN(net290)
);

INV_X8 c305(
.A(net273),
.ZN(net291)
);

INV_X16 c306(
.A(net10199),
.ZN(net292)
);

AND2_X1 c307(
.A1(net288),
.A2(net151),
.ZN(net293)
);

AOI21_X4 c308(
.A(net243),
.B1(net291),
.B2(net262),
.ZN(net294)
);

AND3_X1 c309(
.A1(net294),
.A2(net293),
.A3(net272),
.ZN(net295)
);

NAND2_X1 c310(
.A1(net239),
.A2(net218),
.ZN(net296)
);

NAND3_X1 c311(
.A1(net217),
.A2(net268),
.A3(net67),
.ZN(net297)
);

INV_X32 c312(
.A(net10898),
.ZN(net298)
);

NOR3_X4 c313(
.A1(net262),
.A2(net291),
.A3(net11042),
.ZN(net299)
);

NAND2_X2 c314(
.A1(net299),
.A2(net270),
.ZN(net300)
);

NOR3_X2 c315(
.A1(net293),
.A2(net276),
.A3(net10809),
.ZN(net301)
);

NAND2_X4 c316(
.A1(net237),
.A2(net258),
.ZN(net302)
);

INV_X4 c317(
.A(net10771),
.ZN(net303)
);

AND3_X4 c318(
.A1(net293),
.A2(net303),
.A3(net251),
.ZN(net304)
);

SDFF_X1 c319(
.D(net302),
.SE(net292),
.SI(net179),
.CK(clk),
.Q(net306),
.QN(net305)
);

INV_X1 c320(
.A(net291),
.ZN(net307)
);

AND2_X2 c321(
.A1(net307),
.A2(net257),
.ZN(net308)
);

NAND3_X2 c322(
.A1(net290),
.A2(net300),
.A3(net256),
.ZN(net309)
);

SDFFR_X1 c323(
.D(net240),
.RN(net291),
.SE(net309),
.SI(net277),
.CK(clk),
.Q(net311),
.QN(net310)
);

AOI222_X1 c324(
.A1(net304),
.A2(net311),
.B1(net309),
.B2(net265),
.C1(net251),
.C2(net11042),
.ZN(net312)
);

SDFF_X2 c325(
.D(net224),
.SE(net277),
.SI(net10809),
.CK(clk),
.Q(net314),
.QN(net313)
);

DFFRS_X1 c326(
.D(net264),
.RN(net293),
.SN(net299),
.CK(clk),
.Q(net316),
.QN(net315)
);

INV_X2 c327(
.A(net10806),
.ZN(net317)
);

XOR2_X1 c328(
.A(net300),
.B(net303),
.Z(net318)
);

OR3_X1 c329(
.A1(net318),
.A2(net309),
.ZN(net319)
);

SDFFRS_X1 c330(
.D(net284),
.RN(net290),
.SE(net191),
.SI(net318),
.SN(net10396),
.CK(clk),
.Q(net321),
.QN(net320)
);

AOI221_X4 c331(
.A(net317),
.B1(net187),
.B2(net320),
.C1(net166),
.C2(net10396),
.ZN(net322)
);

INV_X8 c332(
.A(net303),
.ZN(net323)
);

NOR2_X1 c333(
.A1(net132),
.A2(net283),
.ZN(net324)
);

INV_X16 c334(
.A(net159),
.ZN(net325)
);

INV_X32 c335(
.A(net159),
.ZN(net326)
);

OR2_X2 c336(
.A1(net230),
.A2(net151),
.ZN(net327)
);

NOR2_X4 c337(
.A1(net132),
.A2(net282),
.ZN(net328)
);

INV_X4 c338(
.A(net185),
.ZN(net329)
);

INV_X1 c339(
.A(net123),
.ZN(net330)
);

INV_X2 c340(
.A(net10949),
.ZN(net331)
);

INV_X8 c341(
.A(net11074),
.ZN(net332)
);

INV_X16 c342(
.A(net298),
.ZN(net333)
);

INV_X32 c343(
.A(net282),
.ZN(net334)
);

INV_X4 c344(
.A(net263),
.ZN(net335)
);

INV_X1 c345(
.A(net322),
.ZN(net336)
);

INV_X2 c346(
.A(net281),
.ZN(net337)
);

INV_X8 c347(
.A(net10289),
.ZN(net338)
);

INV_X16 c348(
.A(net316),
.ZN(net339)
);

INV_X32 c349(
.A(net313),
.ZN(net340)
);

INV_X4 c350(
.A(net333),
.ZN(net341)
);

INV_X1 c351(
.A(net262),
.ZN(net342)
);

INV_X2 c352(
.A(net265),
.ZN(net343)
);

NOR2_X2 c353(
.A1(net281),
.A2(net274),
.ZN(net344)
);

INV_X8 c354(
.A(net332),
.ZN(net345)
);

XOR2_X2 c355(
.A(net345),
.B(net338),
.Z(net346)
);

INV_X16 c356(
.A(net220),
.ZN(net347)
);

INV_X32 c357(
.A(net193),
.ZN(net348)
);

INV_X4 c358(
.A(in11),
.ZN(net349)
);

XNOR2_X1 c359(
.A(net349),
.B(net151),
.ZN(net350)
);

OR2_X4 c360(
.A1(net344),
.A2(in11),
.ZN(net351)
);

INV_X1 c361(
.A(net346),
.ZN(net352)
);

OR2_X1 c362(
.A1(net314),
.A2(net179),
.ZN(net353)
);

XNOR2_X2 c363(
.A(net349),
.B(net337),
.ZN(net354)
);

INV_X2 c364(
.A(net11074),
.ZN(net355)
);

AND2_X4 c365(
.A1(net233),
.A2(net348),
.ZN(net356)
);

AND2_X1 c366(
.A1(net341),
.A2(net326),
.ZN(net357)
);

INV_X8 c367(
.A(net356),
.ZN(net358)
);

INV_X16 c368(
.A(net9746),
.ZN(net359)
);

NAND2_X1 c369(
.A1(net355),
.A2(net328),
.ZN(net360)
);

NAND2_X2 c370(
.A1(net357),
.A2(net265),
.ZN(net361)
);

INV_X32 c371(
.A(net332),
.ZN(net362)
);

NAND2_X4 c372(
.A1(net216),
.A2(net351),
.ZN(net363)
);

INV_X4 c373(
.A(net274),
.ZN(net364)
);

MUX2_X1 c374(
.A(net329),
.B(net298),
.S(net323),
.Z(net365)
);

INV_X1 c375(
.A(net328),
.ZN(net366)
);

AND2_X2 c376(
.A1(net340),
.A2(net359),
.ZN(net367)
);

XOR2_X1 c377(
.A(net352),
.B(net356),
.Z(net368)
);

NOR2_X1 c378(
.A1(net359),
.A2(net356),
.ZN(net369)
);

INV_X2 c379(
.A(net10743),
.ZN(net370)
);

INV_X8 c380(
.A(net325),
.ZN(net371)
);

OR2_X2 c381(
.A1(net362),
.A2(net325),
.ZN(net372)
);

NOR2_X4 c382(
.A1(net358),
.A2(net355),
.ZN(net373)
);

NOR2_X2 c383(
.A1(net372),
.A2(net366),
.ZN(net374)
);

INV_X16 c384(
.A(net356),
.ZN(net375)
);

INV_X32 c385(
.A(net373),
.ZN(net376)
);

XOR2_X2 c386(
.A(net326),
.B(net370),
.Z(net377)
);

OAI21_X4 c387(
.A(net374),
.B1(net274),
.B2(net344),
.ZN(net378)
);

XNOR2_X1 c388(
.A(net361),
.B(net315),
.ZN(net379)
);

INV_X4 c389(
.A(net334),
.ZN(net380)
);

INV_X1 c390(
.A(net346),
.ZN(net381)
);

OR2_X4 c391(
.A1(net336),
.A2(net324),
.ZN(net382)
);

OR2_X1 c392(
.A1(net380),
.A2(net343),
.ZN(net383)
);

XNOR2_X2 c393(
.A(net348),
.B(net383),
.ZN(net384)
);

AND2_X4 c394(
.A1(net376),
.A2(net351),
.ZN(net385)
);

MUX2_X2 c395(
.A(net333),
.B(net379),
.S(net185),
.Z(net386)
);

NAND3_X4 c396(
.A1(net372),
.A2(net381),
.A3(net339),
.ZN(net387)
);

AND2_X1 c397(
.A1(net378),
.A2(net364),
.ZN(net388)
);

NAND2_X1 c398(
.A1(net384),
.A2(net331),
.ZN(net389)
);

NAND2_X2 c399(
.A1(net364),
.A2(net387),
.ZN(net390)
);

NAND2_X4 c400(
.A1(net360),
.A2(net10441),
.ZN(net391)
);

OR3_X4 c401(
.A1(net366),
.A2(net358),
.A3(net10441),
.ZN(net392)
);

DFFRS_X2 c402(
.D(net347),
.RN(net377),
.SN(net357),
.CK(clk),
.Q(net394),
.QN(net393)
);

AND3_X2 c403(
.A1(net375),
.A2(net382),
.A3(net385),
.ZN(net395)
);

AND2_X2 c404(
.A1(net374),
.A2(net10441),
.ZN(net396)
);

XOR2_X1 c405(
.A(net395),
.B(net344),
.Z(net397)
);

NOR2_X1 c406(
.A1(net387),
.A2(net396),
.ZN(net398)
);

NOR3_X1 c407(
.A1(net390),
.A2(net326),
.A3(net10441),
.ZN(net399)
);

INV_X2 c408(
.A(net10811),
.ZN(net400)
);

SDFF_X1 c409(
.D(net381),
.SE(net396),
.SI(net400),
.CK(clk),
.Q(net402),
.QN(net401)
);

OR4_X4 c410(
.A1(net400),
.A2(net376),
.A3(net402),
.A4(net397),
.ZN(net403)
);

SDFFR_X2 c411(
.D(net369),
.RN(net403),
.SE(net391),
.SI(net400),
.CK(clk),
.Q(net405),
.QN(net404)
);

OAI22_X2 c412(
.A1(net367),
.A2(net396),
.B1(net397),
.B2(net403),
.ZN(net406)
);

OR3_X2 c413(
.A1(net382),
.A2(net367),
.A3(net10728),
.ZN(net407)
);

OAI211_X4 c414(
.A(net379),
.B(net387),
.C1(net397),
.C2(net400),
.ZN(net408)
);

INV_X8 c415(
.A(net301),
.ZN(net409)
);

INV_X16 c416(
.A(net383),
.ZN(net410)
);

INV_X32 c417(
.A(net409),
.ZN(net411)
);

INV_X4 c418(
.A(net9790),
.ZN(net412)
);

OR2_X2 c419(
.A1(net373),
.A2(net392),
.ZN(net413)
);

OAI21_X2 c420(
.A(net397),
.B1(net409),
.B2(net342),
.ZN(net414)
);

INV_X1 c421(
.A(net411),
.ZN(net415)
);

NOR2_X4 c422(
.A1(net405),
.A2(net385),
.ZN(net416)
);

INV_X2 c423(
.A(net415),
.ZN(net417)
);

INV_X8 c424(
.A(net324),
.ZN(net418)
);

NOR2_X2 c425(
.A1(net141),
.A2(net147),
.ZN(net419)
);

INV_X16 c426(
.A(net324),
.ZN(net420)
);

INV_X32 c427(
.A(net383),
.ZN(net421)
);

XOR2_X2 c428(
.A(net420),
.B(net365),
.Z(net422)
);

OAI211_X1 c429(
.A(net404),
.B(net417),
.C1(net295),
.C2(net338),
.ZN(net423)
);

XNOR2_X1 c430(
.A(net329),
.B(net321),
.ZN(net424)
);

INV_X4 c431(
.A(net250),
.ZN(net425)
);

OR2_X4 c432(
.A1(net407),
.A2(net303),
.ZN(net426)
);

INV_X1 c433(
.A(net425),
.ZN(net427)
);

INV_X2 c434(
.A(net295),
.ZN(net428)
);

INV_X8 c435(
.A(net336),
.ZN(net429)
);

INV_X16 c436(
.A(net33),
.ZN(net430)
);

INV_X32 c437(
.A(net429),
.ZN(net431)
);

INV_X4 c438(
.A(net9548),
.ZN(net432)
);

OR2_X1 c439(
.A1(net283),
.A2(net426),
.ZN(net433)
);

INV_X1 c440(
.A(net371),
.ZN(net434)
);

INV_X2 c441(
.A(net254),
.ZN(net435)
);

INV_X8 c442(
.A(net192),
.ZN(net436)
);

INV_X16 c443(
.A(net432),
.ZN(net437)
);

XNOR2_X2 c444(
.A(net162),
.B(net412),
.ZN(net438)
);

AND2_X4 c445(
.A1(net433),
.A2(net429),
.ZN(net439)
);

AND2_X1 c446(
.A1(net426),
.A2(net301),
.ZN(net440)
);

OAI21_X1 c447(
.A(net417),
.B1(net432),
.B2(net426),
.ZN(net441)
);

NAND2_X1 c448(
.A1(net430),
.A2(net435),
.ZN(net442)
);

INV_X32 c449(
.A(net431),
.ZN(net443)
);

NAND2_X2 c450(
.A1(net399),
.A2(net432),
.ZN(net444)
);

AOI21_X2 c451(
.A(net413),
.B1(net428),
.B2(net440),
.ZN(net445)
);

INV_X4 c452(
.A(net9548),
.ZN(net446)
);

INV_X1 c453(
.A(net10380),
.ZN(net447)
);

INV_X2 c454(
.A(net428),
.ZN(net448)
);

INV_X8 c455(
.A(net10380),
.ZN(net449)
);

NAND2_X4 c456(
.A1(net394),
.A2(net435),
.ZN(net450)
);

INV_X16 c457(
.A(net430),
.ZN(net451)
);

INV_X32 c458(
.A(net11060),
.ZN(net452)
);

INV_X4 c459(
.A(net9788),
.ZN(net453)
);

AOI21_X1 c460(
.A(net295),
.B1(net447),
.B2(net436),
.ZN(net454)
);

INV_X1 c461(
.A(net9788),
.ZN(net455)
);

AOI21_X4 c462(
.A(net322),
.B1(net441),
.B2(net443),
.ZN(net456)
);

AND2_X2 c463(
.A1(net446),
.A2(net301),
.ZN(net457)
);

INV_X2 c464(
.A(net456),
.ZN(net458)
);

INV_X8 c465(
.A(net9941),
.ZN(net459)
);

AND3_X1 c466(
.A1(net444),
.A2(net343),
.A3(net425),
.ZN(net460)
);

XOR2_X1 c467(
.A(net429),
.B(net443),
.Z(net461)
);

NOR2_X1 c468(
.A1(net67),
.A2(net423),
.ZN(net462)
);

OR2_X2 c469(
.A1(net413),
.A2(net435),
.ZN(net463)
);

NOR2_X4 c470(
.A1(net448),
.A2(net453),
.ZN(net464)
);

INV_X16 c471(
.A(net452),
.ZN(net465)
);

INV_X32 c472(
.A(net444),
.ZN(net466)
);

NOR2_X2 c473(
.A1(net464),
.A2(net254),
.ZN(net467)
);

NAND3_X1 c474(
.A1(net424),
.A2(net448),
.A3(net415),
.ZN(net468)
);

NOR3_X4 c475(
.A1(net412),
.A2(net322),
.A3(net449),
.ZN(net469)
);

XOR2_X2 c476(
.A(net420),
.B(net399),
.Z(net470)
);

SDFF_X2 c477(
.D(net451),
.SE(net431),
.SI(net393),
.CK(clk),
.Q(net472),
.QN(net471)
);

INV_X4 c478(
.A(net466),
.ZN(net473)
);

NOR3_X2 c479(
.A1(net473),
.A2(net464),
.A3(net471),
.ZN(net474)
);

AND3_X4 c480(
.A1(net416),
.A2(net362),
.A3(net10579),
.ZN(net475)
);

XNOR2_X1 c481(
.A(net439),
.B(net461),
.ZN(net476)
);

INV_X1 c482(
.A(net342),
.ZN(net477)
);

INV_X2 c483(
.A(net477),
.ZN(net478)
);

INV_X8 c484(
.A(net10781),
.ZN(net479)
);

OR2_X4 c485(
.A1(net478),
.A2(net10897),
.ZN(net480)
);

NAND3_X2 c486(
.A1(net470),
.A2(net478),
.A3(net10781),
.ZN(net481)
);

OR3_X1 c487(
.A1(net422),
.A2(net446),
.A3(net473),
.ZN(net482)
);

MUX2_X1 c488(
.A(net475),
.B(net420),
.S(net434),
.Z(net483)
);

OAI21_X4 c489(
.A(net447),
.B1(net350),
.B2(net439),
.ZN(net484)
);

DFFRS_X1 c490(
.D(net469),
.RN(net440),
.SN(net451),
.CK(clk),
.Q(net486),
.QN(net485)
);

MUX2_X2 c491(
.A(net485),
.B(net432),
.S(net10897),
.Z(net487)
);

SDFFRS_X2 c492(
.D(net483),
.RN(net440),
.SE(net481),
.SI(net403),
.SN(net476),
.CK(clk),
.Q(net489),
.QN(net488)
);

OR2_X1 c493(
.A1(net486),
.A2(net446),
.ZN(net490)
);

INV_X16 c494(
.A(net10132),
.ZN(net491)
);

CLKGATETST_X8 c495(
.E(net468),
.SE(net427),
.CK(clk),
.GCK(net492)
);

NAND3_X4 c496(
.A1(net491),
.A2(net490),
.A3(net394),
.ZN(net493)
);

OR3_X4 c497(
.A1(net493),
.A2(net490),
.A3(net481),
.ZN(net494)
);

INV_X32 c498(
.A(net9659),
.ZN(net495)
);

INV_X4 c499(
.A(net385),
.ZN(net496)
);

XNOR2_X2 c500(
.A(net489),
.B(net520),
.ZN(net497)
);

AND2_X4 c501(
.A1(net57),
.A2(net510),
.ZN(net498)
);

INV_X1 c502(
.A(net523),
.ZN(net499)
);

INV_X2 c503(
.A(net498),
.ZN(net500)
);

AND2_X1 c504(
.A1(net512),
.A2(net525),
.ZN(net501)
);

INV_X8 c505(
.A(net338),
.ZN(net502)
);

NAND2_X1 c506(
.A1(net501),
.A2(net494),
.ZN(net503)
);

INV_X16 c507(
.A(net512),
.ZN(net504)
);

NAND2_X2 c508(
.A1(net521),
.A2(net496),
.ZN(net505)
);

NAND2_X4 c509(
.A1(net505),
.A2(net524),
.ZN(net506)
);

INV_X32 c510(
.A(net10830),
.ZN(net507)
);

INV_X4 c511(
.A(net151),
.ZN(net508)
);

INV_X1 c512(
.A(net510),
.ZN(net509)
);

INV_X2 c513(
.A(net9659),
.ZN(net510)
);

AND2_X2 c514(
.A1(net466),
.A2(net251),
.ZN(net511)
);

INV_X8 c515(
.A(net151),
.ZN(net512)
);

INV_X16 c516(
.A(net487),
.ZN(net513)
);

INV_X32 c517(
.A(net457),
.ZN(net514)
);

INV_X4 c518(
.A(net391),
.ZN(net515)
);

INV_X1 c519(
.A(net321),
.ZN(net516)
);

INV_X2 c520(
.A(net511),
.ZN(net517)
);

INV_X8 c521(
.A(net460),
.ZN(net518)
);

INV_X16 c522(
.A(net391),
.ZN(net519)
);

INV_X32 c523(
.A(net9896),
.ZN(net520)
);

XOR2_X1 c524(
.A(net446),
.B(net455),
.Z(net521)
);

INV_X4 c525(
.A(net392),
.ZN(net522)
);

INV_X1 c526(
.A(net470),
.ZN(net523)
);

INV_X2 c527(
.A(net338),
.ZN(net524)
);

DFFR_X1 c528(
.D(net353),
.RN(net517),
.CK(clk),
.Q(net526),
.QN(net525)
);

INV_X8 c529(
.A(net497),
.ZN(net527)
);

DFFRS_X2 c530(
.D(net353),
.RN(net392),
.SN(net355),
.CK(clk),
.Q(net529),
.QN(net528)
);

NOR2_X1 c531(
.A1(net523),
.A2(net524),
.ZN(net530)
);

OR2_X2 c532(
.A1(net433),
.A2(net33),
.ZN(net531)
);

NOR2_X4 c533(
.A1(net524),
.A2(net11047),
.ZN(net532)
);

NOR2_X2 c534(
.A1(net361),
.A2(net514),
.ZN(net533)
);

XOR2_X2 c535(
.A(net533),
.B(net509),
.Z(net534)
);

INV_X16 c536(
.A(net529),
.ZN(net535)
);

AND3_X2 c537(
.A1(net508),
.A2(net351),
.A3(net482),
.ZN(net536)
);

XNOR2_X1 c538(
.A(net532),
.B(net509),
.ZN(net537)
);

INV_X32 c539(
.A(net10345),
.ZN(net538)
);

NOR3_X1 c540(
.A1(net484),
.A2(net437),
.A3(net461),
.ZN(net539)
);

OR2_X4 c541(
.A1(net496),
.A2(net509),
.ZN(net540)
);

OR2_X1 c542(
.A1(net385),
.A2(net504),
.ZN(net541)
);

XNOR2_X2 c543(
.A(net446),
.B(net10518),
.ZN(net542)
);

AND2_X4 c544(
.A1(net462),
.A2(net528),
.ZN(net543)
);

AND2_X1 c545(
.A1(net538),
.A2(net532),
.ZN(net544)
);

NAND2_X1 c546(
.A1(net479),
.A2(net492),
.ZN(net545)
);

INV_X4 c547(
.A(net502),
.ZN(net546)
);

NAND2_X2 c548(
.A1(net541),
.A2(net500),
.ZN(net547)
);

NAND2_X4 c549(
.A1(net10518),
.A2(net11047),
.ZN(net548)
);

AND2_X2 c550(
.A1(net545),
.A2(net538),
.ZN(net549)
);

XOR2_X1 c551(
.A(net509),
.B(net535),
.Z(net550)
);

NOR2_X1 c552(
.A1(net550),
.A2(net547),
.ZN(net551)
);

OR2_X2 c553(
.A1(net547),
.A2(net545),
.ZN(net552)
);

NOR2_X4 c554(
.A1(net549),
.A2(net530),
.ZN(net553)
);

NOR2_X2 c555(
.A1(net541),
.A2(net548),
.ZN(net554)
);

XOR2_X2 c556(
.A(net544),
.B(net426),
.Z(net555)
);

SDFFRS_X1 c557(
.D(net507),
.RN(net521),
.SE(net192),
.SI(net551),
.SN(net459),
.CK(clk),
.Q(net557),
.QN(net556)
);

XNOR2_X1 c558(
.A(net524),
.B(net512),
.ZN(net558)
);

DFFR_X2 c559(
.D(net501),
.RN(net553),
.CK(clk),
.Q(net560),
.QN(net559)
);

AOI222_X4 c560(
.A1(net520),
.A2(net532),
.B1(net508),
.B2(net512),
.C1(net551),
.C2(net559),
.ZN(net561)
);

OR3_X2 c561(
.A1(net526),
.A2(net507),
.A3(net459),
.ZN(net562)
);

OR2_X4 c562(
.A1(net513),
.A2(net550),
.ZN(net563)
);

OR2_X1 c563(
.A1(net456),
.A2(net543),
.ZN(net564)
);

XNOR2_X2 c564(
.A(net497),
.B(net547),
.ZN(net565)
);

INV_X1 c565(
.A(net10830),
.ZN(net566)
);

OAI21_X2 c566(
.A(net563),
.B1(net549),
.B2(net562),
.ZN(net567)
);

AND2_X4 c567(
.A1(net534),
.A2(net527),
.ZN(net568)
);

DFFS_X1 c568(
.D(net565),
.SN(net566),
.CK(clk),
.Q(net570),
.QN(net569)
);

AND2_X1 c569(
.A1(net558),
.A2(net524),
.ZN(net571)
);

INV_X2 c570(
.A(net11088),
.ZN(net572)
);

NAND2_X1 c571(
.A1(net437),
.A2(net556),
.ZN(net573)
);

NAND2_X2 c572(
.A1(net531),
.A2(net11143),
.ZN(net574)
);

NAND2_X4 c573(
.A1(net567),
.A2(net573),
.ZN(net575)
);

OAI21_X1 c574(
.A(net557),
.B1(net575),
.B2(net11142),
.ZN(net576)
);

AND2_X2 c575(
.A1(net334),
.A2(net569),
.ZN(net577)
);

INV_X8 c576(
.A(net11056),
.ZN(net578)
);

SDFF_X1 c577(
.D(net494),
.SE(net565),
.SI(net578),
.CK(clk),
.Q(net580),
.QN(net579)
);

AOI21_X2 c578(
.A(net542),
.B1(net479),
.B2(net575),
.ZN(net581)
);

OAI33_X1 c579(
.A1(net572),
.A2(net487),
.A3(net581),
.B1(net578),
.B2(net551),
.B3(net10804),
.ZN(net582)
);

AOI222_X2 c580(
.A1(net495),
.A2(net574),
.B1(net579),
.B2(net509),
.C1(net578),
.C2(net11145),
.ZN(net583)
);

INV_X16 c581(
.A(net511),
.ZN(net584)
);

INV_X32 c582(
.A(net440),
.ZN(net585)
);

INV_X4 c583(
.A(net9969),
.ZN(net586)
);

INV_X1 c584(
.A(net492),
.ZN(net587)
);

INV_X2 c585(
.A(net368),
.ZN(net588)
);

XOR2_X1 c586(
.A(net577),
.B(net555),
.Z(net589)
);

INV_X8 c587(
.A(net9560),
.ZN(net590)
);

NOR2_X1 c588(
.A1(net562),
.A2(net441),
.ZN(net591)
);

INV_X16 c589(
.A(net566),
.ZN(net592)
);

INV_X32 c590(
.A(net502),
.ZN(net593)
);

OR2_X2 c591(
.A1(net546),
.A2(net354),
.ZN(net594)
);

INV_X4 c592(
.A(net85),
.ZN(net595)
);

NOR2_X4 c593(
.A1(net504),
.A2(net546),
.ZN(net596)
);

INV_X1 c594(
.A(net77),
.ZN(net597)
);

NOR2_X2 c595(
.A1(net555),
.A2(net586),
.ZN(net598)
);

XOR2_X2 c596(
.A(net436),
.B(net580),
.Z(net599)
);

INV_X2 c597(
.A(net461),
.ZN(net600)
);

INV_X8 c598(
.A(net354),
.ZN(net601)
);

INV_X16 c599(
.A(net548),
.ZN(net602)
);

INV_X32 c600(
.A(net596),
.ZN(net603)
);

INV_X4 c601(
.A(net586),
.ZN(net604)
);

INV_X1 c602(
.A(net9560),
.ZN(net605)
);

INV_X2 c603(
.A(net504),
.ZN(net606)
);

INV_X8 c604(
.A(net592),
.ZN(net607)
);

INV_X16 c605(
.A(net597),
.ZN(net608)
);

AOI21_X1 c606(
.A(net426),
.B1(net598),
.B2(net601),
.ZN(net609)
);

XNOR2_X1 c607(
.A(net461),
.B(net586),
.ZN(net610)
);

INV_X32 c608(
.A(net492),
.ZN(net611)
);

OR2_X4 c609(
.A1(net603),
.A2(net586),
.ZN(net612)
);

INV_X4 c610(
.A(net601),
.ZN(net613)
);

INV_X1 c611(
.A(net608),
.ZN(net614)
);

INV_X2 c612(
.A(net580),
.ZN(net615)
);

INV_X8 c613(
.A(net9734),
.ZN(net616)
);

INV_X16 c614(
.A(net613),
.ZN(net617)
);

OR2_X1 c615(
.A1(net603),
.A2(net593),
.ZN(net618)
);

XNOR2_X2 c616(
.A(net593),
.B(net573),
.ZN(net619)
);

AND2_X4 c617(
.A1(net607),
.A2(net535),
.ZN(net620)
);

AND2_X1 c618(
.A1(net602),
.A2(net607),
.ZN(net621)
);

NAND2_X1 c619(
.A1(net604),
.A2(net621),
.ZN(net622)
);

INV_X32 c620(
.A(net537),
.ZN(net623)
);

AOI21_X4 c621(
.A(net610),
.B1(net614),
.B2(net601),
.ZN(net624)
);

INV_X4 c622(
.A(net621),
.ZN(net625)
);

NAND2_X2 c623(
.A1(net591),
.A2(net607),
.ZN(net626)
);

INV_X1 c624(
.A(net9765),
.ZN(net627)
);

NAND2_X4 c625(
.A1(net625),
.A2(net354),
.ZN(net628)
);

DFFS_X2 c626(
.D(net599),
.SN(net502),
.CK(clk),
.Q(net630),
.QN(net629)
);

INV_X2 c627(
.A(net585),
.ZN(net631)
);

AND2_X2 c628(
.A1(net600),
.A2(net594),
.ZN(net632)
);

INV_X8 c629(
.A(net607),
.ZN(net633)
);

INV_X16 c630(
.A(net630),
.ZN(net634)
);

XOR2_X1 c631(
.A(net590),
.B(net581),
.Z(net635)
);

AND3_X1 c632(
.A1(net619),
.A2(net560),
.A3(net587),
.ZN(net636)
);

NOR2_X1 c633(
.A1(net441),
.A2(net602),
.ZN(net637)
);

CLKGATETST_X1 c634(
.E(net628),
.SE(net626),
.CK(clk),
.GCK(net638)
);

INV_X32 c635(
.A(net595),
.ZN(net639)
);

INV_X4 c636(
.A(net9790),
.ZN(net640)
);

NAND3_X1 c637(
.A1(net639),
.A2(net593),
.A3(net626),
.ZN(net641)
);

INV_X1 c638(
.A(net622),
.ZN(net642)
);

INV_X2 c639(
.A(net614),
.ZN(net643)
);

INV_X8 c640(
.A(net10196),
.ZN(net644)
);

INV_X16 c641(
.A(net617),
.ZN(net645)
);

OR2_X2 c642(
.A1(net623),
.A2(net616),
.ZN(net646)
);

NOR2_X4 c643(
.A1(net633),
.A2(net628),
.ZN(net647)
);

NOR3_X4 c644(
.A1(net562),
.A2(net640),
.A3(net633),
.ZN(net648)
);

NOR2_X2 c645(
.A1(net647),
.A2(net624),
.ZN(net649)
);

CLKGATETST_X2 c646(
.E(net617),
.SE(net632),
.CK(clk),
.GCK(net650)
);

CLKGATETST_X4 c647(
.E(net624),
.SE(net434),
.CK(clk),
.GCK(net651)
);

XOR2_X2 c648(
.A(net495),
.B(net640),
.Z(net652)
);

CLKGATETST_X8 c649(
.E(net631),
.SE(net627),
.CK(clk),
.GCK(net653)
);

INV_X32 c650(
.A(net616),
.ZN(net654)
);

NOR3_X2 c651(
.A1(net588),
.A2(net585),
.A3(net368),
.ZN(net655)
);

SDFF_X2 c652(
.D(net655),
.SE(net628),
.SI(net10782),
.CK(clk),
.Q(net657),
.QN(net656)
);

INV_X4 c653(
.A(net652),
.ZN(net658)
);

AND3_X4 c654(
.A1(net658),
.A2(net653),
.A3(net632),
.ZN(net659)
);

INV_X1 c655(
.A(net644),
.ZN(net660)
);

XNOR2_X1 c656(
.A(net642),
.B(net651),
.ZN(net661)
);

NAND3_X2 c657(
.A1(net633),
.A2(net658),
.A3(net661),
.ZN(net662)
);

OR3_X1 c658(
.A1(net436),
.A2(net537),
.A3(net628),
.ZN(net663)
);

AOI221_X2 c659(
.A(net192),
.B1(net655),
.B2(net595),
.C1(net594),
.C2(net607),
.ZN(net664)
);

MUX2_X1 c660(
.A(net589),
.B(net636),
.S(net562),
.Z(net665)
);

DFFRS_X1 c661(
.D(net586),
.RN(net662),
.SN(net609),
.CK(clk),
.Q(net667),
.QN(net666)
);

OAI21_X4 c662(
.A(net351),
.B1(net661),
.B2(net637),
.ZN(net668)
);

NOR4_X4 c663(
.A1(net636),
.A2(net657),
.A3(net654),
.A4(net666),
.ZN(net669)
);

INV_X2 c664(
.A(net11105),
.ZN(net670)
);

INV_X8 c665(
.A(net11145),
.ZN(net671)
);

INV_X16 c666(
.A(net611),
.ZN(net672)
);

OR2_X4 c667(
.A1(net251),
.A2(net650),
.ZN(net673)
);

INV_X32 c668(
.A(net671),
.ZN(net674)
);

INV_X4 c669(
.A(net465),
.ZN(net675)
);

INV_X1 c670(
.A(net648),
.ZN(net676)
);

INV_X2 c671(
.A(net10131),
.ZN(net677)
);

INV_X8 c672(
.A(net673),
.ZN(net678)
);

INV_X16 c673(
.A(net11105),
.ZN(net679)
);

INV_X32 c674(
.A(net611),
.ZN(net680)
);

INV_X4 c675(
.A(net9729),
.ZN(net681)
);

OR2_X1 c676(
.A1(net640),
.A2(net656),
.ZN(net682)
);

INV_X1 c677(
.A(net612),
.ZN(net683)
);

INV_X2 c678(
.A(net10905),
.ZN(net684)
);

INV_X8 c679(
.A(net676),
.ZN(net685)
);

XNOR2_X2 c680(
.A(net658),
.B(net587),
.ZN(net686)
);

INV_X16 c681(
.A(net639),
.ZN(net687)
);

INV_X32 c682(
.A(net365),
.ZN(net688)
);

INV_X4 c683(
.A(net640),
.ZN(net689)
);

INV_X1 c684(
.A(net9793),
.ZN(net690)
);

INV_X2 c685(
.A(net652),
.ZN(net691)
);

AND2_X4 c686(
.A1(net612),
.A2(net10905),
.ZN(net692)
);

INV_X8 c687(
.A(net692),
.ZN(net693)
);

INV_X16 c688(
.A(net671),
.ZN(net694)
);

AND2_X1 c689(
.A1(net645),
.A2(net587),
.ZN(net695)
);

INV_X32 c690(
.A(net587),
.ZN(net696)
);

INV_X4 c691(
.A(net691),
.ZN(net697)
);

INV_X1 c692(
.A(net678),
.ZN(net698)
);

INV_X2 c693(
.A(net524),
.ZN(net699)
);

NAND2_X1 c694(
.A1(net667),
.A2(net672),
.ZN(net700)
);

INV_X8 c695(
.A(net696),
.ZN(net701)
);

INV_X16 c696(
.A(net661),
.ZN(net702)
);

INV_X32 c697(
.A(net692),
.ZN(net703)
);

INV_X4 c698(
.A(net682),
.ZN(net704)
);

INV_X1 c699(
.A(net701),
.ZN(net705)
);

NAND2_X2 c700(
.A1(net677),
.A2(net691),
.ZN(net706)
);

INV_X2 c701(
.A(net690),
.ZN(net707)
);

INV_X8 c702(
.A(net9793),
.ZN(net708)
);

NAND2_X4 c703(
.A1(net697),
.A2(net678),
.ZN(net709)
);

AND2_X2 c704(
.A1(net706),
.A2(net691),
.ZN(net710)
);

INV_X16 c705(
.A(net591),
.ZN(net711)
);

INV_X32 c706(
.A(net687),
.ZN(net712)
);

XOR2_X1 c707(
.A(net705),
.B(net702),
.Z(net713)
);

NOR2_X1 c708(
.A1(net712),
.A2(net674),
.ZN(net714)
);

AOI221_X1 c709(
.A(net657),
.B1(net667),
.B2(net689),
.C1(net708),
.C2(net11144),
.ZN(net715)
);

INV_X4 c710(
.A(net10283),
.ZN(net716)
);

OR2_X2 c711(
.A1(net680),
.A2(net654),
.ZN(net717)
);

INV_X1 c712(
.A(net716),
.ZN(net718)
);

INV_X2 c713(
.A(net706),
.ZN(net719)
);

NOR2_X4 c714(
.A1(net685),
.A2(net709),
.ZN(net720)
);

MUX2_X2 c715(
.A(net718),
.B(net679),
.S(net692),
.Z(net721)
);

NOR2_X2 c716(
.A1(net720),
.A2(net594),
.ZN(net722)
);

XOR2_X2 c717(
.A(net721),
.B(net714),
.Z(net723)
);

INV_X8 c718(
.A(net704),
.ZN(net724)
);

INV_X16 c719(
.A(net715),
.ZN(net725)
);

XNOR2_X1 c720(
.A(net711),
.B(net673),
.ZN(net726)
);

INV_X32 c721(
.A(net675),
.ZN(net727)
);

OR2_X4 c722(
.A1(net700),
.A2(net722),
.ZN(net728)
);

NAND3_X4 c723(
.A1(net434),
.A2(net707),
.A3(net696),
.ZN(net729)
);

OR3_X4 c724(
.A1(net354),
.A2(net717),
.A3(net11146),
.ZN(net730)
);

INV_X4 c725(
.A(net698),
.ZN(net731)
);

AND3_X2 c726(
.A1(net714),
.A2(net620),
.A3(net722),
.ZN(net732)
);

DFFR_X1 c727(
.D(net723),
.RN(net732),
.CK(clk),
.Q(net734),
.QN(net733)
);

SDFFRS_X2 c728(
.D(net627),
.RN(net584),
.SE(net587),
.SI(net710),
.SN(net708),
.CK(clk),
.Q(net736),
.QN(net735)
);

NOR3_X1 c729(
.A1(net717),
.A2(net699),
.A3(net683),
.ZN(net737)
);

INV_X1 c730(
.A(net10120),
.ZN(net738)
);

INV_X2 c731(
.A(net737),
.ZN(net739)
);

OR2_X1 c732(
.A1(net688),
.A2(net730),
.ZN(net740)
);

XNOR2_X2 c733(
.A(net707),
.B(net738),
.ZN(net741)
);

OR3_X2 c734(
.A1(net568),
.A2(net736),
.A3(net674),
.ZN(net742)
);

AND2_X4 c735(
.A1(net672),
.A2(net727),
.ZN(net743)
);

INV_X8 c736(
.A(net713),
.ZN(net744)
);

INV_X16 c737(
.A(net743),
.ZN(net745)
);

INV_X32 c738(
.A(net741),
.ZN(net746)
);

AND2_X1 c739(
.A1(net729),
.A2(net576),
.ZN(net747)
);

OAI21_X2 c740(
.A(net730),
.B1(net747),
.B2(net10930),
.ZN(net748)
);

INV_X4 c741(
.A(net747),
.ZN(net749)
);

OAI21_X1 c742(
.A(net739),
.B1(net712),
.B2(net748),
.ZN(net750)
);

NOR4_X2 c743(
.A1(net749),
.A2(net704),
.A3(net750),
.A4(net715),
.ZN(net751)
);

OAI221_X1 c744(
.A(net742),
.B1(net735),
.B2(net749),
.C1(net687),
.C2(net654),
.ZN(net752)
);

OAI221_X4 c745(
.A(net728),
.B1(net751),
.B2(net744),
.C1(net750),
.C2(net730),
.ZN(net753)
);

NAND2_X1 c746(
.A1(net748),
.A2(net10930),
.ZN(net754)
);

NAND2_X2 c747(
.A1(net337),
.A2(net702),
.ZN(net755)
);

INV_X1 c748(
.A(net9838),
.ZN(net756)
);

INV_X2 c749(
.A(net719),
.ZN(net757)
);

INV_X8 c750(
.A(net654),
.ZN(net758)
);

NAND2_X4 c751(
.A1(net499),
.A2(net757),
.ZN(net759)
);

INV_X16 c752(
.A(net744),
.ZN(net760)
);

AND2_X2 c753(
.A1(net311),
.A2(net710),
.ZN(net761)
);

INV_X32 c754(
.A(net710),
.ZN(net762)
);

INV_X4 c755(
.A(net620),
.ZN(net763)
);

INV_X1 c756(
.A(net651),
.ZN(net764)
);

AOI21_X2 c757(
.A(net278),
.B1(net530),
.B2(net764),
.ZN(net765)
);

INV_X2 c758(
.A(net758),
.ZN(net766)
);

AOI21_X1 c759(
.A(net748),
.B1(net638),
.B2(net686),
.ZN(net767)
);

INV_X8 c760(
.A(net620),
.ZN(net768)
);

INV_X16 c761(
.A(net763),
.ZN(net769)
);

INV_X32 c762(
.A(net734),
.ZN(net770)
);

XOR2_X1 c763(
.A(net70),
.B(net758),
.Z(net771)
);

NOR2_X1 c764(
.A1(net757),
.A2(net708),
.ZN(net772)
);

INV_X4 c765(
.A(net615),
.ZN(net773)
);

INV_X1 c766(
.A(net773),
.ZN(net774)
);

INV_X2 c767(
.A(net11147),
.ZN(net775)
);

INV_X8 c768(
.A(net648),
.ZN(net776)
);

INV_X16 c769(
.A(net724),
.ZN(net777)
);

INV_X32 c770(
.A(net615),
.ZN(net778)
);

INV_X4 c771(
.A(net702),
.ZN(net779)
);

INV_X1 c772(
.A(net770),
.ZN(net780)
);

OR2_X2 c773(
.A1(net57),
.A2(net779),
.ZN(net781)
);

NOR2_X4 c774(
.A1(net768),
.A2(net776),
.ZN(net782)
);

INV_X2 c775(
.A(net764),
.ZN(net783)
);

INV_X8 c776(
.A(net731),
.ZN(net784)
);

INV_X16 c777(
.A(net775),
.ZN(net785)
);

NOR2_X2 c778(
.A1(net761),
.A2(net766),
.ZN(net786)
);

INV_X32 c779(
.A(net9657),
.ZN(net787)
);

XOR2_X2 c780(
.A(net638),
.B(net778),
.Z(net788)
);

XNOR2_X1 c781(
.A(net782),
.B(net719),
.ZN(net789)
);

INV_X4 c782(
.A(net779),
.ZN(net790)
);

OR2_X4 c783(
.A1(net784),
.A2(net785),
.ZN(net791)
);

INV_X1 c784(
.A(net778),
.ZN(net792)
);

AOI21_X4 c785(
.A(net790),
.B1(net781),
.B2(net719),
.ZN(net793)
);

INV_X2 c786(
.A(net774),
.ZN(net794)
);

OR2_X1 c787(
.A1(net638),
.A2(net732),
.ZN(net795)
);

XNOR2_X2 c788(
.A(net709),
.B(net787),
.ZN(net796)
);

AND2_X4 c789(
.A1(net789),
.A2(net10409),
.ZN(net797)
);

INV_X8 c790(
.A(net776),
.ZN(net798)
);

INV_X16 c791(
.A(net794),
.ZN(net799)
);

INV_X32 c792(
.A(out0),
.ZN(net800)
);

INV_X4 c793(
.A(net788),
.ZN(net801)
);

AND2_X1 c794(
.A1(net774),
.A2(net760),
.ZN(net802)
);

NAND2_X1 c795(
.A1(net710),
.A2(net731),
.ZN(net803)
);

INV_X1 c796(
.A(net780),
.ZN(net804)
);

INV_X2 c797(
.A(net790),
.ZN(net805)
);

NAND2_X2 c798(
.A1(net756),
.A2(net778),
.ZN(net806)
);

INV_X8 c799(
.A(net10808),
.ZN(net807)
);

DFFR_X2 c800(
.D(net785),
.RN(net805),
.CK(clk),
.Q(net809),
.QN(net808)
);

INV_X16 c801(
.A(net9657),
.ZN(net810)
);

NAND2_X4 c802(
.A1(net789),
.A2(net794),
.ZN(net811)
);

INV_X32 c803(
.A(net755),
.ZN(net812)
);

AOI211_X4 c804(
.A(net797),
.B(net806),
.C1(net785),
.C2(net807),
.ZN(net813)
);

AND2_X2 c805(
.A1(net763),
.A2(net803),
.ZN(net814)
);

XOR2_X1 c806(
.A(net769),
.B(net648),
.Z(net815)
);

INV_X4 c807(
.A(net10409),
.ZN(net816)
);

INV_X1 c808(
.A(net792),
.ZN(net817)
);

NOR2_X1 c809(
.A1(net703),
.A2(net814),
.ZN(net818)
);

OR2_X2 c810(
.A1(net781),
.A2(net814),
.ZN(net819)
);

NOR4_X1 c811(
.A1(net784),
.A2(net807),
.A3(net781),
.A4(net813),
.ZN(net820)
);

OAI221_X2 c812(
.A(net806),
.B1(net813),
.B2(net648),
.C1(net778),
.C2(net811),
.ZN(net821)
);

NOR2_X4 c813(
.A1(net768),
.A2(net810),
.ZN(net822)
);

INV_X2 c814(
.A(net9893),
.ZN(net823)
);

NOR2_X2 c815(
.A1(net681),
.A2(net811),
.ZN(net824)
);

XOR2_X2 c816(
.A(net791),
.B(net817),
.Z(net825)
);

XNOR2_X1 c817(
.A(net825),
.B(net822),
.ZN(net826)
);

DFFS_X1 c818(
.D(net821),
.SN(net823),
.CK(clk),
.Q(net828),
.QN(net827)
);

OR2_X4 c819(
.A1(net817),
.A2(net702),
.ZN(net829)
);

DFFRS_X2 c820(
.D(net819),
.RN(net826),
.SN(net772),
.CK(clk),
.Q(net831),
.QN(net830)
);

AOI221_X4 c821(
.A(net826),
.B1(net804),
.B2(net790),
.C1(net813),
.C2(net825),
.ZN(net832)
);

AND3_X1 c822(
.A1(net799),
.A2(net814),
.A3(net827),
.ZN(net833)
);

SDFF_X1 c823(
.D(net832),
.SE(net801),
.SI(net792),
.CK(clk),
.Q(net835),
.QN(net834)
);

NAND3_X1 c824(
.A1(net835),
.A2(net654),
.A3(net787),
.ZN(net836)
);

AOI221_X2 c825(
.A(net818),
.B1(net830),
.B2(net833),
.C1(net766),
.C2(net827),
.ZN(net837)
);

AOI211_X2 c826(
.A(net820),
.B(net789),
.C1(net832),
.C2(net813),
.ZN(net838)
);

OR2_X1 c827(
.A1(net824),
.A2(net797),
.ZN(net839)
);

XNOR2_X2 c828(
.A(net829),
.B(net804),
.ZN(net840)
);

SDFFRS_X1 c829(
.D(net840),
.RN(net833),
.SE(net839),
.SI(net813),
.SN(net762),
.CK(clk),
.Q(net842),
.QN(net841)
);

INV_X8 c830(
.A(net813),
.ZN(net843)
);

INV_X16 c831(
.A(net9597),
.ZN(net844)
);

INV_X32 c832(
.A(net459),
.ZN(net845)
);

AND2_X4 c833(
.A1(net581),
.A2(net548),
.ZN(net846)
);

INV_X4 c834(
.A(net351),
.ZN(net847)
);

INV_X1 c835(
.A(net845),
.ZN(net848)
);

INV_X2 c836(
.A(net845),
.ZN(net849)
);

INV_X8 c837(
.A(net847),
.ZN(net850)
);

INV_X16 c838(
.A(net846),
.ZN(net851)
);

AND2_X1 c839(
.A1(net812),
.A2(net811),
.ZN(net852)
);

INV_X32 c840(
.A(net849),
.ZN(net853)
);

INV_X4 c841(
.A(net808),
.ZN(net854)
);

NAND2_X1 c842(
.A1(net854),
.A2(net852),
.ZN(net855)
);

INV_X1 c843(
.A(net10422),
.ZN(net856)
);

INV_X2 c844(
.A(net9597),
.ZN(net857)
);

INV_X8 c845(
.A(net815),
.ZN(net858)
);

NAND2_X2 c846(
.A1(net744),
.A2(net629),
.ZN(net859)
);

SDFF_X2 c847(
.D(net859),
.SE(net815),
.SI(net841),
.CK(clk),
.Q(net861),
.QN(net860)
);

INV_X16 c848(
.A(net847),
.ZN(net862)
);

INV_X32 c849(
.A(net750),
.ZN(net863)
);

DFFRS_X1 c850(
.D(net850),
.RN(net861),
.SN(net760),
.CK(clk),
.Q(net865),
.QN(net864)
);

INV_X4 c851(
.A(net777),
.ZN(net866)
);

NOR3_X4 c852(
.A1(net842),
.A2(net860),
.A3(net776),
.ZN(net867)
);

INV_X1 c853(
.A(net803),
.ZN(net868)
);

INV_X2 c854(
.A(net866),
.ZN(net869)
);

INV_X8 c855(
.A(net856),
.ZN(net870)
);

INV_X16 c856(
.A(net853),
.ZN(net871)
);

INV_X32 c857(
.A(net766),
.ZN(net872)
);

INV_X4 c858(
.A(net812),
.ZN(net873)
);

INV_X1 c859(
.A(net846),
.ZN(net874)
);

NAND2_X4 c860(
.A1(net694),
.A2(net766),
.ZN(net875)
);

AND2_X2 c861(
.A1(net719),
.A2(net767),
.ZN(net876)
);

XOR2_X1 c862(
.A(net856),
.B(net804),
.Z(net877)
);

NOR2_X1 c863(
.A1(net872),
.A2(net813),
.ZN(net878)
);

OR2_X2 c864(
.A1(net514),
.A2(net772),
.ZN(net879)
);

NOR2_X4 c865(
.A1(net877),
.A2(net772),
.ZN(net880)
);

INV_X2 c866(
.A(net871),
.ZN(net881)
);

INV_X8 c867(
.A(net9783),
.ZN(net882)
);

NOR3_X2 c868(
.A1(net848),
.A2(net881),
.A3(net737),
.ZN(net883)
);

AOI22_X1 c869(
.A1(net871),
.A2(net845),
.B1(net488),
.B2(net827),
.ZN(net884)
);

INV_X16 c870(
.A(net737),
.ZN(net885)
);

INV_X32 c871(
.A(net10209),
.ZN(net886)
);

NOR2_X2 c872(
.A1(net870),
.A2(net854),
.ZN(net887)
);

INV_X4 c873(
.A(net858),
.ZN(net888)
);

INV_X1 c874(
.A(net854),
.ZN(net889)
);

XOR2_X2 c875(
.A(net881),
.B(net888),
.Z(net890)
);

INV_X2 c876(
.A(net9783),
.ZN(net891)
);

INV_X8 c877(
.A(net884),
.ZN(net892)
);

AND3_X4 c878(
.A1(net866),
.A2(net888),
.A3(net871),
.ZN(net893)
);

DFFS_X2 c879(
.D(net878),
.SN(net891),
.CK(clk),
.Q(net895),
.QN(net894)
);

NAND3_X2 c880(
.A1(net551),
.A2(net828),
.A3(net629),
.ZN(net896)
);

INV_X16 c881(
.A(net885),
.ZN(net897)
);

INV_X32 c882(
.A(net886),
.ZN(net898)
);

XNOR2_X1 c883(
.A(net892),
.B(net879),
.ZN(net899)
);

OR2_X4 c884(
.A1(net874),
.A2(net842),
.ZN(net900)
);

OR2_X1 c885(
.A1(net898),
.A2(net870),
.ZN(net901)
);

XNOR2_X2 c886(
.A(net844),
.B(net803),
.ZN(net902)
);

INV_X4 c887(
.A(net862),
.ZN(net903)
);

AND2_X4 c888(
.A1(net869),
.A2(net777),
.ZN(net904)
);

INV_X1 c889(
.A(net904),
.ZN(net905)
);

INV_X2 c890(
.A(net857),
.ZN(net906)
);

OR3_X1 c891(
.A1(net868),
.A2(net811),
.A3(net899),
.ZN(net907)
);

MUX2_X1 c892(
.A(net813),
.B(net884),
.S(net871),
.Z(net908)
);

INV_X8 c893(
.A(net901),
.ZN(net909)
);

INV_X16 c894(
.A(net10422),
.ZN(net910)
);

INV_X32 c895(
.A(net9729),
.ZN(net911)
);

INV_X4 c896(
.A(net10130),
.ZN(net912)
);

OAI21_X4 c897(
.A(net907),
.B1(net888),
.B2(net776),
.ZN(net913)
);

AND2_X1 c898(
.A1(net776),
.A2(net879),
.ZN(net914)
);

MUX2_X2 c899(
.A(net861),
.B(net750),
.S(net10856),
.Z(net915)
);

NAND2_X1 c900(
.A1(net906),
.A2(net10856),
.ZN(net916)
);

INV_X1 c901(
.A(net10219),
.ZN(net917)
);

OAI222_X1 c902(
.A1(net911),
.A2(net913),
.B1(net881),
.B2(net888),
.C1(net877),
.C2(net866),
.ZN(net918)
);

NAND2_X2 c903(
.A1(net916),
.A2(net914),
.ZN(net919)
);

INV_X2 c904(
.A(net919),
.ZN(net920)
);

INV_X8 c905(
.A(net11010),
.ZN(net921)
);

NAND3_X4 c906(
.A1(net912),
.A2(net921),
.A3(net887),
.ZN(net922)
);

NAND2_X4 c907(
.A1(net883),
.A2(net804),
.ZN(net923)
);

OR3_X4 c908(
.A1(net917),
.A2(net920),
.A3(net910),
.ZN(net924)
);

AOI221_X1 c909(
.A(net890),
.B1(net865),
.B2(net922),
.C1(net877),
.C2(net551),
.ZN(net925)
);

DFFRS_X2 c910(
.D(net906),
.RN(net921),
.SN(net878),
.CK(clk),
.Q(net927),
.QN(net926)
);

AND3_X2 c911(
.A1(net887),
.A2(net905),
.A3(net10616),
.ZN(net928)
);

AND2_X2 c912(
.A1(net928),
.A2(net10589),
.ZN(net929)
);

INV_X16 c913(
.A(net35),
.ZN(net930)
);

INV_X32 c914(
.A(net9),
.ZN(net931)
);

INV_X4 c915(
.A(net50),
.ZN(net932)
);

INV_X1 c916(
.A(net26),
.ZN(net933)
);

INV_X2 c917(
.A(net47),
.ZN(net934)
);

INV_X8 c918(
.A(net6),
.ZN(net935)
);

INV_X16 c919(
.A(net46),
.ZN(net936)
);

INV_X32 c920(
.A(in23),
.ZN(net937)
);

INV_X4 c921(
.A(in5),
.ZN(net938)
);

INV_X1 c922(
.A(net19),
.ZN(net939)
);

INV_X2 c923(
.A(net6),
.ZN(net940)
);

XOR2_X1 c924(
.A(in12),
.B(net50),
.Z(net941)
);

INV_X8 c925(
.A(net934),
.ZN(net942)
);

INV_X16 c926(
.A(net9670),
.ZN(net943)
);

INV_X32 c927(
.A(net51),
.ZN(net944)
);

INV_X4 c928(
.A(net9670),
.ZN(net945)
);

NOR2_X1 c929(
.A1(in19),
.A2(net940),
.ZN(net946)
);

INV_X1 c930(
.A(net941),
.ZN(net947)
);

INV_X2 c931(
.A(in13),
.ZN(net948)
);

INV_X8 c932(
.A(net941),
.ZN(net949)
);

INV_X16 c933(
.A(net945),
.ZN(net950)
);

INV_X32 c934(
.A(in19),
.ZN(net951)
);

INV_X4 c935(
.A(net948),
.ZN(net952)
);

OR2_X2 c936(
.A1(net947),
.A2(net949),
.ZN(net953)
);

INV_X1 c937(
.A(net945),
.ZN(net954)
);

INV_X2 c938(
.A(net954),
.ZN(net955)
);

NOR2_X4 c939(
.A1(net19),
.A2(net946),
.ZN(net956)
);

INV_X8 c940(
.A(net46),
.ZN(net957)
);

INV_X16 c941(
.A(in7),
.ZN(net958)
);

INV_X32 c942(
.A(net939),
.ZN(net959)
);

INV_X4 c943(
.A(net959),
.ZN(net960)
);

INV_X1 c944(
.A(net938),
.ZN(net961)
);

INV_X2 c945(
.A(net49),
.ZN(net962)
);

INV_X8 c946(
.A(net962),
.ZN(net963)
);

NOR3_X1 c947(
.A1(net949),
.A2(net954),
.A3(net961),
.ZN(net964)
);

INV_X16 c948(
.A(net960),
.ZN(net965)
);

NOR2_X2 c949(
.A1(net51),
.A2(net951),
.ZN(net966)
);

INV_X32 c950(
.A(in9),
.ZN(net967)
);

INV_X4 c951(
.A(net946),
.ZN(net968)
);

INV_X1 c952(
.A(net50),
.ZN(net969)
);

INV_X2 c953(
.A(net967),
.ZN(net970)
);

XOR2_X2 c954(
.A(net933),
.B(net969),
.Z(net971)
);

XNOR2_X1 c955(
.A(net968),
.B(net971),
.ZN(net972)
);

INV_X8 c956(
.A(net963),
.ZN(net973)
);

OR2_X4 c957(
.A1(net964),
.A2(net970),
.ZN(net974)
);

OR2_X1 c958(
.A1(net939),
.A2(net959),
.ZN(net975)
);

OR3_X2 c959(
.A1(net947),
.A2(net962),
.A3(net964),
.ZN(net976)
);

XNOR2_X2 c960(
.A(net958),
.B(net952),
.ZN(net977)
);

INV_X16 c961(
.A(net965),
.ZN(net978)
);

OAI21_X2 c962(
.A(in15),
.B1(net6),
.B2(net937),
.ZN(net979)
);

INV_X32 c963(
.A(net977),
.ZN(net980)
);

AND2_X4 c964(
.A1(net976),
.A2(net6),
.ZN(net981)
);

INV_X4 c965(
.A(net966),
.ZN(net982)
);

AND2_X1 c966(
.A1(net975),
.A2(net965),
.ZN(net983)
);

NAND2_X1 c967(
.A1(net943),
.A2(net978),
.ZN(net984)
);

NAND2_X2 c968(
.A1(net940),
.A2(in23),
.ZN(net985)
);

NAND2_X4 c969(
.A1(net931),
.A2(net980),
.ZN(net986)
);

AND2_X2 c970(
.A1(net973),
.A2(net982),
.ZN(net987)
);

OAI21_X1 c971(
.A(net964),
.B1(net943),
.B2(net954),
.ZN(net988)
);

XOR2_X1 c972(
.A(net934),
.B(net955),
.Z(net989)
);

NOR2_X1 c973(
.A1(net986),
.A2(net977),
.ZN(net990)
);

INV_X1 c974(
.A(net955),
.ZN(net991)
);

INV_X2 c975(
.A(net985),
.ZN(net992)
);

INV_X8 c976(
.A(net990),
.ZN(net993)
);

INV_X16 c977(
.A(in9),
.ZN(net994)
);

AOI21_X2 c978(
.A(net992),
.B1(net993),
.B2(net958),
.ZN(net995)
);

OR2_X2 c979(
.A1(net952),
.A2(net964),
.ZN(net996)
);

INV_X32 c980(
.A(in12),
.ZN(net997)
);

INV_X4 c981(
.A(net982),
.ZN(net998)
);

NOR2_X4 c982(
.A1(net971),
.A2(net973),
.ZN(net999)
);

NOR2_X2 c983(
.A1(net998),
.A2(net990),
.ZN(net1000)
);

XOR2_X2 c984(
.A(net999),
.B(net996),
.Z(net1001)
);

AOI21_X1 c985(
.A(net969),
.B1(net35),
.B2(net989),
.ZN(net1002)
);

XNOR2_X1 c986(
.A(net980),
.B(net959),
.ZN(net1003)
);

OR2_X4 c987(
.A1(net991),
.A2(net10472),
.ZN(net1004)
);

OAI222_X4 c988(
.A1(net992),
.A2(net937),
.B1(net979),
.B2(net1004),
.C1(net961),
.C2(net10472),
.ZN(net1005)
);

OR2_X1 c989(
.A1(net936),
.A2(net10472),
.ZN(net1006)
);

OAI221_X1 c990(
.A(net1000),
.B1(net1005),
.B2(net961),
.C1(net937),
.C2(net10472),
.ZN(net1007)
);

CLKGATETST_X1 c991(
.E(net989),
.SE(net1003),
.CK(clk),
.GCK(net1008)
);

XNOR2_X2 c992(
.A(net1003),
.B(net967),
.ZN(net1009)
);

AND4_X4 c993(
.A1(net1005),
.A2(net1009),
.A3(net1000),
.A4(net1004),
.ZN(net1010)
);

NAND4_X1 c994(
.A1(net1009),
.A2(net996),
.A3(net1000),
.A4(net954),
.ZN(net1011)
);

OR4_X1 c995(
.A1(net984),
.A2(net988),
.A3(net1009),
.A4(net954),
.ZN(net1012)
);

AOI21_X4 c996(
.A(net1071),
.B1(net1069),
.B2(net942),
.ZN(net1013)
);

INV_X1 c997(
.A(net983),
.ZN(net1014)
);

AND2_X4 c998(
.A1(net1073),
.A2(net52),
.ZN(net1015)
);

AND2_X1 c999(
.A1(net108),
.A2(net978),
.ZN(net1016)
);

INV_X2 c1000(
.A(net1058),
.ZN(net1017)
);

INV_X8 c1001(
.A(net117),
.ZN(net1018)
);

NAND2_X1 c1002(
.A1(net1006),
.A2(net1075),
.ZN(net1019)
);

NAND2_X2 c1003(
.A1(net1072),
.A2(net1014),
.ZN(net1020)
);

INV_X16 c1004(
.A(net10536),
.ZN(net1021)
);

INV_X32 c1005(
.A(net1048),
.ZN(net1022)
);

INV_X4 c1006(
.A(net1017),
.ZN(net1023)
);

SDFF_X1 c1007(
.D(net1014),
.SE(net1018),
.SI(net1020),
.CK(clk),
.Q(net1025),
.QN(net1024)
);

INV_X1 c1008(
.A(net972),
.ZN(net1026)
);

INV_X2 c1009(
.A(net938),
.ZN(net1027)
);

AND3_X1 c1010(
.A1(net1021),
.A2(net975),
.A3(net996),
.ZN(net1028)
);

NAND2_X4 c1011(
.A1(net1046),
.A2(net1057),
.ZN(net1029)
);

AND2_X2 c1012(
.A1(net1056),
.A2(net1066),
.ZN(net1030)
);

XOR2_X1 c1013(
.A(net1015),
.B(net1047),
.Z(net1031)
);

NOR2_X1 c1014(
.A1(net1062),
.A2(net1046),
.ZN(net1032)
);

INV_X8 c1015(
.A(net1067),
.ZN(net1033)
);

INV_X16 c1016(
.A(net1057),
.ZN(net1034)
);

OR2_X2 c1017(
.A1(net1033),
.A2(in25),
.ZN(net1035)
);

INV_X32 c1018(
.A(net10399),
.ZN(net1036)
);

SDFF_X2 c1019(
.D(net1018),
.SE(net133),
.SI(net950),
.CK(clk),
.Q(net1038),
.QN(net1037)
);

OAI222_X2 c1020(
.A1(net1036),
.A2(net1030),
.B1(net1059),
.B2(net1053),
.C1(net961),
.C2(net942),
.ZN(net1039)
);

INV_X4 c1021(
.A(net1065),
.ZN(net1040)
);

CLKGATETST_X2 c1022(
.E(net1060),
.SE(net1075),
.CK(clk),
.GCK(net1041)
);

NOR2_X4 c1023(
.A1(net1045),
.A2(net11148),
.ZN(net1042)
);

NOR2_X2 c1024(
.A1(net98),
.A2(net984),
.ZN(net1043)
);

XOR2_X2 c1025(
.A(net1006),
.B(net138),
.Z(net1044)
);

XNOR2_X1 c1026(
.A(net129),
.B(net49),
.ZN(net1045)
);

OR2_X4 c1027(
.A1(net978),
.A2(net122),
.ZN(net1046)
);

OR2_X1 c1028(
.A1(net107),
.A2(net974),
.ZN(net1047)
);

NAND3_X1 c1029(
.A1(net52),
.A2(net138),
.A3(net17),
.ZN(net1048)
);

DFFRS_X1 c1030(
.D(net37),
.RN(net1048),
.SN(net108),
.CK(clk),
.Q(net1050),
.QN(net1049)
);

XNOR2_X2 c1031(
.A(net138),
.B(net136),
.ZN(net1051)
);

INV_X1 c1032(
.A(net9567),
.ZN(net1052)
);

INV_X2 c1033(
.A(net953),
.ZN(net1053)
);

CLKGATETST_X4 c1034(
.E(net112),
.SE(net972),
.CK(clk),
.GCK(net1054)
);

AND2_X4 c1035(
.A1(net1049),
.A2(net52),
.ZN(net1055)
);

INV_X8 c1036(
.A(net62),
.ZN(net1056)
);

CLKGATETST_X8 c1037(
.E(net1044),
.SE(net95),
.CK(clk),
.GCK(net1057)
);

AND2_X1 c1038(
.A1(net974),
.A2(net66),
.ZN(net1058)
);

DFFR_X1 c1039(
.D(net932),
.RN(net133),
.CK(clk),
.Q(net1060),
.QN(net1059)
);

INV_X16 c1040(
.A(net953),
.ZN(net1061)
);

INV_X32 c1041(
.A(net52),
.ZN(net1062)
);

INV_X4 c1042(
.A(net1061),
.ZN(net1063)
);

INV_X1 c1043(
.A(net1044),
.ZN(net1064)
);

INV_X2 c1044(
.A(net1047),
.ZN(net1065)
);

NAND2_X1 c1045(
.A1(net75),
.A2(net70),
.ZN(net1066)
);

INV_X8 c1046(
.A(net9930),
.ZN(net1067)
);

NAND2_X2 c1047(
.A1(net122),
.A2(net1063),
.ZN(net1068)
);

NAND2_X4 c1048(
.A1(net1066),
.A2(net983),
.ZN(net1069)
);

INV_X16 c1049(
.A(net991),
.ZN(net1070)
);

INV_X32 c1050(
.A(net66),
.ZN(net1071)
);

INV_X4 c1051(
.A(net1063),
.ZN(net1072)
);

INV_X1 c1052(
.A(net961),
.ZN(net1073)
);

INV_X2 c1053(
.A(net1062),
.ZN(net1074)
);

AND2_X2 c1054(
.A1(net1068),
.A2(net1047),
.ZN(net1075)
);

INV_X8 c1055(
.A(net1069),
.ZN(net1076)
);

INV_X16 c1056(
.A(net136),
.ZN(net1077)
);

XOR2_X1 c1057(
.A(net1030),
.B(net136),
.Z(net1078)
);

DFFR_X2 c1058(
.D(net1023),
.RN(net954),
.CK(clk),
.Q(net1080),
.QN(net1079)
);

INV_X32 c1059(
.A(net9568),
.ZN(net1081)
);

NOR3_X4 c1060(
.A1(net1040),
.A2(net997),
.A3(net1080),
.ZN(net1082)
);

NOR2_X1 c1061(
.A1(net1050),
.A2(net1042),
.ZN(net1083)
);

OAI22_X1 c1062(
.A1(net1041),
.A2(net1021),
.B1(net1067),
.B2(net1053),
.ZN(net1084)
);

OR2_X2 c1063(
.A1(net1035),
.A2(net961),
.ZN(net1085)
);

NOR2_X4 c1064(
.A1(net122),
.A2(net10536),
.ZN(net1086)
);

DFFS_X1 c1065(
.D(net95),
.SN(net1083),
.CK(clk),
.Q(net1088),
.QN(net1087)
);

NOR2_X2 c1066(
.A1(net1080),
.A2(net10524),
.ZN(net1089)
);

XOR2_X2 c1067(
.A(net1088),
.B(net1024),
.Z(net1090)
);

AND4_X2 c1068(
.A1(net1043),
.A2(net1015),
.A3(net1053),
.A4(net1079),
.ZN(net1091)
);

XNOR2_X1 c1069(
.A(net1080),
.B(net1091),
.ZN(net1092)
);

OR2_X4 c1070(
.A1(net1091),
.A2(net1081),
.ZN(net1093)
);

OAI221_X4 c1071(
.A(net1083),
.B1(net1067),
.B2(net953),
.C1(net1022),
.C2(net1091),
.ZN(net1094)
);

INV_X4 c1072(
.A(net10685),
.ZN(net1095)
);

SDFFS_X1 c1073(
.D(net1090),
.SE(net1094),
.SI(net1079),
.SN(net1091),
.CK(clk),
.Q(net1097),
.QN(net1096)
);

OR2_X1 c1074(
.A1(net133),
.A2(net1095),
.ZN(net1098)
);

XNOR2_X2 c1075(
.A(net1095),
.B(net1032),
.ZN(net1099)
);

AOI222_X1 c1076(
.A1(net1020),
.A2(net1087),
.B1(net1042),
.B2(net1084),
.C1(net1091),
.C2(net11148),
.ZN(net1100)
);

SDFFS_X2 c1077(
.D(net1077),
.SE(net1099),
.SI(net1070),
.SN(net11150),
.CK(clk),
.Q(net1102),
.QN(net1101)
);

AOI222_X4 c1078(
.A1(net972),
.A2(net1101),
.B1(net1091),
.B2(net1070),
.C1(net10536),
.C2(net11150),
.ZN(net1103)
);

INV_X1 c1079(
.A(net9698),
.ZN(net1104)
);

INV_X2 c1080(
.A(net9674),
.ZN(net1105)
);

INV_X8 c1081(
.A(net152),
.ZN(net1106)
);

INV_X16 c1082(
.A(net183),
.ZN(net1107)
);

INV_X32 c1083(
.A(net9674),
.ZN(net1108)
);

INV_X4 c1084(
.A(net1089),
.ZN(net1109)
);

AND2_X4 c1085(
.A1(in25),
.A2(net59),
.ZN(net1110)
);

INV_X1 c1086(
.A(net190),
.ZN(net1111)
);

INV_X2 c1087(
.A(net89),
.ZN(net1112)
);

AND2_X1 c1088(
.A1(net1080),
.A2(net1110),
.ZN(net1113)
);

INV_X8 c1089(
.A(net1034),
.ZN(net1114)
);

INV_X16 c1090(
.A(net1009),
.ZN(net1115)
);

INV_X32 c1091(
.A(net1068),
.ZN(net1116)
);

INV_X4 c1092(
.A(net175),
.ZN(net1117)
);

NOR3_X2 c1093(
.A1(net1117),
.A2(net975),
.A3(net1107),
.ZN(net1118)
);

INV_X1 c1094(
.A(net1052),
.ZN(net1119)
);

INV_X2 c1095(
.A(net9697),
.ZN(net1120)
);

INV_X8 c1096(
.A(net1029),
.ZN(net1121)
);

INV_X16 c1097(
.A(net950),
.ZN(net1122)
);

INV_X32 c1098(
.A(net219),
.ZN(net1123)
);

INV_X4 c1099(
.A(net1031),
.ZN(net1124)
);

INV_X1 c1100(
.A(net214),
.ZN(net1125)
);

INV_X2 c1101(
.A(net1108),
.ZN(net1126)
);

INV_X8 c1102(
.A(net1106),
.ZN(net1127)
);

INV_X16 c1103(
.A(net10172),
.ZN(net1128)
);

NAND2_X1 c1104(
.A1(net1111),
.A2(net11151),
.ZN(net1129)
);

INV_X32 c1105(
.A(net9725),
.ZN(net1130)
);

INV_X4 c1106(
.A(net10636),
.ZN(net1131)
);

INV_X1 c1107(
.A(net9823),
.ZN(net1132)
);

NAND2_X2 c1108(
.A1(net1120),
.A2(net1129),
.ZN(net1133)
);

INV_X2 c1109(
.A(net975),
.ZN(net1134)
);

DFFRS_X2 c1110(
.D(net225),
.RN(net196),
.SN(net932),
.CK(clk),
.Q(net1136),
.QN(net1135)
);

NAND2_X4 c1111(
.A1(net110),
.A2(net1052),
.ZN(net1137)
);

AND2_X2 c1112(
.A1(net1133),
.A2(net1121),
.ZN(net1138)
);

AND3_X4 c1113(
.A1(net1029),
.A2(net1129),
.A3(net11151),
.ZN(net1139)
);

INV_X8 c1114(
.A(net198),
.ZN(net1140)
);

XOR2_X1 c1115(
.A(net1110),
.B(net1132),
.Z(net1141)
);

INV_X16 c1116(
.A(net10633),
.ZN(net1142)
);

INV_X32 c1117(
.A(net161),
.ZN(net1143)
);

SDFF_X1 c1118(
.D(net1143),
.SE(net1138),
.SI(net1121),
.CK(clk),
.Q(net1145),
.QN(net1144)
);

NOR2_X1 c1119(
.A1(net1071),
.A2(net1121),
.ZN(net1146)
);

OR2_X2 c1120(
.A1(net156),
.A2(net1117),
.ZN(net1147)
);

NAND3_X2 c1121(
.A1(net107),
.A2(net1144),
.A3(net1084),
.ZN(net1148)
);

INV_X4 c1122(
.A(net161),
.ZN(net1149)
);

NOR2_X4 c1123(
.A1(net190),
.A2(net89),
.ZN(net1150)
);

DFFS_X2 c1124(
.D(net223),
.SN(net1146),
.CK(clk),
.Q(net1152),
.QN(net1151)
);

NOR2_X2 c1125(
.A1(net1106),
.A2(net1111),
.ZN(net1153)
);

INV_X1 c1126(
.A(net110),
.ZN(net1154)
);

XOR2_X2 c1127(
.A(net68),
.B(net1145),
.Z(net1155)
);

XNOR2_X1 c1128(
.A(net1140),
.B(net1148),
.ZN(net1156)
);

INV_X2 c1129(
.A(net1154),
.ZN(net1157)
);

OR3_X1 c1130(
.A1(net1076),
.A2(net994),
.A3(net11151),
.ZN(net1158)
);

MUX2_X1 c1131(
.A(net1134),
.B(net1150),
.S(net1119),
.Z(net1159)
);

OR2_X4 c1132(
.A1(net189),
.A2(net214),
.ZN(net1160)
);

INV_X8 c1133(
.A(net10810),
.ZN(net1161)
);

OR2_X1 c1134(
.A1(net1131),
.A2(net222),
.ZN(net1162)
);

XNOR2_X2 c1135(
.A(net1162),
.B(net1150),
.ZN(net1163)
);

AND2_X4 c1136(
.A1(net196),
.A2(net1084),
.ZN(net1164)
);

INV_X16 c1137(
.A(net1127),
.ZN(net1165)
);

OAI21_X4 c1138(
.A(net1115),
.B1(net1165),
.B2(net86),
.ZN(net1166)
);

AND2_X1 c1139(
.A1(net59),
.A2(net1141),
.ZN(net1167)
);

NAND2_X1 c1140(
.A1(net1130),
.A2(net1160),
.ZN(net1168)
);

MUX2_X2 c1141(
.A(net1109),
.B(net1114),
.S(net1009),
.Z(net1169)
);

NAND2_X2 c1142(
.A1(net1107),
.A2(net1167),
.ZN(net1170)
);

NAND3_X4 c1143(
.A1(net1120),
.A2(net1160),
.A3(net107),
.ZN(net1171)
);

SDFF_X2 c1144(
.D(net1156),
.SE(net1165),
.SI(net1166),
.CK(clk),
.Q(net1173),
.QN(net1172)
);

OR3_X4 c1145(
.A1(net1171),
.A2(net1162),
.A3(net1170),
.ZN(net1174)
);

NAND2_X4 c1146(
.A1(net1167),
.A2(net1161),
.ZN(net1175)
);

INV_X32 c1147(
.A(net1157),
.ZN(net1176)
);

AND3_X2 c1148(
.A1(net177),
.A2(net1129),
.A3(net1166),
.ZN(net1177)
);

AND2_X2 c1149(
.A1(net1141),
.A2(net1128),
.ZN(net1178)
);

NOR3_X1 c1150(
.A1(net1176),
.A2(net219),
.A3(net1178),
.ZN(net1179)
);

OAI221_X2 c1151(
.A(net1158),
.B1(net1168),
.B2(net1166),
.C1(net942),
.C2(net1179),
.ZN(net1180)
);

OR3_X2 c1152(
.A1(net1166),
.A2(net1122),
.A3(net1151),
.ZN(net1181)
);

OAI21_X2 c1153(
.A(net1168),
.B1(net1179),
.B2(net1115),
.ZN(net1182)
);

OAI21_X1 c1154(
.A(net1152),
.B1(net1179),
.B2(net10868),
.ZN(net1183)
);

XOR2_X1 c1155(
.A(net191),
.B(net10868),
.Z(net1184)
);

NOR2_X1 c1156(
.A1(net1178),
.A2(net1177),
.ZN(net1185)
);

CLKGATETST_X1 c1157(
.E(net1185),
.SE(net189),
.CK(clk),
.GCK(net1186)
);

DFFRS_X1 c1158(
.D(net1184),
.RN(net1179),
.SN(net1185),
.CK(clk),
.Q(net1188),
.QN(net1187)
);

AOI21_X2 c1159(
.A(net1132),
.B1(net1176),
.B2(net1109),
.ZN(net1189)
);

AOI21_X1 c1160(
.A(net1155),
.B1(net1181),
.B2(net1175),
.ZN(net1190)
);

OAI33_X1 c1161(
.A1(net937),
.A2(net1190),
.A3(net1179),
.B1(net1079),
.B2(net1052),
.B3(net10528),
.ZN(net1191)
);

INV_X4 c1162(
.A(net9745),
.ZN(net1192)
);

INV_X1 c1163(
.A(net259),
.ZN(net1193)
);

INV_X2 c1164(
.A(net247),
.ZN(net1194)
);

INV_X8 c1165(
.A(net1122),
.ZN(net1195)
);

INV_X16 c1166(
.A(net994),
.ZN(net1196)
);

INV_X32 c1167(
.A(net10833),
.ZN(net1197)
);

INV_X4 c1168(
.A(net10833),
.ZN(net1198)
);

INV_X1 c1169(
.A(net1195),
.ZN(net1199)
);

INV_X2 c1170(
.A(net1199),
.ZN(net1200)
);

INV_X8 c1171(
.A(net11023),
.ZN(net1201)
);

INV_X16 c1172(
.A(net1181),
.ZN(net1202)
);

OR2_X2 c1173(
.A1(net207),
.A2(net1170),
.ZN(net1203)
);

INV_X32 c1174(
.A(net259),
.ZN(net1204)
);

INV_X4 c1175(
.A(net9983),
.ZN(net1205)
);

INV_X1 c1176(
.A(net1026),
.ZN(net1206)
);

INV_X2 c1177(
.A(net10242),
.ZN(net1207)
);

NOR2_X4 c1178(
.A1(net1084),
.A2(net1070),
.ZN(net1208)
);

NOR2_X2 c1179(
.A1(net1202),
.A2(net1179),
.ZN(net1209)
);

XOR2_X2 c1180(
.A(net1150),
.B(net234),
.Z(net1210)
);

XNOR2_X1 c1181(
.A(net1026),
.B(net1193),
.ZN(net1211)
);

INV_X8 c1182(
.A(net1136),
.ZN(net1212)
);

INV_X16 c1183(
.A(net9984),
.ZN(net1213)
);

INV_X32 c1184(
.A(net248),
.ZN(net1214)
);

INV_X4 c1185(
.A(net10398),
.ZN(net1215)
);

AOI21_X4 c1186(
.A(net1171),
.B1(net1138),
.B2(net1211),
.ZN(net1216)
);

INV_X1 c1187(
.A(net1113),
.ZN(net1217)
);

INV_X2 c1188(
.A(net1205),
.ZN(net1218)
);

OR2_X4 c1189(
.A1(net1137),
.A2(net1197),
.ZN(net1219)
);

AND3_X1 c1190(
.A1(net191),
.A2(net1054),
.A3(net1105),
.ZN(net1220)
);

OR2_X1 c1191(
.A1(net318),
.A2(net1196),
.ZN(net1221)
);

INV_X8 c1192(
.A(net1215),
.ZN(net1222)
);

INV_X16 c1193(
.A(net1215),
.ZN(net1223)
);

INV_X32 c1194(
.A(net1214),
.ZN(net1224)
);

XNOR2_X2 c1195(
.A(net1054),
.B(net57),
.ZN(net1225)
);

AND2_X4 c1196(
.A1(net1198),
.A2(net1207),
.ZN(net1226)
);

AND2_X1 c1197(
.A1(net1217),
.A2(net1226),
.ZN(net1227)
);

INV_X4 c1198(
.A(net1118),
.ZN(net1228)
);

INV_X1 c1199(
.A(net1117),
.ZN(net1229)
);

NAND2_X1 c1200(
.A1(net1192),
.A2(net10869),
.ZN(net1230)
);

NAND2_X2 c1201(
.A1(net1165),
.A2(net1226),
.ZN(net1231)
);

INV_X2 c1202(
.A(net1228),
.ZN(net1232)
);

CLKGATETST_X2 c1203(
.E(net1138),
.SE(net308),
.CK(clk),
.GCK(net1233)
);

INV_X8 c1204(
.A(net9725),
.ZN(net1234)
);

INV_X16 c1205(
.A(net1233),
.ZN(net1235)
);

INV_X32 c1206(
.A(net1206),
.ZN(net1236)
);

NAND2_X4 c1207(
.A1(net932),
.A2(net1226),
.ZN(net1237)
);

NAND3_X1 c1208(
.A1(net1232),
.A2(net1211),
.A3(net1213),
.ZN(net1238)
);

NOR3_X4 c1209(
.A1(net234),
.A2(net1238),
.A3(net1193),
.ZN(net1239)
);

INV_X4 c1210(
.A(net1229),
.ZN(net1240)
);

AND2_X2 c1211(
.A1(net1225),
.A2(net1198),
.ZN(net1241)
);

INV_X1 c1212(
.A(net1218),
.ZN(net1242)
);

AND4_X1 c1213(
.A1(net1160),
.A2(net306),
.A3(net45),
.A4(net1070),
.ZN(net1243)
);

XOR2_X1 c1214(
.A(net1104),
.B(net1229),
.Z(net1244)
);

NOR2_X1 c1215(
.A1(net1231),
.A2(net1237),
.ZN(net1245)
);

INV_X2 c1216(
.A(net10889),
.ZN(net1246)
);

OR2_X2 c1217(
.A1(net1226),
.A2(net1240),
.ZN(net1247)
);

INV_X8 c1218(
.A(net1243),
.ZN(net1248)
);

NOR2_X4 c1219(
.A1(net1202),
.A2(net1231),
.ZN(net1249)
);

NOR2_X2 c1220(
.A1(net1220),
.A2(net1217),
.ZN(net1250)
);

XOR2_X2 c1221(
.A(net1240),
.B(net1226),
.Z(net1251)
);

INV_X16 c1222(
.A(net9992),
.ZN(net1252)
);

XNOR2_X1 c1223(
.A(net1214),
.B(net1237),
.ZN(net1253)
);

OR2_X4 c1224(
.A1(net1227),
.A2(net1228),
.ZN(net1254)
);

NOR3_X2 c1225(
.A1(net1123),
.A2(net305),
.A3(net1254),
.ZN(net1255)
);

AND3_X4 c1226(
.A1(net306),
.A2(net1247),
.A3(net1225),
.ZN(net1256)
);

OR2_X1 c1227(
.A1(net1194),
.A2(net1218),
.ZN(net1257)
);

XNOR2_X2 c1228(
.A(net1250),
.B(net994),
.ZN(net1258)
);

AND2_X4 c1229(
.A1(net1256),
.A2(net10402),
.ZN(net1259)
);

AND2_X1 c1230(
.A1(net1255),
.A2(net1211),
.ZN(net1260)
);

NAND2_X1 c1231(
.A1(net17),
.A2(net1227),
.ZN(net1261)
);

NAND3_X2 c1232(
.A1(net1246),
.A2(net1259),
.A3(net1251),
.ZN(net1262)
);

NAND2_X2 c1233(
.A1(net246),
.A2(net1229),
.ZN(net1263)
);

OR3_X1 c1234(
.A1(net1258),
.A2(net1233),
.A3(net1207),
.ZN(net1264)
);

DFFRS_X2 c1235(
.D(net1238),
.RN(net1214),
.SN(net1202),
.CK(clk),
.Q(net1266),
.QN(net1265)
);

MUX2_X1 c1236(
.A(net1263),
.B(net1250),
.S(net1264),
.Z(net1267)
);

OAI21_X4 c1237(
.A(net1222),
.B1(net1121),
.B2(net10890),
.ZN(net1268)
);

MUX2_X2 c1238(
.A(net1247),
.B(net1241),
.S(net1215),
.Z(net1269)
);

AOI222_X2 c1239(
.A1(net1246),
.A2(net1084),
.B1(net1200),
.B2(net1230),
.C1(net251),
.C2(net11041),
.ZN(net1270)
);

AOI22_X4 c1240(
.A1(net1241),
.A2(net1250),
.B1(net1150),
.B2(net1195),
.ZN(net1271)
);

OAI22_X4 c1241(
.A1(net1269),
.A2(net1238),
.B1(net1264),
.B2(net1233),
.ZN(net1272)
);

OAI222_X1 c1242(
.A1(net296),
.A2(net1242),
.B1(net246),
.B2(net1233),
.C1(net1195),
.C2(net251),
.ZN(net1273)
);

NAND2_X4 c1243(
.A1(net1253),
.A2(net1271),
.ZN(net1274)
);

AND2_X2 c1244(
.A1(net1256),
.A2(net1263),
.ZN(net1275)
);

INV_X32 c1245(
.A(net10825),
.ZN(net1276)
);

INV_X4 c1246(
.A(net331),
.ZN(net1277)
);

INV_X1 c1247(
.A(net1163),
.ZN(net1278)
);

INV_X2 c1248(
.A(net10403),
.ZN(net1279)
);

XOR2_X1 c1249(
.A(net298),
.B(net1147),
.Z(net1280)
);

INV_X8 c1250(
.A(net1211),
.ZN(net1281)
);

INV_X16 c1251(
.A(net1105),
.ZN(net1282)
);

INV_X32 c1252(
.A(net11070),
.ZN(net1283)
);

NOR2_X1 c1253(
.A1(net1279),
.A2(net10637),
.ZN(net1284)
);

INV_X4 c1254(
.A(net9605),
.ZN(net1285)
);

INV_X1 c1255(
.A(net10825),
.ZN(net1286)
);

INV_X2 c1256(
.A(net1281),
.ZN(net1287)
);

OR2_X2 c1257(
.A1(net179),
.A2(net401),
.ZN(net1288)
);

INV_X8 c1258(
.A(net9605),
.ZN(net1289)
);

INV_X16 c1259(
.A(net1285),
.ZN(net1290)
);

INV_X32 c1260(
.A(net1240),
.ZN(net1291)
);

NOR2_X4 c1261(
.A1(net45),
.A2(net1259),
.ZN(net1292)
);

CLKGATETST_X4 c1262(
.E(net396),
.SE(net1177),
.CK(clk),
.GCK(net1293)
);

NAND3_X4 c1263(
.A1(net1242),
.A2(net1200),
.A3(net10728),
.ZN(net1294)
);

INV_X4 c1264(
.A(net1121),
.ZN(net1295)
);

INV_X1 c1265(
.A(net316),
.ZN(net1296)
);

INV_X2 c1266(
.A(net1283),
.ZN(net1297)
);

INV_X8 c1267(
.A(net1122),
.ZN(net1298)
);

INV_X16 c1268(
.A(net1282),
.ZN(net1299)
);

AOI221_X4 c1269(
.A(net220),
.B1(net1298),
.B2(net1195),
.C1(net1070),
.C2(net1230),
.ZN(net1300)
);

INV_X32 c1270(
.A(net262),
.ZN(net1301)
);

INV_X4 c1271(
.A(net1242),
.ZN(net1302)
);

NOR2_X2 c1272(
.A1(net1192),
.A2(net1207),
.ZN(net1303)
);

INV_X1 c1273(
.A(net1142),
.ZN(net1304)
);

INV_X2 c1274(
.A(net1147),
.ZN(net1305)
);

INV_X8 c1275(
.A(net9778),
.ZN(net1306)
);

XOR2_X2 c1276(
.A(net1200),
.B(net10869),
.Z(net1307)
);

INV_X16 c1277(
.A(net382),
.ZN(net1308)
);

INV_X32 c1278(
.A(net1164),
.ZN(net1309)
);

INV_X4 c1279(
.A(net1290),
.ZN(net1310)
);

INV_X1 c1280(
.A(net1303),
.ZN(net1311)
);

SDFFR_X1 c1281(
.D(net1277),
.RN(net1268),
.SE(net1285),
.SI(net401),
.CK(clk),
.Q(net1313),
.QN(net1312)
);

INV_X2 c1282(
.A(net1304),
.ZN(net1314)
);

INV_X8 c1283(
.A(net1311),
.ZN(net1315)
);

XNOR2_X1 c1284(
.A(net1313),
.B(net283),
.ZN(net1316)
);

INV_X16 c1285(
.A(net1284),
.ZN(net1317)
);

OR3_X4 c1286(
.A1(net1309),
.A2(net1211),
.A3(net1298),
.ZN(net1318)
);

INV_X32 c1287(
.A(net1301),
.ZN(net1319)
);

INV_X4 c1288(
.A(net10799),
.ZN(net1320)
);

INV_X1 c1289(
.A(net9761),
.ZN(net1321)
);

INV_X2 c1290(
.A(net10890),
.ZN(net1322)
);

AOI22_X2 c1291(
.A1(net323),
.A2(net1298),
.B1(net1279),
.B2(net10637),
.ZN(net1323)
);

OR2_X4 c1292(
.A1(net1316),
.A2(net1322),
.ZN(net1324)
);

INV_X8 c1293(
.A(net11023),
.ZN(net1325)
);

INV_X16 c1294(
.A(net1302),
.ZN(net1326)
);

INV_X32 c1295(
.A(net1326),
.ZN(net1327)
);

OR2_X1 c1296(
.A1(net1287),
.A2(net1208),
.ZN(net1328)
);

INV_X4 c1297(
.A(net9778),
.ZN(net1329)
);

XNOR2_X2 c1298(
.A(net1310),
.B(net1311),
.ZN(net1330)
);

AND2_X4 c1299(
.A1(net1330),
.A2(net1304),
.ZN(net1331)
);

INV_X1 c1300(
.A(net10717),
.ZN(net1332)
);

AND2_X1 c1301(
.A1(net330),
.A2(net1324),
.ZN(net1333)
);

INV_X2 c1302(
.A(net386),
.ZN(net1334)
);

AND3_X2 c1303(
.A1(net370),
.A2(net1304),
.A3(net10799),
.ZN(net1335)
);

NAND2_X1 c1304(
.A1(net1152),
.A2(net1330),
.ZN(net1336)
);

NAND2_X2 c1305(
.A1(net1278),
.A2(net1332),
.ZN(net1337)
);

NAND2_X4 c1306(
.A1(net1333),
.A2(net1195),
.ZN(net1338)
);

AND2_X2 c1307(
.A1(net1296),
.A2(net1321),
.ZN(net1339)
);

INV_X8 c1308(
.A(net1337),
.ZN(net1340)
);

SDFFR_X2 c1309(
.D(net1294),
.RN(net402),
.SE(net408),
.SI(net1230),
.CK(clk),
.Q(net1342),
.QN(net1341)
);

INV_X16 c1310(
.A(net1323),
.ZN(net1343)
);

INV_X32 c1311(
.A(net10937),
.ZN(net1344)
);

XOR2_X1 c1312(
.A(net363),
.B(net1163),
.Z(net1345)
);

NOR2_X1 c1313(
.A1(net1201),
.A2(net1332),
.ZN(net1346)
);

NOR3_X1 c1314(
.A1(net1344),
.A2(net1339),
.A3(net987),
.ZN(net1347)
);

OR2_X2 c1315(
.A1(net1327),
.A2(net1293),
.ZN(net1348)
);

INV_X4 c1316(
.A(net10811),
.ZN(net1349)
);

NAND4_X4 c1317(
.A1(net1348),
.A2(net1304),
.A3(net1324),
.A4(net10643),
.ZN(net1350)
);

OR3_X2 c1318(
.A1(net1306),
.A2(net1290),
.A3(net1310),
.ZN(net1351)
);

OAI211_X2 c1319(
.A(net1248),
.B(net1195),
.C1(net343),
.C2(net1332),
.ZN(net1352)
);

NOR2_X4 c1320(
.A1(net1312),
.A2(net10955),
.ZN(net1353)
);

OAI21_X2 c1321(
.A(net1349),
.B1(net1350),
.B2(net10955),
.ZN(net1354)
);

NOR2_X2 c1322(
.A1(net1343),
.A2(net1354),
.ZN(net1355)
);

OAI21_X1 c1323(
.A(net1266),
.B1(net1310),
.B2(net10644),
.ZN(net1356)
);

AOI221_X2 c1324(
.A(net1338),
.B1(net1339),
.B2(net1332),
.C1(net1355),
.C2(net1334),
.ZN(net1357)
);

SDFF_X1 c1325(
.D(net1204),
.SE(net1248),
.SI(net1300),
.CK(clk),
.Q(net1359),
.QN(net1358)
);

XOR2_X2 c1326(
.A(net1351),
.B(net1335),
.Z(net1360)
);

AOI21_X2 c1327(
.A(net1357),
.B1(net1358),
.B2(net1360),
.ZN(net1361)
);

INV_X1 c1328(
.A(net9746),
.ZN(net1362)
);

INV_X2 c1329(
.A(net1353),
.ZN(net1363)
);

XNOR2_X1 c1330(
.A(net303),
.B(net416),
.ZN(net1364)
);

INV_X8 c1331(
.A(net10931),
.ZN(net1365)
);

OR2_X4 c1332(
.A1(net1266),
.A2(net1259),
.ZN(net1366)
);

INV_X16 c1333(
.A(net1133),
.ZN(net1367)
);

OR2_X1 c1334(
.A1(net162),
.A2(net1334),
.ZN(net1368)
);

SDFF_X2 c1335(
.D(net301),
.SE(net1208),
.SI(net1295),
.CK(clk),
.Q(net1370),
.QN(net1369)
);

XNOR2_X2 c1336(
.A(net150),
.B(net443),
.ZN(net1371)
);

INV_X32 c1337(
.A(net435),
.ZN(net1372)
);

AND2_X4 c1338(
.A1(net416),
.A2(net320),
.ZN(net1373)
);

AND2_X1 c1339(
.A1(net1371),
.A2(net1298),
.ZN(net1374)
);

INV_X4 c1340(
.A(net493),
.ZN(net1375)
);

NAND2_X1 c1341(
.A1(net1210),
.A2(net1359),
.ZN(net1376)
);

OR4_X2 c1342(
.A1(net424),
.A2(net1376),
.A3(net1317),
.A4(net1354),
.ZN(net1377)
);

INV_X1 c1343(
.A(net1259),
.ZN(net1378)
);

AOI21_X1 c1344(
.A(net1342),
.B1(net1276),
.B2(net442),
.ZN(net1379)
);

INV_X2 c1345(
.A(net432),
.ZN(net1380)
);

INV_X8 c1346(
.A(net449),
.ZN(net1381)
);

NAND2_X2 c1347(
.A1(net1220),
.A2(net1321),
.ZN(net1382)
);

NAND2_X4 c1348(
.A1(net1257),
.A2(net472),
.ZN(net1383)
);

INV_X16 c1349(
.A(net343),
.ZN(net1384)
);

CLKGATETST_X8 c1350(
.E(net1295),
.SE(net476),
.CK(clk),
.GCK(net1385)
);

INV_X32 c1351(
.A(net10362),
.ZN(net1386)
);

INV_X4 c1352(
.A(net1286),
.ZN(net1387)
);

INV_X1 c1353(
.A(net10946),
.ZN(net1388)
);

INV_X2 c1354(
.A(net1376),
.ZN(net1389)
);

AND2_X2 c1355(
.A1(net1265),
.A2(net10740),
.ZN(net1390)
);

INV_X8 c1356(
.A(net1387),
.ZN(net1391)
);

INV_X16 c1357(
.A(net1325),
.ZN(net1392)
);

INV_X32 c1358(
.A(net407),
.ZN(net1393)
);

XOR2_X1 c1359(
.A(net423),
.B(net1383),
.Z(net1394)
);

INV_X4 c1360(
.A(net1373),
.ZN(net1395)
);

NOR2_X1 c1361(
.A1(net1293),
.A2(net1345),
.ZN(net1396)
);

OR2_X2 c1362(
.A1(net453),
.A2(net1392),
.ZN(net1397)
);

NOR2_X4 c1363(
.A1(net480),
.A2(net1394),
.ZN(net1398)
);

NOR2_X2 c1364(
.A1(net427),
.A2(net1341),
.ZN(net1399)
);

INV_X1 c1365(
.A(net10781),
.ZN(net1400)
);

INV_X2 c1366(
.A(net278),
.ZN(net1401)
);

INV_X8 c1367(
.A(net1400),
.ZN(net1402)
);

AOI211_X1 c1368(
.A(net1402),
.B(net1381),
.C1(net455),
.C2(net1070),
.ZN(net1403)
);

AOI21_X4 c1369(
.A(net1362),
.B1(net1375),
.B2(net1385),
.ZN(net1404)
);

INV_X16 c1370(
.A(net10986),
.ZN(net1405)
);

XOR2_X2 c1371(
.A(net472),
.B(net1388),
.Z(net1406)
);

XNOR2_X1 c1372(
.A(net1321),
.B(net435),
.ZN(net1407)
);

INV_X32 c1373(
.A(net1336),
.ZN(net1408)
);

INV_X4 c1374(
.A(net1404),
.ZN(net1409)
);

OR2_X4 c1375(
.A1(net1367),
.A2(net1341),
.ZN(net1410)
);

AND3_X1 c1376(
.A1(net1365),
.A2(net1283),
.A3(net1382),
.ZN(net1411)
);

OR2_X1 c1377(
.A1(net1396),
.A2(net427),
.ZN(net1412)
);

XNOR2_X2 c1378(
.A(net1409),
.B(net424),
.ZN(net1413)
);

INV_X1 c1379(
.A(net1283),
.ZN(net1414)
);

INV_X2 c1380(
.A(net10946),
.ZN(net1415)
);

INV_X8 c1381(
.A(net1377),
.ZN(net1416)
);

INV_X16 c1382(
.A(net1405),
.ZN(net1417)
);

SDFFRS_X2 c1383(
.D(net1378),
.RN(net1387),
.SE(net1400),
.SI(net1208),
.SN(net1392),
.CK(clk),
.Q(net1419),
.QN(net1418)
);

NAND3_X1 c1384(
.A1(net1359),
.A2(net1418),
.A3(net1389),
.ZN(net1420)
);

NAND4_X2 c1385(
.A1(net1420),
.A2(net1390),
.A3(net1408),
.A4(net1380),
.ZN(net1421)
);

DFFRS_X1 c1386(
.D(net1404),
.RN(net450),
.SN(net10644),
.CK(clk),
.Q(net1423),
.QN(net1422)
);

INV_X32 c1387(
.A(net10178),
.ZN(net1424)
);

AND2_X4 c1388(
.A1(net1388),
.A2(net1385),
.ZN(net1425)
);

INV_X4 c1389(
.A(net9888),
.ZN(net1426)
);

INV_X1 c1390(
.A(net9933),
.ZN(net1427)
);

AND2_X1 c1391(
.A1(net1427),
.A2(net1408),
.ZN(net1428)
);

NAND2_X1 c1392(
.A1(net1425),
.A2(net1334),
.ZN(net1429)
);

NOR3_X4 c1393(
.A1(net1397),
.A2(net1354),
.A3(net1422),
.ZN(net1430)
);

NAND2_X2 c1394(
.A1(net1424),
.A2(net10977),
.ZN(net1431)
);

NAND2_X4 c1395(
.A1(net1415),
.A2(net480),
.ZN(net1432)
);

AND2_X2 c1396(
.A1(net1430),
.A2(net1265),
.ZN(net1433)
);

XOR2_X1 c1397(
.A(net1432),
.B(net1355),
.Z(net1434)
);

NOR2_X1 c1398(
.A1(net1413),
.A2(net1388),
.ZN(net1435)
);

OR2_X2 c1399(
.A1(net1417),
.A2(net1411),
.ZN(net1436)
);

NOR3_X2 c1400(
.A1(net1419),
.A2(net1353),
.A3(net10977),
.ZN(net1437)
);

INV_X2 c1401(
.A(net10931),
.ZN(net1438)
);

AOI221_X1 c1402(
.A(net1437),
.B1(net1407),
.B2(net1391),
.C1(net343),
.C2(net1367),
.ZN(net1439)
);

OAI221_X1 c1403(
.A(net1429),
.B1(net1424),
.B2(net1346),
.C1(net1392),
.C2(net1408),
.ZN(net1440)
);

SDFFS_X1 c1404(
.D(net1317),
.SE(net1433),
.SI(net1420),
.SN(net1382),
.CK(clk),
.Q(net1442),
.QN(net1441)
);

OR4_X4 c1405(
.A1(net1399),
.A2(net1436),
.A3(net1441),
.A4(net1298),
.ZN(net1443)
);

INV_X8 c1406(
.A(net11047),
.ZN(net1444)
);

SDFFS_X2 c1407(
.D(net1436),
.SE(net1431),
.SI(net1398),
.SN(net10857),
.CK(clk),
.Q(net1446),
.QN(net1445)
);

AND3_X4 c1408(
.A1(net1346),
.A2(net1444),
.A3(net1425),
.ZN(net1447)
);

NAND3_X2 c1409(
.A1(net1447),
.A2(net276),
.A3(net1437),
.ZN(net1448)
);

OAI222_X4 c1410(
.A1(net1364),
.A2(net1447),
.B1(net1445),
.B2(net1195),
.C1(net1392),
.C2(net10857),
.ZN(net1449)
);

INV_X16 c1411(
.A(net9807),
.ZN(net1450)
);

INV_X32 c1412(
.A(net9621),
.ZN(net1451)
);

NOR2_X4 c1413(
.A1(net543),
.A2(net1380),
.ZN(net1452)
);

NOR2_X2 c1414(
.A1(net392),
.A2(net1384),
.ZN(net1453)
);

OR3_X1 c1415(
.A1(net571),
.A2(net554),
.A3(net1291),
.ZN(net1454)
);

INV_X4 c1416(
.A(net9813),
.ZN(net1455)
);

XOR2_X2 c1417(
.A(net1416),
.B(net10578),
.Z(net1456)
);

XNOR2_X1 c1418(
.A(net1385),
.B(net1345),
.ZN(net1457)
);

INV_X1 c1419(
.A(net11087),
.ZN(net1458)
);

INV_X2 c1420(
.A(net1393),
.ZN(net1459)
);

INV_X8 c1421(
.A(net1419),
.ZN(net1460)
);

OR2_X4 c1422(
.A1(net570),
.A2(net458),
.ZN(net1461)
);

INV_X16 c1423(
.A(net1386),
.ZN(net1462)
);

OAI22_X2 c1424(
.A1(net522),
.A2(net516),
.B1(net368),
.B2(net1392),
.ZN(net1463)
);

MUX2_X1 c1425(
.A(net518),
.B(net500),
.S(net1431),
.Z(net1464)
);

INV_X32 c1426(
.A(net11076),
.ZN(net1465)
);

INV_X4 c1427(
.A(net540),
.ZN(net1466)
);

INV_X1 c1428(
.A(net1389),
.ZN(net1467)
);

INV_X2 c1429(
.A(net11076),
.ZN(net1468)
);

INV_X8 c1430(
.A(net250),
.ZN(net1469)
);

INV_X16 c1431(
.A(net11129),
.ZN(net1470)
);

INV_X32 c1432(
.A(net9761),
.ZN(net1471)
);

OR2_X1 c1433(
.A1(net1468),
.A2(net459),
.ZN(net1472)
);

INV_X4 c1434(
.A(net9765),
.ZN(net1473)
);

XNOR2_X2 c1435(
.A(net1196),
.B(net1276),
.ZN(net1474)
);

INV_X1 c1436(
.A(net1473),
.ZN(net1475)
);

DFFRS_X2 c1437(
.D(net1457),
.RN(net1472),
.SN(net11031),
.CK(clk),
.Q(net1477),
.QN(net1476)
);

INV_X2 c1438(
.A(net533),
.ZN(net1478)
);

INV_X8 c1439(
.A(net1470),
.ZN(net1479)
);

INV_X16 c1440(
.A(net11088),
.ZN(net1480)
);

AND2_X4 c1441(
.A1(net1466),
.A2(net250),
.ZN(net1481)
);

INV_X32 c1442(
.A(net505),
.ZN(net1482)
);

INV_X4 c1443(
.A(net1428),
.ZN(net1483)
);

AND2_X1 c1444(
.A1(net1458),
.A2(net1468),
.ZN(net1484)
);

NAND2_X1 c1445(
.A1(net355),
.A2(net1476),
.ZN(net1485)
);

INV_X1 c1446(
.A(net11075),
.ZN(net1486)
);

OAI21_X4 c1447(
.A(net1482),
.B1(net1462),
.B2(net518),
.ZN(net1487)
);

INV_X2 c1448(
.A(net9807),
.ZN(net1488)
);

MUX2_X2 c1449(
.A(net1453),
.B(net1483),
.S(net530),
.Z(net1489)
);

INV_X8 c1450(
.A(net11002),
.ZN(net1490)
);

OAI211_X4 c1451(
.A(net1276),
.B(net1418),
.C1(net1416),
.C2(net10827),
.ZN(net1491)
);

NAND2_X2 c1452(
.A1(net1451),
.A2(net578),
.ZN(net1492)
);

NAND2_X4 c1453(
.A1(net1442),
.A2(net1469),
.ZN(net1493)
);

INV_X16 c1454(
.A(net1431),
.ZN(net1494)
);

DFFR_X1 c1455(
.D(net1483),
.RN(net517),
.CK(clk),
.Q(net1496),
.QN(net1495)
);

NAND3_X4 c1456(
.A1(net1485),
.A2(net1470),
.A3(net1459),
.ZN(net1497)
);

AND2_X2 c1457(
.A1(net1298),
.A2(net1495),
.ZN(net1498)
);

INV_X32 c1458(
.A(net1390),
.ZN(net1499)
);

XOR2_X1 c1459(
.A(net440),
.B(net1493),
.Z(net1500)
);

INV_X4 c1460(
.A(net11031),
.ZN(net1501)
);

INV_X1 c1461(
.A(net1465),
.ZN(net1502)
);

NOR2_X1 c1462(
.A1(net1474),
.A2(net514),
.ZN(net1503)
);

OR2_X2 c1463(
.A1(net1488),
.A2(net443),
.ZN(net1504)
);

INV_X2 c1464(
.A(net1345),
.ZN(net1505)
);

NOR2_X4 c1465(
.A1(net1499),
.A2(net578),
.ZN(net1506)
);

NOR2_X2 c1466(
.A1(net500),
.A2(net581),
.ZN(net1507)
);

INV_X8 c1467(
.A(net9620),
.ZN(net1508)
);

INV_X16 c1468(
.A(net443),
.ZN(net1509)
);

XOR2_X2 c1469(
.A(net1475),
.B(net1468),
.Z(net1510)
);

OAI222_X2 c1470(
.A1(net554),
.A2(net1482),
.B1(net1510),
.B2(net535),
.C1(net1497),
.C2(net551),
.ZN(net1511)
);

OR3_X4 c1471(
.A1(net1478),
.A2(net578),
.A3(net1369),
.ZN(net1512)
);

XNOR2_X1 c1472(
.A(net1496),
.B(net1434),
.ZN(net1513)
);

AND3_X2 c1473(
.A1(net1186),
.A2(net571),
.A3(net251),
.ZN(net1514)
);

NOR3_X1 c1474(
.A1(net1492),
.A2(net1442),
.A3(net554),
.ZN(net1515)
);

OR2_X4 c1475(
.A1(net1472),
.A2(net1497),
.ZN(net1516)
);

OR3_X2 c1476(
.A1(net517),
.A2(net1504),
.A3(net1508),
.ZN(net1517)
);

OR2_X1 c1477(
.A1(net1516),
.A2(net1497),
.ZN(net1518)
);

OAI21_X2 c1478(
.A(net1477),
.B1(net522),
.B2(net1508),
.ZN(net1519)
);

XNOR2_X2 c1479(
.A(net1490),
.B(net11002),
.ZN(net1520)
);

AND2_X4 c1480(
.A1(net1480),
.A2(net1486),
.ZN(net1521)
);

AND2_X1 c1481(
.A1(net1500),
.A2(net1506),
.ZN(net1522)
);

SDFF_X1 c1482(
.D(net1497),
.SE(net1390),
.SI(net1522),
.CK(clk),
.Q(net1524),
.QN(net1523)
);

OAI21_X1 c1483(
.A(net1496),
.B1(net1523),
.B2(net11069),
.ZN(net1525)
);

AOI222_X1 c1484(
.A1(net1460),
.A2(net1512),
.B1(net1499),
.B2(net1200),
.C1(net1493),
.C2(net578),
.ZN(net1526)
);

SDFF_X2 c1485(
.D(net1366),
.SE(net1477),
.SI(net1522),
.CK(clk),
.Q(net1528),
.QN(net1527)
);

DFFRS_X1 c1486(
.D(net1527),
.RN(net1522),
.SN(net10826),
.CK(clk),
.Q(net1530),
.QN(net1529)
);

DFFRS_X2 c1487(
.D(net1504),
.RN(net1470),
.SN(net1522),
.CK(clk),
.Q(net1532),
.QN(net1531)
);

OAI211_X1 c1488(
.A(net1508),
.B(net1492),
.C1(net1514),
.C2(net1497),
.ZN(net1533)
);

AOI222_X4 c1489(
.A1(net1370),
.A2(net1486),
.B1(net1502),
.B2(net1522),
.C1(net578),
.C2(net551),
.ZN(net1534)
);

AOI21_X2 c1490(
.A(net1514),
.B1(net1531),
.B2(net10815),
.ZN(net1535)
);

SDFF_X1 c1491(
.D(net1501),
.SE(net1522),
.SI(net1535),
.CK(clk),
.Q(net1537),
.QN(net1536)
);

AOI21_X1 c1492(
.A(net1536),
.B1(net1521),
.B2(net10815),
.ZN(net1538)
);

AOI21_X4 c1493(
.A(net1526),
.B1(net1533),
.B2(net11002),
.ZN(net1539)
);

NAND2_X1 c1494(
.A1(net1041),
.A2(net634),
.ZN(net1540)
);

INV_X32 c1495(
.A(net11108),
.ZN(net1541)
);

INV_X4 c1496(
.A(net9782),
.ZN(net1542)
);

NOR4_X4 c1497(
.A1(net573),
.A2(net647),
.A3(net499),
.A4(net650),
.ZN(net1543)
);

INV_X1 c1498(
.A(net1538),
.ZN(net1544)
);

INV_X2 c1499(
.A(net606),
.ZN(net1545)
);

INV_X8 c1500(
.A(net653),
.ZN(net1546)
);

INV_X16 c1501(
.A(net660),
.ZN(net1547)
);

INV_X32 c1502(
.A(net669),
.ZN(net1548)
);

INV_X4 c1503(
.A(net578),
.ZN(net1549)
);

NAND2_X2 c1504(
.A1(net321),
.A2(net618),
.ZN(net1550)
);

INV_X1 c1505(
.A(net1545),
.ZN(net1551)
);

INV_X2 c1506(
.A(net560),
.ZN(net1552)
);

INV_X8 c1507(
.A(net1547),
.ZN(net1553)
);

AND3_X1 c1508(
.A1(net1545),
.A2(net634),
.A3(net1549),
.ZN(net1554)
);

NAND2_X4 c1509(
.A1(net646),
.A2(net339),
.ZN(net1555)
);

AND2_X2 c1510(
.A1(net598),
.A2(net1529),
.ZN(net1556)
);

INV_X16 c1511(
.A(net11108),
.ZN(net1557)
);

INV_X32 c1512(
.A(net1535),
.ZN(net1558)
);

INV_X4 c1513(
.A(net10813),
.ZN(net1559)
);

INV_X1 c1514(
.A(net10813),
.ZN(net1560)
);

INV_X2 c1515(
.A(net11040),
.ZN(net1561)
);

DFFR_X2 c1516(
.D(net1543),
.RN(net455),
.CK(clk),
.Q(net1563),
.QN(net1562)
);

INV_X8 c1517(
.A(net1547),
.ZN(net1564)
);

NAND3_X1 c1518(
.A1(net1554),
.A2(net1562),
.A3(net1540),
.ZN(net1565)
);

XOR2_X1 c1519(
.A(net1307),
.B(net1545),
.Z(net1566)
);

INV_X16 c1520(
.A(net11069),
.ZN(net1567)
);

NOR2_X1 c1521(
.A1(net635),
.A2(net455),
.ZN(net1568)
);

INV_X32 c1522(
.A(net1520),
.ZN(net1569)
);

INV_X4 c1523(
.A(net1530),
.ZN(net1570)
);

DFFS_X1 c1524(
.D(net1556),
.SN(net1563),
.CK(clk),
.Q(net1572),
.QN(net1571)
);

INV_X1 c1525(
.A(net634),
.ZN(net1573)
);

INV_X2 c1526(
.A(net1524),
.ZN(net1574)
);

INV_X8 c1527(
.A(net9782),
.ZN(net1575)
);

OR2_X2 c1528(
.A1(net1550),
.A2(net1427),
.ZN(net1576)
);

NOR2_X4 c1529(
.A1(net1540),
.A2(net605),
.ZN(net1577)
);

NOR2_X2 c1530(
.A1(net662),
.A2(net1354),
.ZN(net1578)
);

XOR2_X2 c1531(
.A(net1541),
.B(net1575),
.Z(net1579)
);

INV_X16 c1532(
.A(net1568),
.ZN(net1580)
);

INV_X32 c1533(
.A(net1565),
.ZN(net1581)
);

INV_X4 c1534(
.A(net625),
.ZN(net1582)
);

INV_X1 c1535(
.A(net368),
.ZN(net1583)
);

XNOR2_X1 c1536(
.A(net1580),
.B(net1509),
.ZN(net1584)
);

OR2_X4 c1537(
.A1(net637),
.A2(net1307),
.ZN(net1585)
);

OR2_X1 c1538(
.A1(net1558),
.A2(net1502),
.ZN(net1586)
);

INV_X2 c1539(
.A(net10084),
.ZN(net1587)
);

XNOR2_X2 c1540(
.A(net1557),
.B(net1584),
.ZN(net1588)
);

AND2_X4 c1541(
.A1(net1509),
.A2(net1558),
.ZN(net1589)
);

AND2_X1 c1542(
.A1(net1578),
.A2(net1581),
.ZN(net1590)
);

NAND2_X1 c1543(
.A1(net1549),
.A2(net1583),
.ZN(net1591)
);

INV_X8 c1544(
.A(net10154),
.ZN(net1592)
);

NOR4_X2 c1545(
.A1(net1573),
.A2(net1583),
.A3(net662),
.A4(net1579),
.ZN(net1593)
);

NAND2_X2 c1546(
.A1(net1559),
.A2(net1585),
.ZN(net1594)
);

OAI221_X4 c1547(
.A(net1406),
.B1(net1589),
.B2(net1570),
.C1(net459),
.C2(net626),
.ZN(net1595)
);

INV_X16 c1548(
.A(net1582),
.ZN(net1596)
);

NAND2_X4 c1549(
.A1(net1462),
.A2(net1530),
.ZN(net1597)
);

AND2_X2 c1550(
.A1(net1577),
.A2(net1545),
.ZN(net1598)
);

INV_X32 c1551(
.A(net1586),
.ZN(net1599)
);

XOR2_X1 c1552(
.A(net1576),
.B(net1406),
.Z(net1600)
);

NOR2_X1 c1553(
.A1(net455),
.A2(net1574),
.ZN(net1601)
);

INV_X4 c1554(
.A(net1555),
.ZN(net1602)
);

OR2_X2 c1555(
.A1(net1546),
.A2(net10772),
.ZN(net1603)
);

NOR2_X4 c1556(
.A1(net605),
.A2(net1570),
.ZN(net1604)
);

NOR2_X2 c1557(
.A1(net1570),
.A2(net1591),
.ZN(net1605)
);

NOR3_X4 c1558(
.A1(net1572),
.A2(net1603),
.A3(net476),
.ZN(net1606)
);

XOR2_X2 c1559(
.A(net1591),
.B(net1577),
.Z(net1607)
);

SDFFR_X1 c1560(
.D(net1597),
.RN(net1526),
.SE(net626),
.SI(net1579),
.CK(clk),
.Q(net1609),
.QN(net1608)
);

NOR3_X2 c1561(
.A1(net1602),
.A2(net1576),
.A3(net1580),
.ZN(net1610)
);

INV_X1 c1562(
.A(net9861),
.ZN(net1611)
);

AND3_X4 c1563(
.A1(net1600),
.A2(net1604),
.A3(net1571),
.ZN(net1612)
);

XNOR2_X1 c1564(
.A(net1592),
.B(net1406),
.ZN(net1613)
);

OR2_X4 c1565(
.A1(net1603),
.A2(net1610),
.ZN(net1614)
);

INV_X2 c1566(
.A(net1605),
.ZN(net1615)
);

SDFFR_X2 c1567(
.D(net1581),
.RN(net1607),
.SE(net1610),
.SI(net1615),
.CK(clk),
.Q(net1617),
.QN(net1616)
);

SDFFRS_X1 c1568(
.D(net1546),
.RN(net1554),
.SE(net1041),
.SI(net1566),
.SN(net1584),
.CK(clk),
.Q(net1619),
.QN(net1618)
);

OR2_X1 c1569(
.A1(net1611),
.A2(net10529),
.ZN(net1620)
);

AOI211_X4 c1570(
.A(net1610),
.B(net1619),
.C1(net1569),
.C2(net1615),
.ZN(net1621)
);

XNOR2_X2 c1571(
.A(net1600),
.B(net10530),
.ZN(net1622)
);

NAND3_X2 c1572(
.A1(net576),
.A2(net1620),
.A3(net10772),
.ZN(net1623)
);

OR3_X1 c1573(
.A1(net1552),
.A2(net1623),
.A3(net1579),
.ZN(net1624)
);

NOR4_X1 c1574(
.A1(net1596),
.A2(net1620),
.A3(net1564),
.A4(net1579),
.ZN(net1625)
);

AND2_X4 c1575(
.A1(net1607),
.A2(net1618),
.ZN(net1626)
);

MUX2_X1 c1576(
.A(net1569),
.B(net1479),
.S(net1624),
.Z(net1627)
);

INV_X8 c1577(
.A(net577),
.ZN(net1628)
);

INV_X16 c1578(
.A(net654),
.ZN(net1629)
);

OAI21_X4 c1579(
.A(net339),
.B1(net1354),
.B2(net1557),
.ZN(net1630)
);

INV_X32 c1580(
.A(net684),
.ZN(net1631)
);

INV_X4 c1581(
.A(net698),
.ZN(net1632)
);

INV_X1 c1582(
.A(net651),
.ZN(net1633)
);

INV_X2 c1583(
.A(net1200),
.ZN(net1634)
);

INV_X8 c1584(
.A(net1634),
.ZN(net1635)
);

AND2_X1 c1585(
.A1(net677),
.A2(net699),
.ZN(net1636)
);

AOI211_X2 c1586(
.A(net350),
.B(net1634),
.C1(net715),
.C2(net1579),
.ZN(net1637)
);

INV_X16 c1587(
.A(net1636),
.ZN(net1638)
);

INV_X32 c1588(
.A(net1619),
.ZN(net1639)
);

INV_X4 c1589(
.A(net727),
.ZN(net1640)
);

INV_X1 c1590(
.A(net592),
.ZN(net1641)
);

INV_X2 c1591(
.A(net1486),
.ZN(net1642)
);

NAND2_X1 c1592(
.A1(net1628),
.A2(net1625),
.ZN(net1643)
);

INV_X8 c1593(
.A(net661),
.ZN(net1644)
);

INV_X16 c1594(
.A(net1557),
.ZN(net1645)
);

NAND2_X2 c1595(
.A1(net1645),
.A2(net1623),
.ZN(net1646)
);

INV_X32 c1596(
.A(net1553),
.ZN(net1647)
);

INV_X4 c1597(
.A(net10964),
.ZN(net1648)
);

INV_X1 c1598(
.A(net1566),
.ZN(net1649)
);

INV_X2 c1599(
.A(net527),
.ZN(net1650)
);

INV_X8 c1600(
.A(net1629),
.ZN(net1651)
);

INV_X16 c1601(
.A(net722),
.ZN(net1652)
);

INV_X32 c1602(
.A(net10964),
.ZN(net1653)
);

INV_X4 c1603(
.A(net1548),
.ZN(net1654)
);

INV_X1 c1604(
.A(net704),
.ZN(net1655)
);

NAND2_X4 c1605(
.A1(net594),
.A2(net722),
.ZN(net1656)
);

MUX2_X2 c1606(
.A(net727),
.B(net686),
.S(net10773),
.Z(net1657)
);

INV_X2 c1607(
.A(net1656),
.ZN(net1658)
);

AND2_X2 c1608(
.A1(net1630),
.A2(net1655),
.ZN(net1659)
);

INV_X8 c1609(
.A(net1628),
.ZN(net1660)
);

INV_X16 c1610(
.A(net1652),
.ZN(net1661)
);

XOR2_X1 c1611(
.A(net1604),
.B(net1631),
.Z(net1662)
);

NOR2_X1 c1612(
.A1(net1592),
.A2(net1635),
.ZN(net1663)
);

OR2_X2 c1613(
.A1(net1544),
.A2(net748),
.ZN(net1664)
);

INV_X32 c1614(
.A(net1634),
.ZN(net1665)
);

INV_X4 c1615(
.A(net535),
.ZN(net1666)
);

NOR2_X4 c1616(
.A1(net1583),
.A2(net1620),
.ZN(net1667)
);

INV_X1 c1617(
.A(net9830),
.ZN(net1668)
);

NOR2_X2 c1618(
.A1(net1639),
.A2(net514),
.ZN(net1669)
);

XOR2_X2 c1619(
.A(net1651),
.B(net1652),
.Z(net1670)
);

INV_X2 c1620(
.A(net11065),
.ZN(net1671)
);

INV_X8 c1621(
.A(net11030),
.ZN(net1672)
);

INV_X16 c1622(
.A(net730),
.ZN(net1673)
);

INV_X32 c1623(
.A(net1644),
.ZN(net1674)
);

INV_X4 c1624(
.A(net9839),
.ZN(net1675)
);

DFFS_X2 c1625(
.D(net1658),
.SN(net1661),
.CK(clk),
.Q(net1677),
.QN(net1676)
);

INV_X1 c1626(
.A(net1632),
.ZN(net1678)
);

XNOR2_X1 c1627(
.A(net1662),
.B(net1663),
.ZN(net1679)
);

NAND3_X4 c1628(
.A1(net1641),
.A2(net1661),
.A3(net751),
.ZN(net1680)
);

OR3_X4 c1629(
.A1(net1649),
.A2(net1666),
.A3(net1678),
.ZN(net1681)
);

OR2_X4 c1630(
.A1(net725),
.A2(net1666),
.ZN(net1682)
);

OR2_X1 c1631(
.A1(net745),
.A2(net1681),
.ZN(net1683)
);

CLKGATETST_X1 c1632(
.E(net1674),
.SE(net1661),
.CK(clk),
.GCK(net1684)
);

XNOR2_X2 c1633(
.A(net1645),
.B(net1631),
.ZN(net1685)
);

INV_X2 c1634(
.A(net10249),
.ZN(net1686)
);

AND2_X4 c1635(
.A1(net1567),
.A2(net1630),
.ZN(net1687)
);

AOI22_X1 c1636(
.A1(net1668),
.A2(net1236),
.B1(net693),
.B2(net654),
.ZN(net1688)
);

AND2_X1 c1637(
.A1(net650),
.A2(net1583),
.ZN(net1689)
);

CLKGATETST_X2 c1638(
.E(net1688),
.SE(net1649),
.CK(clk),
.GCK(net1690)
);

NAND2_X1 c1639(
.A1(net1664),
.A2(net735),
.ZN(net1691)
);

AND3_X2 c1640(
.A1(net1654),
.A2(net1398),
.A3(net746),
.ZN(net1692)
);

INV_X8 c1641(
.A(net10367),
.ZN(net1693)
);

NAND2_X2 c1642(
.A1(net1635),
.A2(net1690),
.ZN(net1694)
);

INV_X16 c1643(
.A(net9842),
.ZN(net1695)
);

AND4_X4 c1644(
.A1(net1633),
.A2(net1693),
.A3(net1678),
.A4(net689),
.ZN(net1696)
);

NAND2_X4 c1645(
.A1(net1663),
.A2(net1562),
.ZN(net1697)
);

AND2_X2 c1646(
.A1(net1693),
.A2(net10995),
.ZN(net1698)
);

INV_X32 c1647(
.A(net1648),
.ZN(net1699)
);

XOR2_X1 c1648(
.A(net1656),
.B(net1681),
.Z(net1700)
);

NOR3_X1 c1649(
.A1(net1697),
.A2(net1686),
.A3(net1699),
.ZN(net1701)
);

NOR2_X1 c1650(
.A1(net1698),
.A2(net1673),
.ZN(net1702)
);

OR3_X2 c1651(
.A1(net1689),
.A2(net1694),
.A3(net650),
.ZN(net1703)
);

OAI21_X2 c1652(
.A(net1637),
.B1(net535),
.B2(net1697),
.ZN(net1704)
);

OAI21_X1 c1653(
.A(net683),
.B1(net1698),
.B2(net1561),
.ZN(net1705)
);

OR2_X2 c1654(
.A1(net1695),
.A2(net1630),
.ZN(net1706)
);

NOR2_X4 c1655(
.A1(net1705),
.A2(net1592),
.ZN(net1707)
);

NOR2_X2 c1656(
.A1(net1699),
.A2(net674),
.ZN(net1708)
);

CLKGATETST_X4 c1657(
.E(net1704),
.SE(net1686),
.CK(clk),
.GCK(net1709)
);

OAI33_X1 c1658(
.A1(net1703),
.A2(net1656),
.A3(net1709),
.B1(net1394),
.B2(net708),
.B3(net1615),
.ZN(net1710)
);

NAND4_X1 c1659(
.A1(net576),
.A2(net1707),
.A3(net1652),
.A4(net1681),
.ZN(net1711)
);

AOI21_X2 c1660(
.A(net794),
.B1(net822),
.B2(net1666),
.ZN(net1712)
);

INV_X4 c1661(
.A(net1496),
.ZN(net1713)
);

XOR2_X2 c1662(
.A(net804),
.B(net11087),
.Z(net1714)
);

XNOR2_X1 c1663(
.A(net1601),
.B(net834),
.ZN(net1715)
);

AOI21_X1 c1664(
.A(net1696),
.B1(net762),
.B2(net11147),
.ZN(net1716)
);

INV_X1 c1665(
.A(net1650),
.ZN(net1717)
);

OR2_X4 c1666(
.A1(net1498),
.A2(net1394),
.ZN(net1718)
);

OR2_X1 c1667(
.A1(net672),
.A2(net767),
.ZN(net1719)
);

INV_X2 c1668(
.A(net10793),
.ZN(net1720)
);

INV_X8 c1669(
.A(net1620),
.ZN(net1721)
);

INV_X16 c1670(
.A(net1563),
.ZN(net1722)
);

INV_X32 c1671(
.A(net1721),
.ZN(net1723)
);

INV_X4 c1672(
.A(net9566),
.ZN(net1724)
);

XNOR2_X2 c1673(
.A(net833),
.B(net1575),
.ZN(net1725)
);

OAI221_X2 c1674(
.A(net738),
.B1(net618),
.B2(net1495),
.C1(net1579),
.C2(net1720),
.ZN(net1726)
);

INV_X1 c1675(
.A(net1561),
.ZN(net1727)
);

SDFF_X2 c1676(
.D(net839),
.SE(net1684),
.SI(net801),
.CK(clk),
.Q(net1729),
.QN(net1728)
);

AND2_X4 c1677(
.A1(net1724),
.A2(net1627),
.ZN(net1730)
);

INV_X2 c1678(
.A(net1674),
.ZN(net1731)
);

INV_X8 c1679(
.A(net1731),
.ZN(net1732)
);

INV_X16 c1680(
.A(net11025),
.ZN(net1733)
);

INV_X32 c1681(
.A(net9758),
.ZN(net1734)
);

INV_X4 c1682(
.A(net783),
.ZN(net1735)
);

SDFFS_X1 c1683(
.D(net1733),
.SE(net1734),
.SI(net759),
.SN(net822),
.CK(clk),
.Q(net1737),
.QN(net1736)
);

DFFRS_X1 c1684(
.D(net759),
.RN(net1734),
.SN(net733),
.CK(clk),
.Q(net1739),
.QN(net1738)
);

AND2_X1 c1685(
.A1(net1722),
.A2(net1694),
.ZN(net1740)
);

INV_X1 c1686(
.A(net758),
.ZN(net1741)
);

INV_X2 c1687(
.A(net796),
.ZN(net1742)
);

AOI21_X4 c1688(
.A(net835),
.B1(net1608),
.B2(net1728),
.ZN(net1743)
);

NAND2_X1 c1689(
.A1(net1742),
.A2(net1708),
.ZN(net1744)
);

NAND2_X2 c1690(
.A1(net1702),
.A2(net814),
.ZN(net1745)
);

NAND2_X4 c1691(
.A1(net1717),
.A2(net822),
.ZN(net1746)
);

INV_X8 c1692(
.A(net1716),
.ZN(net1747)
);

AND2_X2 c1693(
.A1(net1678),
.A2(net1732),
.ZN(net1748)
);

INV_X16 c1694(
.A(net801),
.ZN(net1749)
);

INV_X32 c1695(
.A(net9758),
.ZN(net1750)
);

INV_X4 c1696(
.A(net1723),
.ZN(net1751)
);

XOR2_X1 c1697(
.A(net1747),
.B(net1744),
.Z(net1752)
);

INV_X1 c1698(
.A(net787),
.ZN(net1753)
);

INV_X2 c1699(
.A(net1725),
.ZN(net1754)
);

INV_X8 c1700(
.A(net1734),
.ZN(net1755)
);

INV_X16 c1701(
.A(net1750),
.ZN(net1756)
);

INV_X32 c1702(
.A(net9789),
.ZN(net1757)
);

AOI222_X2 c1703(
.A1(net1679),
.A2(net783),
.B1(net1734),
.B2(net1727),
.C1(net1693),
.C2(net1720),
.ZN(net1758)
);

INV_X4 c1704(
.A(net9789),
.ZN(net1759)
);

INV_X1 c1705(
.A(net9764),
.ZN(net1760)
);

NOR2_X1 c1706(
.A1(net1684),
.A2(net1650),
.ZN(net1761)
);

AOI221_X4 c1707(
.A(net1757),
.B1(net1761),
.B2(net1200),
.C1(net1720),
.C2(net10443),
.ZN(net1762)
);

INV_X2 c1708(
.A(net10817),
.ZN(net1763)
);

INV_X8 c1709(
.A(net1755),
.ZN(net1764)
);

INV_X16 c1710(
.A(net1749),
.ZN(net1765)
);

OR2_X2 c1711(
.A1(net1763),
.A2(net682),
.ZN(net1766)
);

NOR2_X4 c1712(
.A1(net1740),
.A2(net1738),
.ZN(net1767)
);

INV_X32 c1713(
.A(net1726),
.ZN(net1768)
);

INV_X4 c1714(
.A(net810),
.ZN(net1769)
);

NOR2_X2 c1715(
.A1(net1629),
.A2(net1766),
.ZN(net1770)
);

AND3_X1 c1716(
.A1(net736),
.A2(net1757),
.A3(net651),
.ZN(net1771)
);

OR4_X1 c1717(
.A1(net1743),
.A2(net1726),
.A3(net1667),
.A4(net1720),
.ZN(net1772)
);

INV_X1 c1718(
.A(net1764),
.ZN(net1773)
);

NAND3_X1 c1719(
.A1(net1745),
.A2(net1479),
.A3(net10444),
.ZN(net1774)
);

INV_X2 c1720(
.A(net1686),
.ZN(net1775)
);

XOR2_X2 c1721(
.A(net1775),
.B(net1766),
.Z(net1776)
);

INV_X8 c1722(
.A(net1760),
.ZN(net1777)
);

XNOR2_X1 c1723(
.A(net1609),
.B(net1745),
.ZN(net1778)
);

OR2_X4 c1724(
.A1(net1766),
.A2(net1763),
.ZN(net1779)
);

INV_X16 c1725(
.A(net1712),
.ZN(net1780)
);

NOR3_X4 c1726(
.A1(net1713),
.A2(net1763),
.A3(net488),
.ZN(net1781)
);

NOR3_X2 c1727(
.A1(net1751),
.A2(net1780),
.A3(net771),
.ZN(net1782)
);

OR2_X1 c1728(
.A1(net1774),
.A2(net1741),
.ZN(net1783)
);

INV_X32 c1729(
.A(net9764),
.ZN(net1784)
);

XNOR2_X2 c1730(
.A(net1761),
.B(net1781),
.ZN(net1785)
);

AND2_X4 c1731(
.A1(net1772),
.A2(net1769),
.ZN(net1786)
);

AND2_X1 c1732(
.A1(net1770),
.A2(net1601),
.ZN(net1787)
);

INV_X4 c1733(
.A(net9566),
.ZN(net1788)
);

AND3_X4 c1734(
.A1(net1785),
.A2(net1679),
.A3(net1768),
.ZN(net1789)
);

NAND2_X1 c1735(
.A1(net1773),
.A2(net1756),
.ZN(net1790)
);

NAND3_X2 c1736(
.A1(net1746),
.A2(net1790),
.A3(net1765),
.ZN(net1791)
);

NAND2_X2 c1737(
.A1(net1790),
.A2(net1763),
.ZN(net1792)
);

OR3_X1 c1738(
.A1(net1575),
.A2(net1714),
.A3(net651),
.ZN(net1793)
);

NAND2_X4 c1739(
.A1(net786),
.A2(net1782),
.ZN(net1794)
);

MUX2_X1 c1740(
.A(net1781),
.B(net1794),
.S(net1766),
.Z(net1795)
);

OAI21_X4 c1741(
.A(net1788),
.B1(net1789),
.B2(net1794),
.ZN(net1796)
);

INV_X1 c1742(
.A(net10912),
.ZN(net1797)
);

INV_X2 c1743(
.A(net1776),
.ZN(net1798)
);

INV_X8 c1744(
.A(net1762),
.ZN(net1799)
);

AND2_X2 c1745(
.A1(net1765),
.A2(net1615),
.ZN(net1800)
);

INV_X16 c1746(
.A(net1791),
.ZN(net1801)
);

INV_X32 c1747(
.A(net1394),
.ZN(net1802)
);

XOR2_X1 c1748(
.A(net1732),
.B(net928),
.Z(net1803)
);

INV_X4 c1749(
.A(net10257),
.ZN(net1804)
);

INV_X1 c1750(
.A(net1781),
.ZN(net1805)
);

CLKGATETST_X8 c1751(
.E(net929),
.SE(net889),
.CK(clk),
.GCK(net1806)
);

NOR2_X1 c1752(
.A1(net1806),
.A2(net1741),
.ZN(net1807)
);

OR2_X2 c1753(
.A1(net1802),
.A2(net1765),
.ZN(net1808)
);

NOR2_X4 c1754(
.A1(net804),
.A2(net875),
.ZN(net1809)
);

NOR2_X2 c1755(
.A1(net1809),
.A2(net893),
.ZN(net1810)
);

INV_X2 c1756(
.A(net9547),
.ZN(net1811)
);

INV_X8 c1757(
.A(net880),
.ZN(net1812)
);

XOR2_X2 c1758(
.A(net1804),
.B(net807),
.Z(net1813)
);

INV_X16 c1759(
.A(net836),
.ZN(net1814)
);

XNOR2_X1 c1760(
.A(net879),
.B(net1811),
.ZN(net1815)
);

OR2_X4 c1761(
.A1(net809),
.A2(net894),
.ZN(net1816)
);

INV_X32 c1762(
.A(net849),
.ZN(net1817)
);

OR2_X1 c1763(
.A1(net1811),
.A2(net1574),
.ZN(net1818)
);

SDFFS_X2 c1764(
.D(net1799),
.SE(net929),
.SI(net851),
.SN(net877),
.CK(clk),
.Q(net1820),
.QN(net1819)
);

XNOR2_X2 c1765(
.A(net893),
.B(net1693),
.ZN(net1821)
);

INV_X4 c1766(
.A(net1818),
.ZN(net1822)
);

AND2_X4 c1767(
.A1(net873),
.A2(net1801),
.ZN(net1823)
);

AND2_X1 c1768(
.A1(net903),
.A2(net1800),
.ZN(net1824)
);

INV_X1 c1769(
.A(net10716),
.ZN(net1825)
);

NAND2_X1 c1770(
.A1(net1741),
.A2(net1819),
.ZN(net1826)
);

MUX2_X2 c1771(
.A(net694),
.B(net887),
.S(net1801),
.Z(net1827)
);

SDFFR_X1 c1772(
.D(net915),
.RN(net1810),
.SE(net893),
.SI(net1801),
.CK(clk),
.Q(net1829),
.QN(net1828)
);

NAND2_X2 c1773(
.A1(net1715),
.A2(net1816),
.ZN(net1830)
);

NAND2_X4 c1774(
.A1(net874),
.A2(net1806),
.ZN(net1831)
);

AND2_X2 c1775(
.A1(net923),
.A2(net1814),
.ZN(net1832)
);

INV_X2 c1776(
.A(net875),
.ZN(net1833)
);

INV_X8 c1777(
.A(net1694),
.ZN(net1834)
);

XOR2_X1 c1778(
.A(net1815),
.B(net1819),
.Z(net1835)
);

NOR2_X1 c1779(
.A1(net1829),
.A2(net903),
.ZN(net1836)
);

NAND3_X4 c1780(
.A1(net1291),
.A2(net1776),
.A3(net772),
.ZN(net1837)
);

INV_X16 c1781(
.A(net1826),
.ZN(net1838)
);

OR2_X2 c1782(
.A1(net882),
.A2(net922),
.ZN(net1839)
);

INV_X32 c1783(
.A(net9546),
.ZN(net1840)
);

NOR2_X4 c1784(
.A1(net1693),
.A2(net1822),
.ZN(net1841)
);

OR3_X4 c1785(
.A1(net1822),
.A2(net1806),
.A3(net849),
.ZN(net1842)
);

NOR2_X2 c1786(
.A1(net1842),
.A2(net1813),
.ZN(net1843)
);

XOR2_X2 c1787(
.A(net1831),
.B(net836),
.Z(net1844)
);

AND3_X2 c1788(
.A1(net1832),
.A2(net1817),
.A3(net1825),
.ZN(net1845)
);

XNOR2_X1 c1789(
.A(net1837),
.B(net1813),
.ZN(net1846)
);

OR2_X4 c1790(
.A1(net686),
.A2(net1806),
.ZN(net1847)
);

OR2_X1 c1791(
.A1(net877),
.A2(net10817),
.ZN(net1848)
);

XNOR2_X2 c1792(
.A(net1824),
.B(net837),
.ZN(net1849)
);

AND2_X4 c1793(
.A1(net889),
.A2(net10716),
.ZN(net1850)
);

AND2_X1 c1794(
.A1(net1838),
.A2(net1825),
.ZN(net1851)
);

NAND2_X1 c1795(
.A1(net1735),
.A2(net1732),
.ZN(net1852)
);

NOR3_X1 c1796(
.A1(net899),
.A2(net928),
.A3(net1833),
.ZN(net1853)
);

NAND2_X2 c1797(
.A1(net1798),
.A2(net811),
.ZN(net1854)
);

NAND2_X4 c1798(
.A1(net1818),
.A2(net10817),
.ZN(net1855)
);

AND2_X2 c1799(
.A1(net754),
.A2(net1817),
.ZN(net1856)
);

INV_X4 c1800(
.A(net9932),
.ZN(net1857)
);

OAI222_X1 c1801(
.A1(net1821),
.A2(net926),
.B1(net864),
.B2(net851),
.C1(net1801),
.C2(net10762),
.ZN(net1858)
);

XOR2_X1 c1802(
.A(net1851),
.B(net1818),
.Z(net1859)
);

OR3_X2 c1803(
.A1(net1830),
.A2(net1498),
.A3(net1844),
.ZN(net1860)
);

DFFR_X1 c1804(
.D(net1825),
.RN(net1732),
.CK(clk),
.Q(net1862),
.QN(net1861)
);

DFFRS_X2 c1805(
.D(net928),
.RN(net1856),
.SN(net1820),
.CK(clk),
.Q(net1864),
.QN(net1863)
);

OAI21_X2 c1806(
.A(net1854),
.B1(net1842),
.B2(net915),
.ZN(net1865)
);

NOR2_X1 c1807(
.A1(net1498),
.A2(net1848),
.ZN(net1866)
);

OAI21_X1 c1808(
.A(net1859),
.B1(net1791),
.B2(net1861),
.ZN(net1867)
);

SDFF_X1 c1809(
.D(net1867),
.SE(net895),
.SI(net1856),
.CK(clk),
.Q(net1869),
.QN(net1868)
);

AOI21_X2 c1810(
.A(net923),
.B1(net1866),
.B2(net10590),
.ZN(net1870)
);

AOI221_X2 c1811(
.A(net1835),
.B1(net1801),
.B2(net1866),
.C1(net902),
.C2(net864),
.ZN(net1871)
);

AOI21_X1 c1812(
.A(net1855),
.B1(net1868),
.B2(net10971),
.ZN(net1872)
);

AOI21_X4 c1813(
.A(net1870),
.B1(net1864),
.B2(net1857),
.ZN(net1873)
);

OR2_X2 c1814(
.A1(net1870),
.A2(net10766),
.ZN(net1874)
);

OAI22_X1 c1815(
.A1(net1872),
.A2(net1813),
.B1(net1863),
.B2(net864),
.ZN(net1875)
);

NOR2_X4 c1816(
.A1(net1848),
.A2(net1735),
.ZN(net1876)
);

NOR2_X2 c1817(
.A1(net1876),
.A2(net1822),
.ZN(net1877)
);

AND4_X2 c1818(
.A1(net1875),
.A2(net1828),
.A3(net1809),
.A4(net1846),
.ZN(net1878)
);

XOR2_X2 c1819(
.A(net1812),
.B(net11156),
.Z(net1879)
);

AOI221_X1 c1820(
.A(net1800),
.B1(net882),
.B2(net1862),
.C1(net1806),
.C2(net864),
.ZN(net1880)
);

XNOR2_X1 c1821(
.A(net853),
.B(net1844),
.ZN(net1881)
);

OR2_X4 c1822(
.A1(net1880),
.A2(net10616),
.ZN(net1882)
);

AND4_X1 c1823(
.A1(net1866),
.A2(net1878),
.A3(net1857),
.A4(net1816),
.ZN(net1883)
);

SDFF_X2 c1824(
.D(net1883),
.SE(net1880),
.SI(net10971),
.CK(clk),
.Q(net1885),
.QN(net1884)
);

DFFRS_X1 c1825(
.D(net1810),
.RN(net1884),
.SN(net10576),
.CK(clk),
.Q(net1887),
.QN(net1886)
);

INV_X1 c1826(
.A(net944),
.ZN(net1888)
);

INV_X2 c1827(
.A(net1888),
.ZN(net1889)
);

INV_X8 c1828(
.A(net15),
.ZN(net1890)
);

INV_X16 c1829(
.A(net1890),
.ZN(net1891)
);

INV_X32 c1830(
.A(net56),
.ZN(net1892)
);

INV_X4 c1831(
.A(net9683),
.ZN(net1893)
);

DFFR_X2 c1832(
.D(net931),
.RN(net942),
.CK(clk),
.Q(net1895),
.QN(net1894)
);

INV_X1 c1833(
.A(net7),
.ZN(net1896)
);

INV_X2 c1834(
.A(net1889),
.ZN(net1897)
);

INV_X8 c1835(
.A(net1896),
.ZN(net1898)
);

INV_X16 c1836(
.A(net1012),
.ZN(net1899)
);

INV_X32 c1837(
.A(net9682),
.ZN(net1900)
);

INV_X4 c1838(
.A(net981),
.ZN(net1901)
);

INV_X1 c1839(
.A(net995),
.ZN(net1902)
);

OR2_X1 c1840(
.A1(net997),
.A2(net1902),
.ZN(net1903)
);

INV_X2 c1841(
.A(net1900),
.ZN(net1904)
);

XNOR2_X2 c1842(
.A(net966),
.B(net1903),
.ZN(net1905)
);

INV_X8 c1843(
.A(net1895),
.ZN(net1906)
);

AND2_X4 c1844(
.A1(net956),
.A2(net1889),
.ZN(net1907)
);

AND3_X1 c1845(
.A1(net1900),
.A2(net7),
.A3(net10397),
.ZN(net1908)
);

INV_X16 c1846(
.A(net9755),
.ZN(net1909)
);

AND2_X1 c1847(
.A1(net995),
.A2(net1896),
.ZN(net1910)
);

INV_X32 c1848(
.A(net935),
.ZN(net1911)
);

INV_X4 c1849(
.A(net56),
.ZN(net1912)
);

NAND3_X1 c1850(
.A1(net944),
.A2(net1906),
.A3(net984),
.ZN(net1913)
);

INV_X1 c1851(
.A(net1904),
.ZN(net1914)
);

NAND2_X1 c1852(
.A1(net968),
.A2(net1899),
.ZN(net1915)
);

NAND2_X2 c1853(
.A1(net957),
.A2(net1902),
.ZN(net1916)
);

NAND2_X4 c1854(
.A1(net1012),
.A2(net1899),
.ZN(net1917)
);

INV_X2 c1855(
.A(net21),
.ZN(net1918)
);

NOR3_X4 c1856(
.A1(net1912),
.A2(net1910),
.A3(net942),
.ZN(net1919)
);

NOR3_X2 c1857(
.A1(net1902),
.A2(net1000),
.A3(net29),
.ZN(net1920)
);

DFFS_X1 c1858(
.D(net1917),
.SN(net1894),
.CK(clk),
.Q(net1922),
.QN(net1921)
);

AND2_X2 c1859(
.A1(net1899),
.A2(net1921),
.ZN(net1923)
);

INV_X8 c1860(
.A(net9865),
.ZN(net1924)
);

DFFRS_X2 c1861(
.D(net1901),
.RN(net1892),
.SN(net1007),
.CK(clk),
.Q(net1926),
.QN(net1925)
);

INV_X16 c1862(
.A(net1926),
.ZN(net1927)
);

XOR2_X1 c1863(
.A(net1916),
.B(net10397),
.Z(net1928)
);

DFFS_X2 c1864(
.D(net1915),
.SN(net1924),
.CK(clk),
.Q(net1930),
.QN(net1929)
);

CLKGATETST_X1 c1865(
.E(net1889),
.SE(net1923),
.CK(clk),
.GCK(net1931)
);

INV_X32 c1866(
.A(net9866),
.ZN(net1932)
);

NOR2_X1 c1867(
.A1(net1918),
.A2(net1924),
.ZN(net1933)
);

INV_X4 c1868(
.A(net1907),
.ZN(net1934)
);

INV_X1 c1869(
.A(net981),
.ZN(net1935)
);

OR2_X2 c1870(
.A1(net1913),
.A2(net937),
.ZN(net1936)
);

INV_X2 c1871(
.A(net1914),
.ZN(net1937)
);

NOR2_X4 c1872(
.A1(net1893),
.A2(net935),
.ZN(net1938)
);

NOR2_X2 c1873(
.A1(net1910),
.A2(net995),
.ZN(net1939)
);

INV_X8 c1874(
.A(net1888),
.ZN(net1940)
);

CLKGATETST_X2 c1875(
.E(net1917),
.SE(net1004),
.CK(clk),
.GCK(net1941)
);

XOR2_X2 c1876(
.A(net1929),
.B(net1938),
.Z(net1942)
);

XNOR2_X1 c1877(
.A(net1938),
.B(net1904),
.ZN(net1943)
);

AND3_X4 c1878(
.A1(net970),
.A2(net1938),
.A3(net1902),
.ZN(net1944)
);

INV_X16 c1879(
.A(net9738),
.ZN(net1945)
);

CLKGATETST_X4 c1880(
.E(net1940),
.SE(net1944),
.CK(clk),
.GCK(net1946)
);

NAND3_X2 c1881(
.A1(net1924),
.A2(net1904),
.A3(net999),
.ZN(net1947)
);

INV_X32 c1882(
.A(net1943),
.ZN(net1948)
);

CLKGATETST_X8 c1883(
.E(net1935),
.SE(net1921),
.CK(clk),
.GCK(net1949)
);

DFFR_X1 c1884(
.D(net1901),
.RN(net1949),
.CK(clk),
.Q(net1951),
.QN(net1950)
);

OR2_X4 c1885(
.A1(net1948),
.A2(net1913),
.ZN(net1952)
);

INV_X4 c1886(
.A(net1943),
.ZN(net1953)
);

INV_X1 c1887(
.A(net1945),
.ZN(net1954)
);

OR2_X1 c1888(
.A1(net1895),
.A2(net1924),
.ZN(net1955)
);

XNOR2_X2 c1889(
.A(net1911),
.B(net1914),
.ZN(net1956)
);

AND2_X4 c1890(
.A1(net1955),
.A2(net1952),
.ZN(net1957)
);

OR3_X1 c1891(
.A1(net1956),
.A2(net1948),
.A3(net1000),
.ZN(net1958)
);

DFFR_X2 c1892(
.D(net1000),
.RN(net1939),
.CK(clk),
.Q(net1960),
.QN(net1959)
);

DFFS_X1 c1893(
.D(net1939),
.SN(net1932),
.CK(clk),
.Q(net1962),
.QN(net1961)
);

AND2_X1 c1894(
.A1(net1962),
.A2(net1941),
.ZN(net1963)
);

OAI221_X1 c1895(
.A(net960),
.B1(net1958),
.B2(net56),
.C1(net1936),
.C2(net45),
.ZN(net1964)
);

MUX2_X1 c1896(
.A(net1937),
.B(net1925),
.S(net10540),
.Z(net1965)
);

SDFF_X1 c1897(
.D(net1953),
.SE(net1923),
.SI(net1965),
.CK(clk),
.Q(net1967),
.QN(net1966)
);

NAND2_X1 c1898(
.A1(net21),
.A2(net1953),
.ZN(net1968)
);

SDFF_X2 c1899(
.D(net1941),
.SE(net1967),
.SI(net1917),
.CK(clk),
.Q(net1970),
.QN(net1969)
);

OAI21_X4 c1900(
.A(net1969),
.B1(net1942),
.B2(net10665),
.ZN(net1971)
);

DFFS_X2 c1901(
.D(net1892),
.SN(net1935),
.CK(clk),
.Q(net1973),
.QN(net1972)
);

DFFRS_X1 c1902(
.D(net1970),
.RN(net1957),
.SN(net1968),
.CK(clk),
.Q(net1975),
.QN(net1974)
);

NAND2_X2 c1903(
.A1(net1957),
.A2(net1975),
.ZN(net1976)
);

DFFRS_X2 c1904(
.D(net1930),
.RN(net1955),
.SN(net1958),
.CK(clk),
.Q(net1978),
.QN(net1977)
);

NAND2_X4 c1905(
.A1(net1932),
.A2(net10531),
.ZN(net1979)
);

OAI222_X4 c1906(
.A1(in25),
.A2(net1955),
.B1(net1974),
.B2(net942),
.C1(net954),
.C2(net1898),
.ZN(net1980)
);

MUX2_X2 c1907(
.A(net1937),
.B(net1949),
.S(net1979),
.Z(net1981)
);

AOI22_X4 c1908(
.A1(net1975),
.A2(net1971),
.B1(net1981),
.B2(net1920),
.ZN(net1982)
);

INV_X2 c1909(
.A(net1086),
.ZN(net1983)
);

AND2_X2 c1910(
.A1(net45),
.A2(net57),
.ZN(net1984)
);

INV_X8 c1911(
.A(net1938),
.ZN(net1985)
);

XOR2_X1 c1912(
.A(net1979),
.B(net1037),
.Z(net1986)
);

INV_X16 c1913(
.A(net100),
.ZN(net1987)
);

INV_X32 c1914(
.A(net1985),
.ZN(net1988)
);

INV_X4 c1915(
.A(net114),
.ZN(net1989)
);

NOR2_X1 c1916(
.A1(net1986),
.A2(net11149),
.ZN(net1990)
);

INV_X1 c1917(
.A(net9693),
.ZN(net1991)
);

OR2_X2 c1918(
.A1(net954),
.A2(net1979),
.ZN(net1992)
);

INV_X2 c1919(
.A(net9608),
.ZN(net1993)
);

NOR2_X4 c1920(
.A1(net1993),
.A2(net1099),
.ZN(net1994)
);

INV_X8 c1921(
.A(net9608),
.ZN(net1995)
);

INV_X16 c1922(
.A(net1933),
.ZN(net1996)
);

INV_X32 c1923(
.A(net1973),
.ZN(net1997)
);

INV_X4 c1924(
.A(net1987),
.ZN(net1998)
);

INV_X1 c1925(
.A(net1981),
.ZN(net1999)
);

SDFF_X1 c1926(
.D(net100),
.SE(net1075),
.SI(net1990),
.CK(clk),
.Q(net2001),
.QN(net2000)
);

INV_X2 c1927(
.A(net9711),
.ZN(net2002)
);

NOR2_X2 c1928(
.A1(net1963),
.A2(net1997),
.ZN(net2003)
);

XOR2_X2 c1929(
.A(net1075),
.B(net1933),
.Z(net2004)
);

INV_X8 c1930(
.A(net9712),
.ZN(net2005)
);

INV_X16 c1931(
.A(net9712),
.ZN(net2006)
);

XNOR2_X1 c1932(
.A(net1986),
.B(net984),
.ZN(net2007)
);

OR2_X4 c1933(
.A1(net1074),
.A2(net45),
.ZN(net2008)
);

INV_X32 c1934(
.A(net1949),
.ZN(net2009)
);

OR2_X1 c1935(
.A1(net1989),
.A2(net1972),
.ZN(net2010)
);

INV_X4 c1936(
.A(net984),
.ZN(net2011)
);

CLKGATETST_X1 c1937(
.E(net1074),
.SE(net2010),
.CK(clk),
.GCK(net2012)
);

INV_X1 c1938(
.A(net10175),
.ZN(net2013)
);

INV_X2 c1939(
.A(net1996),
.ZN(net2014)
);

INV_X8 c1940(
.A(net9929),
.ZN(net2015)
);

NAND3_X4 c1941(
.A1(net2011),
.A2(net2014),
.A3(net1028),
.ZN(net2016)
);

OR3_X4 c1942(
.A1(net1984),
.A2(net2003),
.A3(net1968),
.ZN(net2017)
);

INV_X16 c1943(
.A(net1991),
.ZN(net2018)
);

INV_X32 c1944(
.A(net1990),
.ZN(net2019)
);

XNOR2_X2 c1945(
.A(net1902),
.B(net86),
.ZN(net2020)
);

SDFF_X2 c1946(
.D(net1997),
.SE(net1916),
.SI(net10532),
.CK(clk),
.Q(net2022),
.QN(net2021)
);

INV_X4 c1947(
.A(net2008),
.ZN(net2023)
);

INV_X1 c1948(
.A(net2016),
.ZN(net2024)
);

INV_X2 c1949(
.A(net1099),
.ZN(net2025)
);

AND2_X4 c1950(
.A1(net2006),
.A2(net1987),
.ZN(net2026)
);

AND3_X2 c1951(
.A1(net978),
.A2(net1985),
.A3(net1963),
.ZN(net2027)
);

INV_X8 c1952(
.A(net2007),
.ZN(net2028)
);

INV_X16 c1953(
.A(net2008),
.ZN(net2029)
);

INV_X32 c1954(
.A(net996),
.ZN(net2030)
);

INV_X4 c1955(
.A(net10006),
.ZN(net2031)
);

INV_X1 c1956(
.A(net2003),
.ZN(net2032)
);

AND2_X1 c1957(
.A1(net2032),
.A2(net10665),
.ZN(net2033)
);

INV_X2 c1958(
.A(net1897),
.ZN(net2034)
);

CLKGATETST_X2 c1959(
.E(net2026),
.SE(net1011),
.CK(clk),
.GCK(net2035)
);

INV_X8 c1960(
.A(net1028),
.ZN(net2036)
);

NOR3_X1 c1961(
.A1(net2031),
.A2(net1074),
.A3(net1949),
.ZN(net2037)
);

CLKGATETST_X4 c1962(
.E(net2014),
.SE(net1920),
.CK(clk),
.GCK(net2038)
);

NAND2_X1 c1963(
.A1(net1988),
.A2(net1997),
.ZN(net2039)
);

NAND2_X2 c1964(
.A1(net2034),
.A2(net2036),
.ZN(net2040)
);

INV_X16 c1965(
.A(net2011),
.ZN(net2041)
);

NAND2_X4 c1966(
.A1(net1997),
.A2(net2035),
.ZN(net2042)
);

AND2_X2 c1967(
.A1(net1086),
.A2(net2000),
.ZN(net2043)
);

XOR2_X1 c1968(
.A(net2035),
.B(net2017),
.Z(net2044)
);

NOR2_X1 c1969(
.A1(net2030),
.A2(net2038),
.ZN(net2045)
);

INV_X32 c1970(
.A(net2017),
.ZN(net2046)
);

INV_X4 c1971(
.A(net10685),
.ZN(net2047)
);

CLKGATETST_X8 c1972(
.E(net2044),
.SE(net1983),
.CK(clk),
.GCK(net2048)
);

OR2_X2 c1973(
.A1(net1983),
.A2(net2038),
.ZN(net2049)
);

OR3_X2 c1974(
.A1(net2020),
.A2(net2048),
.A3(net2043),
.ZN(net2050)
);

NOR2_X4 c1975(
.A1(net2039),
.A2(net2041),
.ZN(net2051)
);

NOR2_X2 c1976(
.A1(net2043),
.A2(net2038),
.ZN(net2052)
);

DFFR_X1 c1977(
.D(net2025),
.RN(net2037),
.CK(clk),
.Q(net2054),
.QN(net2053)
);

OAI21_X2 c1978(
.A(net2009),
.B1(net2049),
.B2(net954),
.ZN(net2055)
);

OAI21_X1 c1979(
.A(net1998),
.B1(net2035),
.B2(net1965),
.ZN(net2056)
);

XOR2_X2 c1980(
.A(net2048),
.B(net10717),
.Z(net2057)
);

OAI222_X2 c1981(
.A1(net2055),
.A2(net2047),
.B1(net1986),
.B2(net1908),
.C1(net1022),
.C2(net1988),
.ZN(net2058)
);

XNOR2_X1 c1982(
.A(net2002),
.B(net2054),
.ZN(net2059)
);

AOI21_X2 c1983(
.A(net2052),
.B1(net2058),
.B2(net2037),
.ZN(net2060)
);

AOI21_X1 c1984(
.A(net1027),
.B1(net2058),
.B2(net2035),
.ZN(net2061)
);

AOI21_X4 c1985(
.A(net120),
.B1(net2053),
.B2(net2056),
.ZN(net2062)
);

OR2_X4 c1986(
.A1(net2061),
.A2(net1096),
.ZN(net2063)
);

OR2_X1 c1987(
.A1(net2042),
.A2(net2056),
.ZN(net2064)
);

XNOR2_X2 c1988(
.A(net2033),
.B(net2063),
.ZN(net2065)
);

AND3_X1 c1989(
.A1(net1984),
.A2(net2064),
.A3(net2056),
.ZN(net2066)
);

NAND3_X1 c1990(
.A1(net2024),
.A2(net2066),
.A3(net11149),
.ZN(net2067)
);

NOR3_X4 c1991(
.A1(net2066),
.A2(net2054),
.A3(net10470),
.ZN(net2068)
);

INV_X1 c1992(
.A(net2149),
.ZN(net2069)
);

INV_X2 c1993(
.A(net1979),
.ZN(net2070)
);

INV_X8 c1994(
.A(net1126),
.ZN(net2071)
);

INV_X16 c1995(
.A(net2154),
.ZN(net2072)
);

DFFR_X2 c1996(
.D(net2144),
.RN(net1128),
.CK(clk),
.Q(net2074),
.QN(net2073)
);

INV_X32 c1997(
.A(net1145),
.ZN(net2075)
);

INV_X4 c1998(
.A(net10346),
.ZN(net2076)
);

AND2_X4 c1999(
.A1(net2073),
.A2(net10629),
.ZN(net2077)
);

INV_X1 c2000(
.A(net1173),
.ZN(net2078)
);

NOR3_X2 c2001(
.A1(net2078),
.A2(net2070),
.A3(net1936),
.ZN(net2079)
);

AND2_X1 c2002(
.A1(net2076),
.A2(net2137),
.ZN(net2080)
);

NAND2_X1 c2003(
.A1(net2079),
.A2(net207),
.ZN(net2081)
);

INV_X2 c2004(
.A(net9565),
.ZN(net2082)
);

INV_X8 c2005(
.A(net9565),
.ZN(net2083)
);

OAI221_X4 c2006(
.A(net1112),
.B1(net1146),
.B2(net2075),
.C1(net2129),
.C2(net185),
.ZN(net2084)
);

NAND2_X2 c2007(
.A1(net2154),
.A2(net2149),
.ZN(net2085)
);

INV_X16 c2008(
.A(net2069),
.ZN(net2086)
);

INV_X32 c2009(
.A(net9711),
.ZN(net2087)
);

NAND2_X4 c2010(
.A1(net2080),
.A2(net2087),
.ZN(net2088)
);

OAI221_X2 c2011(
.A(net2086),
.B1(net114),
.B2(net229),
.C1(net1084),
.C2(net2129),
.ZN(net2089)
);

AND2_X2 c2012(
.A1(net2083),
.A2(net1968),
.ZN(net2090)
);

AND3_X4 c2013(
.A1(net2070),
.A2(net1125),
.A3(net1927),
.ZN(net2091)
);

XOR2_X1 c2014(
.A(net2085),
.B(net2077),
.Z(net2092)
);

NOR2_X1 c2015(
.A1(net2134),
.A2(net2087),
.ZN(net2093)
);

NAND3_X2 c2016(
.A1(net2059),
.A2(net2085),
.A3(net1149),
.ZN(net2094)
);

INV_X4 c2017(
.A(net10048),
.ZN(net2095)
);

OR2_X2 c2018(
.A1(net2141),
.A2(net1965),
.ZN(net2096)
);

OR3_X1 c2019(
.A1(net2092),
.A2(net2080),
.A3(net1085),
.ZN(net2097)
);

NOR2_X4 c2020(
.A1(net2087),
.A2(net2154),
.ZN(net2098)
);

NOR2_X2 c2021(
.A1(net1161),
.A2(net2078),
.ZN(net2099)
);

XOR2_X2 c2022(
.A(net2096),
.B(net2142),
.Z(net2100)
);

INV_X1 c2023(
.A(net2088),
.ZN(net2101)
);

INV_X2 c2024(
.A(net2101),
.ZN(net2102)
);

XNOR2_X1 c2025(
.A(net2089),
.B(net2095),
.ZN(net2103)
);

MUX2_X1 c2026(
.A(net2091),
.B(net2096),
.S(net10806),
.Z(net2104)
);

OR2_X4 c2027(
.A1(net2028),
.A2(net1169),
.ZN(net2105)
);

OAI21_X4 c2028(
.A(net1128),
.B1(net2096),
.B2(net2142),
.ZN(net2106)
);

INV_X8 c2029(
.A(net2099),
.ZN(net2107)
);

INV_X16 c2030(
.A(net2074),
.ZN(net2108)
);

OR2_X1 c2031(
.A1(net2150),
.A2(net2080),
.ZN(net2109)
);

INV_X32 c2032(
.A(net9955),
.ZN(net2110)
);

MUX2_X2 c2033(
.A(net2091),
.B(net2088),
.S(net1034),
.Z(net2111)
);

INV_X4 c2034(
.A(net9786),
.ZN(net2112)
);

DFFRS_X1 c2035(
.D(net2105),
.RN(net2107),
.SN(net1161),
.CK(clk),
.Q(net2114),
.QN(net2113)
);

NAND3_X4 c2036(
.A1(net2077),
.A2(net2109),
.A3(net2147),
.ZN(net2115)
);

OAI22_X4 c2037(
.A1(net1119),
.A2(net2114),
.B1(net2097),
.B2(net2147),
.ZN(net2116)
);

XNOR2_X2 c2038(
.A(net2100),
.B(net2114),
.ZN(net2117)
);

OR3_X4 c2039(
.A1(net2106),
.A2(net2074),
.A3(net2012),
.ZN(net2118)
);

AND2_X4 c2040(
.A1(net207),
.A2(net2109),
.ZN(net2119)
);

AND3_X2 c2041(
.A1(net1085),
.A2(net2069),
.A3(net11070),
.ZN(net2120)
);

NOR3_X1 c2042(
.A1(net2098),
.A2(net57),
.A3(net10975),
.ZN(net2121)
);

OR3_X2 c2043(
.A1(net2104),
.A2(net2120),
.A3(net10975),
.ZN(net2122)
);

SDFFRS_X2 c2044(
.D(net2082),
.RN(net2111),
.SE(net1934),
.SI(net1174),
.SN(net1091),
.CK(clk),
.Q(net2124),
.QN(net2123)
);

AOI22_X2 c2045(
.A1(net2108),
.A2(net2146),
.B1(net2123),
.B2(net2121),
.ZN(net2125)
);

AND2_X1 c2046(
.A1(net2102),
.A2(net2124),
.ZN(net2126)
);

AOI221_X4 c2047(
.A(net2124),
.B1(net2089),
.B2(net1187),
.C1(net2126),
.C2(net120),
.ZN(net2127)
);

AOI221_X2 c2048(
.A(net2097),
.B1(net1186),
.B2(net2123),
.C1(net2126),
.C2(net1988),
.ZN(net2128)
);

INV_X1 c2049(
.A(net1134),
.ZN(net2129)
);

OAI21_X2 c2050(
.A(net2065),
.B1(net1153),
.B2(net1891),
.ZN(net2130)
);

INV_X2 c2051(
.A(net9864),
.ZN(net2131)
);

NAND2_X1 c2052(
.A1(net1111),
.A2(net207),
.ZN(net2132)
);

INV_X8 c2053(
.A(net9823),
.ZN(net2133)
);

INV_X16 c2054(
.A(net1188),
.ZN(net2134)
);

INV_X32 c2055(
.A(net11084),
.ZN(net2135)
);

OAI21_X1 c2056(
.A(net1146),
.B1(net1189),
.B2(net1128),
.ZN(net2136)
);

INV_X4 c2057(
.A(net1143),
.ZN(net2137)
);

AOI221_X1 c2058(
.A(net206),
.B1(net1936),
.B2(net2047),
.C1(net1144),
.C2(net2137),
.ZN(net2138)
);

INV_X1 c2059(
.A(net2137),
.ZN(net2139)
);

NAND2_X2 c2060(
.A1(net1091),
.A2(net1112),
.ZN(net2140)
);

NAND2_X4 c2061(
.A1(net1053),
.A2(net2137),
.ZN(net2141)
);

AND2_X2 c2062(
.A1(net1175),
.A2(net2129),
.ZN(net2142)
);

AOI21_X2 c2063(
.A(net86),
.B1(net1172),
.B2(net2139),
.ZN(net2143)
);

XOR2_X1 c2064(
.A(net2142),
.B(net2032),
.Z(net2144)
);

INV_X2 c2065(
.A(net2143),
.ZN(net2145)
);

NOR2_X1 c2066(
.A1(net2143),
.A2(net1126),
.ZN(net2146)
);

OR2_X2 c2067(
.A1(net2133),
.A2(net1965),
.ZN(net2147)
);

NOR2_X4 c2068(
.A1(net1148),
.A2(net2145),
.ZN(net2148)
);

INV_X8 c2069(
.A(net9700),
.ZN(net2149)
);

INV_X16 c2070(
.A(net2145),
.ZN(net2150)
);

NOR2_X2 c2071(
.A1(net2129),
.A2(net2132),
.ZN(net2151)
);

AOI21_X1 c2072(
.A(net1149),
.B1(net1965),
.B2(net1979),
.ZN(net2152)
);

INV_X32 c2073(
.A(net10129),
.ZN(net2153)
);

INV_X4 c2074(
.A(net10047),
.ZN(net2154)
);

INV_X1 c2075(
.A(net10739),
.ZN(net2155)
);

INV_X2 c2076(
.A(net230),
.ZN(net2156)
);

INV_X8 c2077(
.A(net10927),
.ZN(net2157)
);

XOR2_X2 c2078(
.A(net1246),
.B(net1135),
.Z(net2158)
);

XNOR2_X1 c2079(
.A(net2158),
.B(net2112),
.ZN(net2159)
);

INV_X16 c2080(
.A(net307),
.ZN(net2160)
);

OR2_X4 c2081(
.A1(net1051),
.A2(net1270),
.ZN(net2161)
);

INV_X32 c2082(
.A(net2078),
.ZN(net2162)
);

INV_X4 c2083(
.A(net1219),
.ZN(net2163)
);

INV_X1 c2084(
.A(net1241),
.ZN(net2164)
);

AOI21_X4 c2085(
.A(net2072),
.B1(net2012),
.B2(net2107),
.ZN(net2165)
);

OR2_X1 c2086(
.A1(net1137),
.A2(net1898),
.ZN(net2166)
);

INV_X2 c2087(
.A(net2162),
.ZN(net2167)
);

INV_X8 c2088(
.A(net2158),
.ZN(net2168)
);

INV_X16 c2089(
.A(net2120),
.ZN(net2169)
);

INV_X32 c2090(
.A(net1170),
.ZN(net2170)
);

INV_X4 c2091(
.A(net1273),
.ZN(net2171)
);

XNOR2_X2 c2092(
.A(net1244),
.B(net2155),
.ZN(net2172)
);

INV_X1 c2093(
.A(net2160),
.ZN(net2173)
);

INV_X2 c2094(
.A(net2012),
.ZN(net2174)
);

INV_X8 c2095(
.A(net10174),
.ZN(net2175)
);

INV_X16 c2096(
.A(net10927),
.ZN(net2176)
);

DFFRS_X2 c2097(
.D(net1254),
.RN(net2126),
.SN(net310),
.CK(clk),
.Q(net2178),
.QN(net2177)
);

AND2_X4 c2098(
.A1(net2071),
.A2(net70),
.ZN(net2179)
);

DFFS_X1 c2099(
.D(net1189),
.SN(net2137),
.CK(clk),
.Q(net2181),
.QN(net2180)
);

AND2_X1 c2100(
.A1(net2173),
.A2(net2000),
.ZN(net2182)
);

INV_X32 c2101(
.A(net2075),
.ZN(net2183)
);

INV_X4 c2102(
.A(net2163),
.ZN(net2184)
);

NAND2_X1 c2103(
.A1(net1275),
.A2(net2169),
.ZN(net2185)
);

INV_X1 c2104(
.A(net2179),
.ZN(net2186)
);

AOI222_X1 c2105(
.A1(net2186),
.A2(net2173),
.B1(net2167),
.B2(net2075),
.C1(net1208),
.C2(net1200),
.ZN(net2187)
);

INV_X2 c2106(
.A(net1261),
.ZN(net2188)
);

NAND2_X2 c2107(
.A1(net2185),
.A2(net10739),
.ZN(net2189)
);

NAND2_X4 c2108(
.A1(net1213),
.A2(net1070),
.ZN(net2190)
);

AND2_X2 c2109(
.A1(net1891),
.A2(net2156),
.ZN(net2191)
);

XOR2_X1 c2110(
.A(net2183),
.B(net2170),
.Z(net2192)
);

NOR2_X1 c2111(
.A1(net2169),
.A2(net2018),
.ZN(net2193)
);

OR2_X2 c2112(
.A1(net2193),
.A2(net2180),
.ZN(net2194)
);

INV_X8 c2113(
.A(net10889),
.ZN(net2195)
);

AND3_X1 c2114(
.A1(net2184),
.A2(net2174),
.A3(net2126),
.ZN(net2196)
);

INV_X16 c2115(
.A(net9730),
.ZN(net2197)
);

INV_X32 c2116(
.A(net10841),
.ZN(net2198)
);

NOR2_X4 c2117(
.A1(net2131),
.A2(net307),
.ZN(net2199)
);

NOR2_X2 c2118(
.A1(net2197),
.A2(net2191),
.ZN(net2200)
);

NAND3_X1 c2119(
.A1(net2018),
.A2(net1934),
.A3(net10633),
.ZN(net2201)
);

INV_X4 c2120(
.A(net2175),
.ZN(net2202)
);

INV_X1 c2121(
.A(net2168),
.ZN(net2203)
);

INV_X2 c2122(
.A(net2156),
.ZN(net2204)
);

XOR2_X2 c2123(
.A(net1223),
.B(net2203),
.Z(net2205)
);

NOR3_X4 c2124(
.A1(net247),
.A2(net1223),
.A3(net307),
.ZN(net2206)
);

NAND4_X4 c2125(
.A1(net2187),
.A2(net2176),
.A3(net1246),
.A4(net1988),
.ZN(net2207)
);

XNOR2_X1 c2126(
.A(net2206),
.B(net10740),
.ZN(net2208)
);

OAI211_X2 c2127(
.A(net308),
.B(net2203),
.C1(net2176),
.C2(net2160),
.ZN(net2209)
);

OR2_X4 c2128(
.A1(net2200),
.A2(net2160),
.ZN(net2210)
);

SDFF_X1 c2129(
.D(net1224),
.SE(net2187),
.SI(net2206),
.CK(clk),
.Q(net2212),
.QN(net2211)
);

INV_X8 c2130(
.A(net10974),
.ZN(net2213)
);

INV_X16 c2131(
.A(net10658),
.ZN(net2214)
);

DFFS_X2 c2132(
.D(net2212),
.SN(net1179),
.CK(clk),
.Q(net2216),
.QN(net2215)
);

OR2_X1 c2133(
.A1(net2213),
.A2(net2163),
.ZN(net2217)
);

XNOR2_X2 c2134(
.A(net2194),
.B(net2208),
.ZN(net2218)
);

OR4_X2 c2135(
.A1(net2178),
.A2(net2205),
.A3(net1245),
.A4(net2208),
.ZN(net2219)
);

AND2_X4 c2136(
.A1(net2182),
.A2(net2216),
.ZN(net2220)
);

AND2_X1 c2137(
.A1(net2190),
.A2(net2220),
.ZN(net2221)
);

NOR3_X2 c2138(
.A1(net2170),
.A2(net2211),
.A3(net2147),
.ZN(net2222)
);

AND3_X4 c2139(
.A1(net2218),
.A2(net2208),
.A3(net2197),
.ZN(net2223)
);

SDFF_X2 c2140(
.D(net2214),
.SE(net2220),
.SI(net1189),
.CK(clk),
.Q(net2225),
.QN(net2224)
);

NAND3_X2 c2141(
.A1(net2198),
.A2(net2188),
.A3(net2113),
.ZN(net2226)
);

NAND2_X1 c2142(
.A1(net2191),
.A2(net2218),
.ZN(net2227)
);

NAND2_X2 c2143(
.A1(net1237),
.A2(net2125),
.ZN(net2228)
);

NAND2_X4 c2144(
.A1(net2210),
.A2(net2227),
.ZN(net2229)
);

OR3_X1 c2145(
.A1(net283),
.A2(net2217),
.A3(net2209),
.ZN(net2230)
);

MUX2_X1 c2146(
.A(net2174),
.B(net2219),
.S(net2225),
.Z(net2231)
);

OAI21_X4 c2147(
.A(net2217),
.B1(net1934),
.B2(net11023),
.ZN(net2232)
);

AND2_X2 c2148(
.A1(net2221),
.A2(net2072),
.ZN(net2233)
);

XOR2_X1 c2149(
.A(net2176),
.B(net10845),
.Z(net2234)
);

MUX2_X2 c2150(
.A(net2217),
.B(net2205),
.S(net2156),
.Z(net2235)
);

NOR2_X1 c2151(
.A1(net2219),
.A2(net2178),
.ZN(net2236)
);

OR2_X2 c2152(
.A1(net2199),
.A2(net2075),
.ZN(net2237)
);

NOR2_X4 c2153(
.A1(net2236),
.A2(net2200),
.ZN(net2238)
);

DFFRS_X1 c2154(
.D(net2237),
.RN(net2234),
.SN(net2238),
.CK(clk),
.Q(net2240),
.QN(net2239)
);

NOR2_X2 c2155(
.A1(net1245),
.A2(net2186),
.ZN(net2241)
);

XOR2_X2 c2156(
.A(net1169),
.B(net2156),
.Z(net2242)
);

XNOR2_X1 c2157(
.A(net2241),
.B(net2177),
.ZN(net2243)
);

INV_X32 c2158(
.A(net2058),
.ZN(net2244)
);

INV_X4 c2159(
.A(net193),
.ZN(net2245)
);

OR2_X4 c2160(
.A1(net1339),
.A2(net327),
.ZN(net2246)
);

INV_X1 c2161(
.A(net33),
.ZN(net2247)
);

INV_X2 c2162(
.A(net2116),
.ZN(net2248)
);

INV_X8 c2163(
.A(net9591),
.ZN(net2249)
);

OR2_X1 c2164(
.A1(net1210),
.A2(net2204),
.ZN(net2250)
);

NAND3_X4 c2165(
.A1(net1262),
.A2(net2107),
.A3(net2247),
.ZN(net2251)
);

INV_X16 c2166(
.A(net2246),
.ZN(net2252)
);

XNOR2_X2 c2167(
.A(net2249),
.B(net1322),
.ZN(net2253)
);

CLKGATETST_X1 c2168(
.E(net1356),
.SE(net2228),
.CK(clk),
.GCK(net2254)
);

AND2_X4 c2169(
.A1(net2245),
.A2(net10874),
.ZN(net2255)
);

AND2_X1 c2170(
.A1(net2243),
.A2(net283),
.ZN(net2256)
);

NAND2_X1 c2171(
.A1(net2216),
.A2(net370),
.ZN(net2257)
);

INV_X32 c2172(
.A(net10824),
.ZN(net2258)
);

NAND2_X2 c2173(
.A1(net2258),
.A2(net1297),
.ZN(net2259)
);

NAND2_X4 c2174(
.A1(net2248),
.A2(net1186),
.ZN(net2260)
);

AND2_X2 c2175(
.A1(net1331),
.A2(net1355),
.ZN(net2261)
);

INV_X4 c2176(
.A(net311),
.ZN(net2262)
);

XOR2_X1 c2177(
.A(net310),
.B(net10727),
.Z(net2263)
);

INV_X1 c2178(
.A(net9591),
.ZN(net2264)
);

NOR2_X1 c2179(
.A1(net2264),
.A2(net2263),
.ZN(net2265)
);

INV_X2 c2180(
.A(net1340),
.ZN(net2266)
);

OR2_X2 c2181(
.A1(net344),
.A2(net2244),
.ZN(net2267)
);

INV_X8 c2182(
.A(net10254),
.ZN(net2268)
);

OR3_X4 c2183(
.A1(net1197),
.A2(net1332),
.A3(net1174),
.ZN(net2269)
);

NOR2_X4 c2184(
.A1(net2155),
.A2(net1299),
.ZN(net2270)
);

NOR2_X2 c2185(
.A1(net2250),
.A2(net1331),
.ZN(net2271)
);

XOR2_X2 c2186(
.A(net2107),
.B(net2267),
.Z(net2272)
);

XNOR2_X1 c2187(
.A(net1289),
.B(net1299),
.ZN(net2273)
);

OR2_X4 c2188(
.A1(net2252),
.A2(net2271),
.ZN(net2274)
);

INV_X16 c2189(
.A(net9940),
.ZN(net2275)
);

INV_X32 c2190(
.A(net1236),
.ZN(net2276)
);

OR2_X1 c2191(
.A1(net1084),
.A2(net2268),
.ZN(net2277)
);

XNOR2_X2 c2192(
.A(net1299),
.B(net327),
.ZN(net2278)
);

INV_X4 c2193(
.A(net377),
.ZN(net2279)
);

AND2_X4 c2194(
.A1(net2274),
.A2(net1324),
.ZN(net2280)
);

INV_X1 c2195(
.A(net2256),
.ZN(net2281)
);

AND2_X1 c2196(
.A1(net2270),
.A2(net2248),
.ZN(net2282)
);

NAND2_X1 c2197(
.A1(net1350),
.A2(net2250),
.ZN(net2283)
);

NAND2_X2 c2198(
.A1(net2253),
.A2(net2204),
.ZN(net2284)
);

NAND2_X4 c2199(
.A1(net2265),
.A2(net2227),
.ZN(net2285)
);

AND2_X2 c2200(
.A1(net2282),
.A2(net2250),
.ZN(net2286)
);

XOR2_X1 c2201(
.A(net10727),
.B(net10854),
.Z(net2287)
);

AND3_X2 c2202(
.A1(net2270),
.A2(net2283),
.A3(net10821),
.ZN(net2288)
);

NOR2_X1 c2203(
.A1(net402),
.A2(net2287),
.ZN(net2289)
);

INV_X2 c2204(
.A(net10058),
.ZN(net2290)
);

NOR3_X1 c2205(
.A1(net2260),
.A2(net2281),
.A3(net2271),
.ZN(net2291)
);

OR2_X2 c2206(
.A1(net1314),
.A2(net2254),
.ZN(net2292)
);

SDFFRS_X1 c2207(
.D(net2172),
.RN(net2215),
.SE(net1292),
.SI(net2224),
.SN(net1360),
.CK(clk),
.Q(net2294),
.QN(net2293)
);

NOR2_X4 c2208(
.A1(net2262),
.A2(net2290),
.ZN(net2295)
);

AOI222_X4 c2209(
.A1(net1174),
.A2(net1342),
.B1(net2259),
.B2(net2268),
.C1(net2244),
.C2(net2248),
.ZN(net2296)
);

NOR2_X2 c2210(
.A1(net2288),
.A2(net10854),
.ZN(net2297)
);

XOR2_X2 c2211(
.A(net2018),
.B(net2271),
.Z(net2298)
);

XNOR2_X1 c2212(
.A(net1335),
.B(net2273),
.ZN(net2299)
);

OR2_X4 c2213(
.A1(net2181),
.A2(net2284),
.ZN(net2300)
);

OR2_X1 c2214(
.A1(net2292),
.A2(net2287),
.ZN(net2301)
);

SDFFRS_X2 c2215(
.D(net2298),
.RN(net2275),
.SE(net1329),
.SI(net401),
.SN(net11152),
.CK(clk),
.Q(net2303),
.QN(net2302)
);

OR3_X2 c2216(
.A1(net2276),
.A2(net1207),
.A3(net11121),
.ZN(net2304)
);

XNOR2_X2 c2217(
.A(net2270),
.B(net11028),
.ZN(net2305)
);

AND2_X4 c2218(
.A1(net327),
.A2(net1319),
.ZN(net2306)
);

AND2_X1 c2219(
.A1(net2289),
.A2(net2305),
.ZN(net2307)
);

OAI21_X2 c2220(
.A(net2268),
.B1(net2270),
.B2(net2244),
.ZN(net2308)
);

DFFRS_X2 c2221(
.D(net2272),
.RN(net2268),
.SN(net10816),
.CK(clk),
.Q(net2310),
.QN(net2309)
);

NAND2_X1 c2222(
.A1(net1207),
.A2(net2208),
.ZN(net2311)
);

NAND2_X2 c2223(
.A1(net370),
.A2(net2292),
.ZN(net2312)
);

NAND2_X4 c2224(
.A1(net1308),
.A2(net1230),
.ZN(net2313)
);

AND2_X2 c2225(
.A1(net2287),
.A2(net2254),
.ZN(net2314)
);

CLKGATETST_X2 c2226(
.E(net2272),
.SE(net2292),
.CK(clk),
.GCK(net2315)
);

XOR2_X1 c2227(
.A(net2311),
.B(net2309),
.Z(net2316)
);

OAI21_X1 c2228(
.A(net2247),
.B1(net276),
.B2(net2301),
.ZN(net2317)
);

OAI33_X1 c2229(
.A1(net2310),
.A2(net1252),
.A3(net2287),
.B1(net1230),
.B2(net2248),
.B3(net1210),
.ZN(net2318)
);

AOI21_X2 c2230(
.A(net2259),
.B1(net1210),
.B2(net1356),
.ZN(net2319)
);

NOR2_X1 c2231(
.A1(net2319),
.A2(net2301),
.ZN(net2320)
);

AOI222_X2 c2232(
.A1(net2319),
.A2(net2302),
.B1(net2254),
.B2(net1070),
.C1(net2317),
.C2(net10806),
.ZN(net2321)
);

SDFF_X1 c2233(
.D(net2167),
.SE(net2288),
.SI(net2267),
.CK(clk),
.Q(net2323),
.QN(net2322)
);

SDFF_X2 c2234(
.D(net2126),
.SE(net2323),
.SI(net2320),
.CK(clk),
.Q(net2325),
.QN(net2324)
);

AOI21_X1 c2235(
.A(net2316),
.B1(net2325),
.B2(net2116),
.ZN(net2326)
);

AOI21_X4 c2236(
.A(net1329),
.B1(net2303),
.B2(net11038),
.ZN(net2327)
);

DFFRS_X1 c2237(
.D(net2318),
.RN(net2320),
.SN(net2058),
.CK(clk),
.Q(net2329),
.QN(net2328)
);

OAI222_X1 c2238(
.A1(net2326),
.A2(net2301),
.B1(net1350),
.B2(net2320),
.C1(net2302),
.C2(net2224),
.ZN(net2330)
);

AOI211_X1 c2239(
.A(net2135),
.B(net2295),
.C1(net2301),
.C2(net1292),
.ZN(net2331)
);

AND3_X1 c2240(
.A1(net1084),
.A2(net2320),
.A3(net10992),
.ZN(net2332)
);

INV_X8 c2241(
.A(net2267),
.ZN(net2333)
);

INV_X16 c2242(
.A(net11013),
.ZN(net2334)
);

INV_X32 c2243(
.A(net10803),
.ZN(net2335)
);

INV_X4 c2244(
.A(net2327),
.ZN(net2336)
);

OR2_X2 c2245(
.A1(net2277),
.A2(net2336),
.ZN(net2337)
);

NAND3_X1 c2246(
.A1(net2228),
.A2(net2277),
.A3(net2322),
.ZN(net2338)
);

INV_X1 c2247(
.A(net2301),
.ZN(net2339)
);

NOR3_X4 c2248(
.A1(net1403),
.A2(net1360),
.A3(net350),
.ZN(net2340)
);

OAI221_X1 c2249(
.A(net2306),
.B1(net2339),
.B2(net2225),
.C1(net1382),
.C2(net1408),
.ZN(net2341)
);

NOR2_X4 c2250(
.A1(net2315),
.A2(net425),
.ZN(net2342)
);

INV_X2 c2251(
.A(net10986),
.ZN(net2343)
);

NOR3_X2 c2252(
.A1(net2227),
.A2(net1408),
.A3(net1446),
.ZN(net2344)
);

NOR2_X2 c2253(
.A1(net1384),
.A2(net10816),
.ZN(net2345)
);

INV_X8 c2254(
.A(net1136),
.ZN(net2346)
);

INV_X16 c2255(
.A(net2323),
.ZN(net2347)
);

INV_X32 c2256(
.A(net2347),
.ZN(net2348)
);

XOR2_X2 c2257(
.A(net457),
.B(net1444),
.Z(net2349)
);

AND3_X4 c2258(
.A1(net1440),
.A2(net442),
.A3(net1355),
.ZN(net2350)
);

INV_X4 c2259(
.A(net9629),
.ZN(net2351)
);

INV_X1 c2260(
.A(net2341),
.ZN(net2352)
);

INV_X2 c2261(
.A(net9629),
.ZN(net2353)
);

INV_X8 c2262(
.A(net2283),
.ZN(net2354)
);

XNOR2_X1 c2263(
.A(net2204),
.B(net2346),
.ZN(net2355)
);

OR2_X4 c2264(
.A1(net2335),
.A2(net2339),
.ZN(net2356)
);

OR2_X1 c2265(
.A1(net2220),
.A2(net418),
.ZN(net2357)
);

XNOR2_X2 c2266(
.A(net2340),
.B(net2349),
.ZN(net2358)
);

CLKGATETST_X4 c2267(
.E(net2352),
.SE(net2228),
.CK(clk),
.GCK(net2359)
);

AND2_X4 c2268(
.A1(net2357),
.A2(net2248),
.ZN(net2360)
);

INV_X16 c2269(
.A(net1447),
.ZN(net2361)
);

NAND3_X2 c2270(
.A1(net442),
.A2(net1423),
.A3(net2312),
.ZN(net2362)
);

AND2_X1 c2271(
.A1(net2343),
.A2(net2348),
.ZN(net2363)
);

NAND2_X1 c2272(
.A1(net1424),
.A2(net2225),
.ZN(net2364)
);

NAND2_X2 c2273(
.A1(net2363),
.A2(net2255),
.ZN(net2365)
);

NAND2_X4 c2274(
.A1(net1360),
.A2(net10502),
.ZN(net2366)
);

AND2_X2 c2275(
.A1(net2353),
.A2(net2356),
.ZN(net2367)
);

XOR2_X1 c2276(
.A(net2367),
.B(net2356),
.Z(net2368)
);

NOR2_X1 c2277(
.A1(net2365),
.A2(net2308),
.ZN(net2369)
);

OR2_X2 c2278(
.A1(net2255),
.A2(net1210),
.ZN(net2370)
);

NOR2_X4 c2279(
.A1(net1360),
.A2(net1414),
.ZN(net2371)
);

NOR2_X2 c2280(
.A1(net1324),
.A2(net2365),
.ZN(net2372)
);

DFFRS_X2 c2281(
.D(net2369),
.RN(net2342),
.SN(net1208),
.CK(clk),
.Q(net2374),
.QN(net2373)
);

INV_X32 c2282(
.A(net425),
.ZN(net2375)
);

INV_X4 c2283(
.A(net11078),
.ZN(net2376)
);

XOR2_X2 c2284(
.A(net2359),
.B(net2349),
.Z(net2377)
);

XNOR2_X1 c2285(
.A(net2125),
.B(net2319),
.ZN(net2378)
);

OR2_X4 c2286(
.A1(net2371),
.A2(net1444),
.ZN(net2379)
);

OR3_X1 c2287(
.A1(net1426),
.A2(net2359),
.A3(net2376),
.ZN(net2380)
);

OR2_X1 c2288(
.A1(net2342),
.A2(net2380),
.ZN(net2381)
);

XNOR2_X2 c2289(
.A(net2381),
.B(net2356),
.ZN(net2382)
);

AND2_X4 c2290(
.A1(net1375),
.A2(net1324),
.ZN(net2383)
);

OAI221_X4 c2291(
.A(net2368),
.B1(net442),
.B2(net2209),
.C1(net2356),
.C2(net11013),
.ZN(net2384)
);

AND2_X1 c2292(
.A1(net2336),
.A2(net2303),
.ZN(net2385)
);

NAND2_X1 c2293(
.A1(net2375),
.A2(net10502),
.ZN(net2386)
);

NAND2_X2 c2294(
.A1(net2361),
.A2(net1279),
.ZN(net2387)
);

CLKGATETST_X8 c2295(
.E(net2378),
.SE(net2333),
.CK(clk),
.GCK(net2388)
);

INV_X1 c2296(
.A(net2387),
.ZN(net2389)
);

NAND2_X4 c2297(
.A1(net1070),
.A2(net2358),
.ZN(net2390)
);

INV_X2 c2298(
.A(net11132),
.ZN(net2391)
);

INV_X8 c2299(
.A(net10857),
.ZN(net2392)
);

AND2_X2 c2300(
.A1(net2390),
.A2(net2376),
.ZN(net2393)
);

XOR2_X1 c2301(
.A(net2358),
.B(net425),
.Z(net2394)
);

SDFF_X1 c2302(
.D(net1410),
.SE(net421),
.SI(net2315),
.CK(clk),
.Q(net2396),
.QN(net2395)
);

INV_X16 c2303(
.A(net2388),
.ZN(net2397)
);

MUX2_X1 c2304(
.A(net2394),
.B(net2388),
.S(net2368),
.Z(net2398)
);

NOR2_X1 c2305(
.A1(net2372),
.A2(net2340),
.ZN(net2399)
);

OR2_X2 c2306(
.A1(net1391),
.A2(net2391),
.ZN(net2400)
);

NOR2_X4 c2307(
.A1(net2383),
.A2(net2377),
.ZN(net2401)
);

NOR2_X2 c2308(
.A1(net2339),
.A2(net2358),
.ZN(net2402)
);

SDFF_X2 c2309(
.D(net2344),
.SE(net2401),
.SI(net2402),
.CK(clk),
.Q(net2404),
.QN(net2403)
);

INV_X32 c2310(
.A(net10355),
.ZN(net2405)
);

XOR2_X2 c2311(
.A(net2351),
.B(net2396),
.Z(net2406)
);

NAND4_X2 c2312(
.A1(net2396),
.A2(net1411),
.A3(net2403),
.A4(net2402),
.ZN(net2407)
);

OAI222_X4 c2313(
.A1(net2225),
.A2(net2373),
.B1(net2406),
.B2(net2317),
.C1(net2401),
.C2(net2333),
.ZN(net2408)
);

XNOR2_X1 c2314(
.A(net1411),
.B(net2389),
.ZN(net2409)
);

SDFFR_X2 c2315(
.D(net2407),
.RN(net2319),
.SE(net2401),
.SI(net10670),
.CK(clk),
.Q(net2411),
.QN(net2410)
);

OAI21_X4 c2316(
.A(net2393),
.B1(net2399),
.B2(net2403),
.ZN(net2412)
);

OAI222_X2 c2317(
.A1(net2392),
.A2(net2404),
.B1(net2412),
.B2(net2395),
.C1(net2401),
.C2(net1070),
.ZN(net2413)
);

OAI221_X2 c2318(
.A(net2401),
.B1(net2396),
.B2(net2400),
.C1(net2356),
.C2(net2402),
.ZN(net2414)
);

MUX2_X2 c2319(
.A(net1423),
.B(net2401),
.S(net1291),
.Z(net2415)
);

OR4_X4 c2320(
.A1(net2412),
.A2(net2391),
.A3(net2401),
.A4(net11164),
.ZN(net2416)
);

AOI221_X4 c2321(
.A(net2308),
.B1(net2407),
.B2(net2412),
.C1(net2401),
.C2(net2203),
.ZN(net2417)
);

AOI222_X1 c2322(
.A1(net2315),
.A2(net2402),
.B1(net2412),
.B2(net2395),
.C1(net2410),
.C2(net10657),
.ZN(net2418)
);

DFFRS_X1 c2323(
.D(net2405),
.RN(net2412),
.SN(net10552),
.CK(clk),
.Q(net2420),
.QN(net2419)
);

INV_X4 c2324(
.A(net1488),
.ZN(net2421)
);

INV_X1 c2325(
.A(net11075),
.ZN(net2422)
);

OR2_X4 c2326(
.A1(net2415),
.A2(net2386),
.ZN(net2423)
);

INV_X2 c2327(
.A(net527),
.ZN(net2424)
);

INV_X8 c2328(
.A(net2422),
.ZN(net2425)
);

AOI222_X4 c2329(
.A1(net2334),
.A2(net1380),
.B1(net1506),
.B2(net1408),
.C1(net1493),
.C2(net10826),
.ZN(net2426)
);

NAND3_X4 c2330(
.A1(net2319),
.A2(net2329),
.A3(net1355),
.ZN(net2427)
);

INV_X16 c2331(
.A(net11048),
.ZN(net2428)
);

INV_X32 c2332(
.A(net10442),
.ZN(net2429)
);

INV_X4 c2333(
.A(net2406),
.ZN(net2430)
);

OR2_X1 c2334(
.A1(net1510),
.A2(net11002),
.ZN(net2431)
);

XNOR2_X2 c2335(
.A(net2429),
.B(net2415),
.ZN(net2432)
);

INV_X1 c2336(
.A(net10442),
.ZN(net2433)
);

AND2_X4 c2337(
.A1(net1480),
.A2(net2426),
.ZN(net2434)
);

AND2_X1 c2338(
.A1(net2431),
.A2(net489),
.ZN(net2435)
);

NAND2_X1 c2339(
.A1(net1195),
.A2(net1459),
.ZN(net2436)
);

INV_X2 c2340(
.A(net2366),
.ZN(net2437)
);

INV_X8 c2341(
.A(net2433),
.ZN(net2438)
);

NAND2_X2 c2342(
.A1(net2437),
.A2(net2110),
.ZN(net2439)
);

NAND2_X4 c2343(
.A1(net2312),
.A2(net11162),
.ZN(net2440)
);

INV_X16 c2344(
.A(net2439),
.ZN(net2441)
);

AND2_X2 c2345(
.A1(net2391),
.A2(net2435),
.ZN(net2442)
);

INV_X32 c2346(
.A(net10343),
.ZN(net2443)
);

XOR2_X1 c2347(
.A(net2386),
.B(net2380),
.Z(net2444)
);

DFFR_X1 c2348(
.D(net2423),
.RN(net1505),
.CK(clk),
.Q(net2446),
.QN(net2445)
);

NOR2_X1 c2349(
.A1(net2428),
.A2(net2445),
.ZN(net2447)
);

DFFR_X2 c2350(
.D(net1537),
.RN(net2434),
.CK(clk),
.Q(net2449),
.QN(net2448)
);

OR2_X2 c2351(
.A1(net2424),
.A2(net2428),
.ZN(net2450)
);

NOR2_X4 c2352(
.A1(net2450),
.A2(net2440),
.ZN(net2451)
);

OR3_X4 c2353(
.A1(net2446),
.A2(net2279),
.A3(net1506),
.ZN(net2452)
);

INV_X4 c2354(
.A(net1499),
.ZN(net2453)
);

NOR2_X2 c2355(
.A1(net2430),
.A2(net2450),
.ZN(net2454)
);

INV_X1 c2356(
.A(net2440),
.ZN(net2455)
);

INV_X2 c2357(
.A(net1512),
.ZN(net2456)
);

DFFRS_X2 c2358(
.D(net1532),
.RN(net2439),
.SN(net1398),
.CK(clk),
.Q(net2458),
.QN(net2457)
);

AOI221_X2 c2359(
.A(net2325),
.B1(net2430),
.B2(net2451),
.C1(net2440),
.C2(net1493),
.ZN(net2459)
);

INV_X8 c2360(
.A(net10916),
.ZN(net2460)
);

XOR2_X2 c2361(
.A(net2426),
.B(net2443),
.Z(net2461)
);

DFFS_X1 c2362(
.D(net2443),
.SN(net2337),
.CK(clk),
.Q(net2463),
.QN(net2462)
);

XNOR2_X1 c2363(
.A(net2380),
.B(net2415),
.ZN(net2464)
);

OR2_X4 c2364(
.A1(net2436),
.A2(net2457),
.ZN(net2465)
);

INV_X16 c2365(
.A(net10442),
.ZN(net2466)
);

OR2_X1 c2366(
.A1(net2290),
.A2(net2421),
.ZN(net2467)
);

INV_X32 c2367(
.A(net2379),
.ZN(net2468)
);

XNOR2_X2 c2368(
.A(net2328),
.B(net11038),
.ZN(net2469)
);

AND2_X4 c2369(
.A1(net2447),
.A2(net11155),
.ZN(net2470)
);

AND3_X2 c2370(
.A1(net1448),
.A2(net2446),
.A3(net2334),
.ZN(net2471)
);

AND2_X1 c2371(
.A1(net2443),
.A2(net339),
.ZN(net2472)
);

NAND2_X1 c2372(
.A1(net2459),
.A2(net2380),
.ZN(net2473)
);

INV_X4 c2373(
.A(net2463),
.ZN(net2474)
);

NAND2_X2 c2374(
.A1(net1469),
.A2(net2464),
.ZN(net2475)
);

NAND2_X4 c2375(
.A1(net2370),
.A2(net2449),
.ZN(net2476)
);

INV_X1 c2376(
.A(net1521),
.ZN(net2477)
);

AND2_X2 c2377(
.A1(net516),
.A2(net11154),
.ZN(net2478)
);

XOR2_X1 c2378(
.A(net1450),
.B(net2345),
.Z(net2479)
);

INV_X2 c2379(
.A(net2471),
.ZN(net2480)
);

NOR2_X1 c2380(
.A1(net1528),
.A2(net2440),
.ZN(net2481)
);

INV_X8 c2381(
.A(net10003),
.ZN(net2482)
);

OR2_X2 c2382(
.A1(net2466),
.A2(net2463),
.ZN(net2483)
);

OAI33_X1 c2383(
.A1(net2456),
.A2(net2452),
.A3(net2370),
.B1(net2443),
.B2(net1380),
.B3(net2447),
.ZN(net2484)
);

NOR3_X1 c2384(
.A1(net514),
.A2(net2441),
.A3(net1493),
.ZN(net2485)
);

NOR2_X4 c2385(
.A1(net2479),
.A2(net2478),
.ZN(net2486)
);

INV_X16 c2386(
.A(net10810),
.ZN(net2487)
);

OR3_X2 c2387(
.A1(net2468),
.A2(net2437),
.A3(net2454),
.ZN(net2488)
);

NOR2_X2 c2388(
.A1(net2482),
.A2(net2447),
.ZN(net2489)
);

XOR2_X2 c2389(
.A(net2489),
.B(net2445),
.Z(net2490)
);

SDFF_X1 c2390(
.D(net2488),
.SE(net2465),
.SI(net1521),
.CK(clk),
.Q(net2492),
.QN(net2491)
);

OAI21_X2 c2391(
.A(net2428),
.B1(net2443),
.B2(net2490),
.ZN(net2493)
);

XNOR2_X1 c2392(
.A(net2439),
.B(net2490),
.ZN(net2494)
);

OR2_X4 c2393(
.A1(net2480),
.A2(net2487),
.ZN(net2495)
);

OR2_X1 c2394(
.A1(net2451),
.A2(net459),
.ZN(net2496)
);

XNOR2_X2 c2395(
.A(net2452),
.B(net2494),
.ZN(net2497)
);

SDFFRS_X1 c2396(
.D(net2444),
.RN(net2492),
.SE(net2493),
.SI(net1521),
.SN(net2425),
.CK(clk),
.Q(net2499),
.QN(net2498)
);

AND2_X4 c2397(
.A1(net2442),
.A2(net2497),
.ZN(net2500)
);

AOI222_X2 c2398(
.A1(net2476),
.A2(net2462),
.B1(net2490),
.B2(net1493),
.C1(net1355),
.C2(net11165),
.ZN(net2501)
);

INV_X32 c2399(
.A(net11048),
.ZN(net2502)
);

AND2_X1 c2400(
.A1(net2502),
.A2(net2443),
.ZN(net2503)
);

OAI21_X1 c2401(
.A(net2495),
.B1(net2271),
.B2(net2425),
.ZN(net2504)
);

AOI21_X2 c2402(
.A(net2503),
.B1(net2458),
.B2(net2464),
.ZN(net2505)
);

INV_X4 c2403(
.A(net10782),
.ZN(net2506)
);

INV_X1 c2404(
.A(net10243),
.ZN(net2507)
);

SDFF_X2 c2405(
.D(net2507),
.SE(net2486),
.SI(net2504),
.CK(clk),
.Q(net2509),
.QN(net2508)
);

AOI221_X1 c2406(
.A(net2464),
.B1(net2485),
.B2(net1493),
.C1(net2508),
.C2(net2491),
.ZN(net2510)
);

INV_X2 c2407(
.A(net9947),
.ZN(net2511)
);

INV_X8 c2408(
.A(net1624),
.ZN(net2512)
);

NAND2_X1 c2409(
.A1(net1484),
.A2(net2494),
.ZN(net2513)
);

INV_X16 c2410(
.A(net9604),
.ZN(net2514)
);

INV_X32 c2411(
.A(net1427),
.ZN(net2515)
);

INV_X4 c2412(
.A(net2513),
.ZN(net2516)
);

INV_X1 c2413(
.A(net9734),
.ZN(net2517)
);

AOI21_X1 c2414(
.A(net2110),
.B1(net2517),
.B2(net1493),
.ZN(net2518)
);

INV_X2 c2415(
.A(net10100),
.ZN(net2519)
);

INV_X8 c2416(
.A(net1611),
.ZN(net2520)
);

AOI21_X4 c2417(
.A(net2511),
.B1(net2519),
.B2(net10670),
.ZN(net2521)
);

INV_X16 c2418(
.A(net588),
.ZN(net2522)
);

INV_X32 c2419(
.A(net1560),
.ZN(net2523)
);

NAND2_X2 c2420(
.A1(net2521),
.A2(net1599),
.ZN(net2524)
);

NAND2_X4 c2421(
.A1(net1564),
.A2(net2518),
.ZN(net2525)
);

AND2_X2 c2422(
.A1(net2467),
.A2(net11163),
.ZN(net2526)
);

XOR2_X1 c2423(
.A(net2271),
.B(net2521),
.Z(net2527)
);

INV_X4 c2424(
.A(net9728),
.ZN(net2528)
);

INV_X1 c2425(
.A(net2522),
.ZN(net2529)
);

OAI22_X2 c2426(
.A1(net2512),
.A2(net1587),
.B1(net1612),
.B2(net2425),
.ZN(net2530)
);

NOR2_X1 c2427(
.A1(net2529),
.A2(net2519),
.ZN(net2531)
);

OR2_X2 c2428(
.A1(net2523),
.A2(net1626),
.ZN(net2532)
);

NOR2_X4 c2429(
.A1(net2493),
.A2(net2474),
.ZN(net2533)
);

NOR2_X2 c2430(
.A1(net597),
.A2(net2435),
.ZN(net2534)
);

INV_X2 c2431(
.A(net647),
.ZN(net2535)
);

INV_X8 c2432(
.A(net10144),
.ZN(net2536)
);

AND3_X1 c2433(
.A1(net2447),
.A2(net2527),
.A3(net2421),
.ZN(net2537)
);

INV_X16 c2434(
.A(net11085),
.ZN(net2538)
);

XOR2_X2 c2435(
.A(net2435),
.B(net2534),
.Z(net2539)
);

DFFRS_X1 c2436(
.D(net2527),
.RN(net2530),
.SN(net2531),
.CK(clk),
.Q(net2541),
.QN(net2540)
);

XNOR2_X1 c2437(
.A(net608),
.B(net2517),
.ZN(net2542)
);

OR2_X4 c2438(
.A1(net2536),
.A2(net1574),
.ZN(net2543)
);

INV_X32 c2439(
.A(net10150),
.ZN(net2544)
);

OR2_X1 c2440(
.A1(net2526),
.A2(net2541),
.ZN(net2545)
);

XNOR2_X2 c2441(
.A(net2542),
.B(net2421),
.ZN(net2546)
);

NAND3_X1 c2442(
.A1(net2543),
.A2(net2529),
.A3(net2545),
.ZN(net2547)
);

AND2_X4 c2443(
.A1(net2438),
.A2(net10392),
.ZN(net2548)
);

AND2_X1 c2444(
.A1(net2538),
.A2(net2271),
.ZN(net2549)
);

INV_X4 c2445(
.A(net9604),
.ZN(net2550)
);

INV_X1 c2446(
.A(net10366),
.ZN(net2551)
);

NOR3_X4 c2447(
.A1(net2517),
.A2(net2511),
.A3(net1584),
.ZN(net2552)
);

INV_X2 c2448(
.A(net10299),
.ZN(net2553)
);

OAI211_X4 c2449(
.A(net1408),
.B(net2551),
.C1(net2545),
.C2(net2346),
.ZN(net2554)
);

NAND2_X1 c2450(
.A1(net2467),
.A2(net1587),
.ZN(net2555)
);

NOR3_X2 c2451(
.A1(net2453),
.A2(net2475),
.A3(net10859),
.ZN(net2556)
);

DFFS_X2 c2452(
.D(net2465),
.SN(net10782),
.CK(clk),
.Q(net2558),
.QN(net2557)
);

NAND2_X2 c2453(
.A1(net2535),
.A2(net459),
.ZN(net2559)
);

NAND2_X4 c2454(
.A1(net2541),
.A2(net2493),
.ZN(net2560)
);

AND2_X2 c2455(
.A1(net2551),
.A2(net2472),
.ZN(net2561)
);

XOR2_X1 c2456(
.A(net2545),
.B(net1627),
.Z(net2562)
);

NOR2_X1 c2457(
.A1(net2560),
.A2(net2517),
.ZN(net2563)
);

INV_X8 c2458(
.A(net2432),
.ZN(net2564)
);

AND3_X4 c2459(
.A1(net2555),
.A2(net2544),
.A3(net2519),
.ZN(net2565)
);

NAND3_X2 c2460(
.A1(net2528),
.A2(net2545),
.A3(net1589),
.ZN(net2566)
);

OR2_X2 c2461(
.A1(net1613),
.A2(net1626),
.ZN(net2567)
);

NOR2_X4 c2462(
.A1(net2400),
.A2(net1624),
.ZN(net2568)
);

NOR2_X2 c2463(
.A1(net1612),
.A2(net1408),
.ZN(net2569)
);

INV_X16 c2464(
.A(net2568),
.ZN(net2570)
);

XOR2_X2 c2465(
.A(net1598),
.B(net10834),
.Z(net2571)
);

XNOR2_X1 c2466(
.A(net2563),
.B(net1615),
.ZN(net2572)
);

INV_X32 c2467(
.A(net2548),
.ZN(net2573)
);

OR2_X4 c2468(
.A1(net2511),
.A2(net2545),
.ZN(net2574)
);

INV_X4 c2469(
.A(net10392),
.ZN(net2575)
);

OR2_X1 c2470(
.A1(net2575),
.A2(net630),
.ZN(net2576)
);

XNOR2_X2 c2471(
.A(net2421),
.B(net1560),
.ZN(net2577)
);

AND2_X4 c2472(
.A1(net2576),
.A2(net2574),
.ZN(net2578)
);

AND2_X1 c2473(
.A1(net350),
.A2(net2346),
.ZN(net2579)
);

NAND2_X1 c2474(
.A1(net2474),
.A2(net2540),
.ZN(net2580)
);

NAND2_X2 c2475(
.A1(net2571),
.A2(net2568),
.ZN(net2581)
);

NAND2_X4 c2476(
.A1(net1598),
.A2(net2544),
.ZN(net2582)
);

AND2_X2 c2477(
.A1(net2580),
.A2(net2568),
.ZN(net2583)
);

SDFFS_X1 c2478(
.D(net643),
.SE(net2583),
.SI(net2493),
.SN(net1615),
.CK(clk),
.Q(net2585),
.QN(net2584)
);

OAI211_X1 c2479(
.A(net2577),
.B(net1623),
.C1(net1615),
.C2(net11165),
.ZN(net2586)
);

XOR2_X1 c2480(
.A(net2559),
.B(net2572),
.Z(net2587)
);

INV_X1 c2481(
.A(net9812),
.ZN(net2588)
);

OR3_X1 c2482(
.A1(net2519),
.A2(net2580),
.A3(net2535),
.ZN(net2589)
);

NOR4_X4 c2483(
.A1(net2586),
.A2(net2584),
.A3(net2589),
.A4(net2557),
.ZN(net2590)
);

NOR2_X1 c2484(
.A1(net2562),
.A2(net2572),
.ZN(net2591)
);

NOR4_X2 c2485(
.A1(net2588),
.A2(net2574),
.A3(net2467),
.A4(net647),
.ZN(net2592)
);

MUX2_X1 c2486(
.A(net2202),
.B(net2536),
.S(net2521),
.Z(net2593)
);

AOI211_X4 c2487(
.A(net2588),
.B(net2582),
.C1(net2593),
.C2(net10617),
.ZN(net2594)
);

OAI21_X4 c2488(
.A(net2579),
.B1(net2587),
.B2(net10834),
.ZN(net2595)
);

MUX2_X2 c2489(
.A(net2592),
.B(net2573),
.S(net10773),
.Z(net2596)
);

CLKGATETST_X1 c2490(
.E(net740),
.SE(net2510),
.CK(clk),
.GCK(net2597)
);

OR2_X2 c2491(
.A1(net1631),
.A2(net1622),
.ZN(net2598)
);

NOR2_X4 c2492(
.A1(net2524),
.A2(net2518),
.ZN(net2599)
);

INV_X2 c2493(
.A(net2426),
.ZN(net2600)
);

INV_X8 c2494(
.A(net1673),
.ZN(net2601)
);

NOR2_X2 c2495(
.A1(net2572),
.A2(net2520),
.ZN(net2602)
);

XOR2_X2 c2496(
.A(net2460),
.B(net2483),
.Z(net2603)
);

INV_X16 c2497(
.A(net9681),
.ZN(net2604)
);

NAND3_X4 c2498(
.A1(net2602),
.A2(net1579),
.A3(net695),
.ZN(net2605)
);

XNOR2_X1 c2499(
.A(net2603),
.B(net1673),
.ZN(net2606)
);

OR2_X4 c2500(
.A1(net1624),
.A2(net2606),
.ZN(net2607)
);

OR2_X1 c2501(
.A1(net2514),
.A2(net2600),
.ZN(net2608)
);

INV_X32 c2502(
.A(net11065),
.ZN(net2609)
);

XNOR2_X2 c2503(
.A(net2607),
.B(net2279),
.ZN(net2610)
);

INV_X4 c2504(
.A(net1354),
.ZN(net2611)
);

INV_X1 c2505(
.A(net1646),
.ZN(net2612)
);

AND2_X4 c2506(
.A1(net1622),
.A2(net695),
.ZN(net2613)
);

AND2_X1 c2507(
.A1(net2279),
.A2(net2572),
.ZN(net2614)
);

NAND2_X1 c2508(
.A1(net1682),
.A2(net1708),
.ZN(net2615)
);

OR3_X4 c2509(
.A1(net1503),
.A2(net1615),
.A3(net2441),
.ZN(net2616)
);

INV_X2 c2510(
.A(net10050),
.ZN(net2617)
);

NAND2_X2 c2511(
.A1(net2589),
.A2(net10860),
.ZN(net2618)
);

NAND2_X4 c2512(
.A1(net2532),
.A2(net2514),
.ZN(net2619)
);

AND2_X2 c2513(
.A1(net674),
.A2(net2589),
.ZN(net2620)
);

XOR2_X1 c2514(
.A(net1665),
.B(net2447),
.Z(net2621)
);

NOR2_X1 c2515(
.A1(net2438),
.A2(net2534),
.ZN(net2622)
);

INV_X8 c2516(
.A(net10883),
.ZN(net2623)
);

INV_X16 c2517(
.A(net11047),
.ZN(net2624)
);

OR2_X2 c2518(
.A1(net1675),
.A2(net2612),
.ZN(net2625)
);

NOR2_X4 c2519(
.A1(net1672),
.A2(net1696),
.ZN(net2626)
);

INV_X32 c2520(
.A(net10098),
.ZN(net2627)
);

AND3_X2 c2521(
.A1(net2520),
.A2(net2601),
.A3(net2610),
.ZN(net2628)
);

NOR2_X2 c2522(
.A1(net2617),
.A2(net1676),
.ZN(net2629)
);

XOR2_X2 c2523(
.A(net2619),
.B(net2532),
.Z(net2630)
);

INV_X4 c2524(
.A(net9681),
.ZN(net2631)
);

INV_X1 c2525(
.A(net9843),
.ZN(net2632)
);

INV_X2 c2526(
.A(net2469),
.ZN(net2633)
);

XNOR2_X1 c2527(
.A(net1709),
.B(net2629),
.ZN(net2634)
);

NOR4_X1 c2528(
.A1(net2611),
.A2(net1672),
.A3(net2632),
.A4(net2612),
.ZN(net2635)
);

INV_X8 c2529(
.A(net1669),
.ZN(net2636)
);

OR2_X4 c2530(
.A1(net2636),
.A2(net1711),
.ZN(net2637)
);

OR2_X1 c2531(
.A1(net2629),
.A2(net10439),
.ZN(net2638)
);

INV_X16 c2532(
.A(net10271),
.ZN(net2639)
);

XNOR2_X2 c2533(
.A(net2638),
.B(net2425),
.ZN(net2640)
);

OAI221_X1 c2534(
.A(net2441),
.B1(net2633),
.B2(net2623),
.C1(net1709),
.C2(net1380),
.ZN(net2641)
);

AND2_X4 c2535(
.A1(net1599),
.A2(net2518),
.ZN(net2642)
);

NOR3_X1 c2536(
.A1(net2599),
.A2(net2616),
.A3(net674),
.ZN(net2643)
);

AND2_X1 c2537(
.A1(net693),
.A2(net2603),
.ZN(net2644)
);

NAND2_X1 c2538(
.A1(net2640),
.A2(net2633),
.ZN(net2645)
);

NAND2_X2 c2539(
.A1(net2483),
.A2(net2633),
.ZN(net2646)
);

NAND2_X4 c2540(
.A1(net2627),
.A2(net2621),
.ZN(net2647)
);

CLKGATETST_X2 c2541(
.E(net2623),
.SE(net1683),
.CK(clk),
.GCK(net2648)
);

OR3_X2 c2542(
.A1(net2534),
.A2(net1669),
.A3(net2648),
.ZN(net2649)
);

CLKGATETST_X4 c2543(
.E(net2610),
.SE(net693),
.CK(clk),
.GCK(net2650)
);

AND2_X2 c2544(
.A1(net2374),
.A2(net2642),
.ZN(net2651)
);

XOR2_X1 c2545(
.A(net1640),
.B(net2648),
.Z(net2652)
);

INV_X32 c2546(
.A(net10870),
.ZN(net2653)
);

NOR2_X1 c2547(
.A1(net2518),
.A2(net2648),
.ZN(net2654)
);

OAI21_X2 c2548(
.A(net2654),
.B1(net2627),
.B2(net2642),
.ZN(net2655)
);

OR2_X2 c2549(
.A1(net1642),
.A2(net2607),
.ZN(net2656)
);

INV_X4 c2550(
.A(net10963),
.ZN(net2657)
);

NOR2_X4 c2551(
.A1(net2622),
.A2(net2649),
.ZN(net2658)
);

NOR2_X2 c2552(
.A1(net979),
.A2(net2648),
.ZN(net2659)
);

XOR2_X2 c2553(
.A(net1685),
.B(net2642),
.Z(net2660)
);

XNOR2_X1 c2554(
.A(net1690),
.B(net2634),
.ZN(net2661)
);

OR2_X4 c2555(
.A1(net2650),
.A2(net10882),
.ZN(net2662)
);

OR2_X1 c2556(
.A1(net2609),
.A2(net1681),
.ZN(net2663)
);

DFFRS_X2 c2557(
.D(net2635),
.RN(net2617),
.SN(net11039),
.CK(clk),
.Q(net2665),
.QN(net2664)
);

INV_X1 c2558(
.A(net10287),
.ZN(net2666)
);

XNOR2_X2 c2559(
.A(net2631),
.B(net2652),
.ZN(net2667)
);

OAI221_X4 c2560(
.A(net2666),
.B1(net2667),
.B2(net2447),
.C1(net687),
.C2(net2633),
.ZN(net2668)
);

INV_X2 c2561(
.A(net10097),
.ZN(net2669)
);

OAI21_X1 c2562(
.A(net2669),
.B1(net618),
.B2(net10930),
.ZN(net2670)
);

AND2_X4 c2563(
.A1(net2658),
.A2(net2657),
.ZN(net2671)
);

AOI21_X2 c2564(
.A(net2671),
.B1(net2670),
.B2(net2653),
.ZN(net2672)
);

OAI222_X1 c2565(
.A1(net2621),
.A2(net2667),
.B1(net746),
.B2(net1579),
.C1(net2658),
.C2(net2670),
.ZN(net2673)
);

AOI21_X1 c2566(
.A(net2539),
.B1(net2664),
.B2(net10930),
.ZN(net2674)
);

AOI21_X4 c2567(
.A(net2645),
.B1(net2673),
.B2(net11122),
.ZN(net2675)
);

AND2_X1 c2568(
.A1(net2648),
.A2(net2617),
.ZN(net2676)
);

AND3_X1 c2569(
.A1(net2669),
.A2(net2670),
.A3(net1707),
.ZN(net2677)
);

OAI221_X2 c2570(
.A(net2670),
.B1(net2653),
.B2(net2612),
.C1(net10654),
.C2(net11122),
.ZN(net2678)
);

NAND2_X1 c2571(
.A1(net2673),
.A2(net2646),
.ZN(net2679)
);

INV_X8 c2572(
.A(net10338),
.ZN(net2680)
);

INV_X16 c2573(
.A(net11025),
.ZN(net2681)
);

NAND2_X2 c2574(
.A1(net1777),
.A2(net2601),
.ZN(net2682)
);

INV_X32 c2575(
.A(net11109),
.ZN(net2683)
);

INV_X4 c2576(
.A(net800),
.ZN(net2684)
);

INV_X1 c2577(
.A(net2641),
.ZN(net2685)
);

INV_X2 c2578(
.A(net2615),
.ZN(net2686)
);

AOI211_X2 c2579(
.A(net1778),
.B(net1787),
.C1(net2544),
.C2(net2653),
.ZN(net2687)
);

NAND2_X4 c2580(
.A1(net1797),
.A2(net2634),
.ZN(net2688)
);

AND2_X2 c2581(
.A1(net2668),
.A2(net1777),
.ZN(net2689)
);

INV_X8 c2582(
.A(net1786),
.ZN(net2690)
);

NAND3_X1 c2583(
.A1(net2682),
.A2(net1681),
.A3(net1787),
.ZN(net2691)
);

INV_X16 c2584(
.A(net10330),
.ZN(net2692)
);

INV_X32 c2585(
.A(net9633),
.ZN(net2693)
);

INV_X4 c2586(
.A(net2604),
.ZN(net2694)
);

INV_X1 c2587(
.A(net10201),
.ZN(net2695)
);

XOR2_X1 c2588(
.A(net1479),
.B(net2498),
.Z(net2696)
);

NOR2_X1 c2589(
.A1(net2653),
.A2(net1729),
.ZN(net2697)
);

INV_X2 c2590(
.A(net2688),
.ZN(net2698)
);

INV_X8 c2591(
.A(net2652),
.ZN(net2699)
);

INV_X16 c2592(
.A(net2662),
.ZN(net2700)
);

NOR3_X4 c2593(
.A1(net2684),
.A2(net2686),
.A3(net2700),
.ZN(net2701)
);

INV_X32 c2594(
.A(net2601),
.ZN(net2702)
);

INV_X4 c2595(
.A(net11056),
.ZN(net2703)
);

OR2_X2 c2596(
.A1(net2543),
.A2(net1737),
.ZN(net2704)
);

NOR2_X4 c2597(
.A1(net2703),
.A2(net2653),
.ZN(net2705)
);

INV_X1 c2598(
.A(net11010),
.ZN(net2706)
);

INV_X2 c2599(
.A(net10439),
.ZN(net2707)
);

NOR2_X2 c2600(
.A1(net2697),
.A2(net1777),
.ZN(net2708)
);

NOR3_X2 c2601(
.A1(net2510),
.A2(net2650),
.A3(net2685),
.ZN(net2709)
);

XOR2_X2 c2602(
.A(net2692),
.B(net1575),
.Z(net2710)
);

XNOR2_X1 c2603(
.A(net1714),
.B(net798),
.ZN(net2711)
);

OR2_X4 c2604(
.A1(net822),
.A2(net2543),
.ZN(net2712)
);

OR2_X1 c2605(
.A1(net1780),
.A2(net2712),
.ZN(net2713)
);

INV_X8 c2606(
.A(net1769),
.ZN(net2714)
);

XNOR2_X2 c2607(
.A(net2707),
.B(net1753),
.ZN(net2715)
);

AND2_X4 c2608(
.A1(net1729),
.A2(net2670),
.ZN(net2716)
);

AND2_X1 c2609(
.A1(net2682),
.A2(net11033),
.ZN(net2717)
);

NAND2_X1 c2610(
.A1(net2676),
.A2(net1666),
.ZN(net2718)
);

INV_X16 c2611(
.A(net9633),
.ZN(net2719)
);

NAND2_X2 c2612(
.A1(net2718),
.A2(net687),
.ZN(net2720)
);

INV_X32 c2613(
.A(net10808),
.ZN(net2721)
);

NAND2_X4 c2614(
.A1(net2706),
.A2(net2544),
.ZN(net2722)
);

AND2_X2 c2615(
.A1(net2600),
.A2(net1714),
.ZN(net2723)
);

XOR2_X1 c2616(
.A(net2719),
.B(net11037),
.Z(net2724)
);

CLKGATETST_X8 c2617(
.E(net1795),
.SE(net2719),
.CK(clk),
.GCK(net2725)
);

NOR2_X1 c2618(
.A1(net2683),
.A2(net2719),
.ZN(net2726)
);

OR2_X2 c2619(
.A1(net2629),
.A2(net2726),
.ZN(net2727)
);

NOR2_X4 c2620(
.A1(net1792),
.A2(net618),
.ZN(net2728)
);

NOR2_X2 c2621(
.A1(net2698),
.A2(net2713),
.ZN(net2729)
);

XOR2_X2 c2622(
.A(net2713),
.B(net2634),
.Z(net2730)
);

AOI22_X1 c2623(
.A1(net2699),
.A2(net2712),
.B1(net2724),
.B2(net2714),
.ZN(net2731)
);

XNOR2_X1 c2624(
.A(net2730),
.B(net2729),
.ZN(net2732)
);

OR2_X4 c2625(
.A1(net2618),
.A2(net1786),
.ZN(net2733)
);

AOI221_X4 c2626(
.A(net2728),
.B1(net2689),
.B2(net1777),
.C1(net1720),
.C2(net2710),
.ZN(net2734)
);

AND3_X4 c2627(
.A1(net2689),
.A2(net2719),
.A3(net10913),
.ZN(net2735)
);

OR2_X1 c2628(
.A1(net2722),
.A2(net2729),
.ZN(net2736)
);

XNOR2_X2 c2629(
.A(net1771),
.B(net2653),
.ZN(net2737)
);

AND2_X4 c2630(
.A1(net2704),
.A2(net2702),
.ZN(net2738)
);

NAND3_X2 c2631(
.A1(net2735),
.A2(net2719),
.A3(net2684),
.ZN(net2739)
);

SDFF_X1 c2632(
.D(net2736),
.SE(net2732),
.SI(net2738),
.CK(clk),
.Q(net2741),
.QN(net2740)
);

AND2_X1 c2633(
.A1(net2701),
.A2(net2700),
.ZN(net2742)
);

NAND2_X1 c2634(
.A1(net2742),
.A2(net2740),
.ZN(net2743)
);

NAND2_X2 c2635(
.A1(net2702),
.A2(net2720),
.ZN(net2744)
);

INV_X4 c2636(
.A(net10808),
.ZN(net2745)
);

NAND2_X4 c2637(
.A1(net2717),
.A2(net11037),
.ZN(net2746)
);

SDFFS_X2 c2638(
.D(net2746),
.SE(net2725),
.SI(net2733),
.SN(net2719),
.CK(clk),
.Q(net2748),
.QN(net2747)
);

OR3_X1 c2639(
.A1(net2743),
.A2(net2472),
.A3(net2543),
.ZN(net2749)
);

AND2_X2 c2640(
.A1(net2329),
.A2(net2747),
.ZN(net2750)
);

AND4_X4 c2641(
.A1(net2659),
.A2(net2634),
.A3(net2747),
.A4(net2715),
.ZN(net2751)
);

XOR2_X1 c2642(
.A(net2717),
.B(net2751),
.Z(net2752)
);

AOI221_X2 c2643(
.A(net695),
.B1(net2558),
.B2(net2714),
.C1(net2710),
.C2(net11033),
.ZN(net2753)
);

NOR2_X1 c2644(
.A1(net2689),
.A2(net2746),
.ZN(net2754)
);

OR2_X2 c2645(
.A1(net2753),
.A2(net1647),
.ZN(net2755)
);

DFFR_X1 c2646(
.D(net2726),
.RN(net2754),
.CK(clk),
.Q(net2757),
.QN(net2756)
);

INV_X1 c2647(
.A(net11034),
.ZN(net2758)
);

NOR2_X4 c2648(
.A1(net2758),
.A2(net2748),
.ZN(net2759)
);

AOI221_X1 c2649(
.A(net2749),
.B1(net2746),
.B2(net2742),
.C1(net2759),
.C2(net2710),
.ZN(net2760)
);

NOR2_X2 c2650(
.A1(net2744),
.A2(net2713),
.ZN(net2761)
);

XOR2_X2 c2651(
.A(net2752),
.B(net2754),
.Z(net2762)
);

XNOR2_X1 c2652(
.A(net2734),
.B(net2756),
.ZN(net2763)
);

OR2_X4 c2653(
.A1(net2720),
.A2(net2757),
.ZN(net2764)
);

OR2_X1 c2654(
.A1(net1542),
.A2(net10729),
.ZN(net2765)
);

XNOR2_X2 c2655(
.A(net2756),
.B(net11037),
.ZN(net2766)
);

AND2_X4 c2656(
.A1(net1877),
.A2(net1836),
.ZN(net2767)
);

AND2_X1 c2657(
.A1(net1739),
.A2(net1814),
.ZN(net2768)
);

NAND2_X1 c2658(
.A1(net1807),
.A2(net2729),
.ZN(net2769)
);

MUX2_X1 c2659(
.A(net2695),
.B(net1863),
.S(net1727),
.Z(net2770)
);

OAI221_X1 c2660(
.A(net1696),
.B1(net927),
.B2(net851),
.C1(net2712),
.C2(net772),
.ZN(net2771)
);

DFFR_X2 c2661(
.D(net2587),
.RN(net10577),
.CK(clk),
.Q(net2773),
.QN(net2772)
);

NAND2_X2 c2662(
.A1(net922),
.A2(net2768),
.ZN(net2774)
);

INV_X2 c2663(
.A(net9644),
.ZN(net2775)
);

NAND2_X4 c2664(
.A1(net1847),
.A2(net2773),
.ZN(net2776)
);

AND2_X2 c2665(
.A1(net2774),
.A2(net1846),
.ZN(net2777)
);

XOR2_X1 c2666(
.A(net1593),
.B(net888),
.Z(net2778)
);

DFFS_X1 c2667(
.D(net767),
.SN(net2587),
.CK(clk),
.Q(net2780),
.QN(net2779)
);

DFFS_X2 c2668(
.D(net2778),
.SN(net1821),
.CK(clk),
.Q(net2782),
.QN(net2781)
);

NOR2_X1 c2669(
.A1(net870),
.A2(net877),
.ZN(net2783)
);

OR2_X2 c2670(
.A1(net2346),
.A2(net888),
.ZN(net2784)
);

NOR2_X4 c2671(
.A1(net927),
.A2(net1833),
.ZN(net2785)
);

NOR2_X2 c2672(
.A1(net2757),
.A2(net1784),
.ZN(net2786)
);

XOR2_X2 c2673(
.A(net921),
.B(net888),
.Z(net2787)
);

XNOR2_X1 c2674(
.A(net788),
.B(net1836),
.ZN(net2788)
);

OAI21_X4 c2675(
.A(net687),
.B1(net2745),
.B2(net902),
.ZN(net2789)
);

OR2_X4 c2676(
.A1(net889),
.A2(net2778),
.ZN(net2790)
);

OR2_X1 c2677(
.A1(net900),
.A2(net2772),
.ZN(net2791)
);

XNOR2_X2 c2678(
.A(net2773),
.B(net2786),
.ZN(net2792)
);

AND2_X4 c2679(
.A1(net1647),
.A2(net2774),
.ZN(net2793)
);

AND2_X1 c2680(
.A1(net2727),
.A2(net922),
.ZN(net2794)
);

NAND2_X1 c2681(
.A1(net1856),
.A2(net2771),
.ZN(net2795)
);

INV_X8 c2682(
.A(net2716),
.ZN(net2796)
);

NAND2_X2 c2683(
.A1(net2616),
.A2(net2771),
.ZN(net2797)
);

INV_X16 c2684(
.A(net10279),
.ZN(net2798)
);

NAND2_X4 c2685(
.A1(net1839),
.A2(net2789),
.ZN(net2799)
);

AND2_X2 c2686(
.A1(net1737),
.A2(net2784),
.ZN(net2800)
);

XOR2_X1 c2687(
.A(net2748),
.B(net2775),
.Z(net2801)
);

NOR2_X1 c2688(
.A1(net865),
.A2(net10401),
.ZN(net2802)
);

SDFF_X2 c2689(
.D(net2785),
.SE(net1844),
.SI(net1847),
.CK(clk),
.Q(net2804),
.QN(net2803)
);

OR2_X2 c2690(
.A1(net920),
.A2(net1784),
.ZN(net2805)
);

MUX2_X2 c2691(
.A(net1820),
.B(net2750),
.S(net1816),
.Z(net2806)
);

NOR2_X4 c2692(
.A1(net1864),
.A2(net2806),
.ZN(net2807)
);

NOR2_X2 c2693(
.A1(net888),
.A2(net2798),
.ZN(net2808)
);

XOR2_X2 c2694(
.A(net2801),
.B(net2799),
.Z(net2809)
);

XNOR2_X1 c2695(
.A(net914),
.B(net2806),
.ZN(net2810)
);

OAI221_X4 c2696(
.A(net2750),
.B1(net1843),
.B2(net1727),
.C1(net2799),
.C2(net2808),
.ZN(net2811)
);

DFFRS_X1 c2697(
.D(net2811),
.RN(net2787),
.SN(net914),
.CK(clk),
.Q(net2813),
.QN(net2812)
);

OR2_X4 c2698(
.A1(net1817),
.A2(net2812),
.ZN(net2814)
);

OR2_X1 c2699(
.A1(net811),
.A2(net1846),
.ZN(net2815)
);

XNOR2_X2 c2700(
.A(net2807),
.B(net870),
.ZN(net2816)
);

NAND3_X4 c2701(
.A1(net2729),
.A2(net2796),
.A3(net1736),
.ZN(net2817)
);

AND2_X4 c2702(
.A1(net897),
.A2(net1739),
.ZN(net2818)
);

SDFFRS_X2 c2703(
.D(net910),
.RN(net2587),
.SE(net2740),
.SI(net2774),
.SN(net1846),
.CK(clk),
.Q(net2820),
.QN(net2819)
);

CLKGATETST_X1 c2704(
.E(net2650),
.SE(net2817),
.CK(clk),
.GCK(net2821)
);

OR3_X4 c2705(
.A1(net2794),
.A2(net2821),
.A3(net851),
.ZN(net2822)
);

NAND4_X1 c2706(
.A1(net2818),
.A2(net1869),
.A3(net921),
.A4(net2809),
.ZN(net2823)
);

AND2_X1 c2707(
.A1(net2798),
.A2(net10763),
.ZN(net2824)
);

INV_X32 c2708(
.A(net9794),
.ZN(net2825)
);

INV_X4 c2709(
.A(net10272),
.ZN(net2826)
);

CLKGATETST_X2 c2710(
.E(net2790),
.SE(net2810),
.CK(clk),
.GCK(net2827)
);

NAND2_X1 c2711(
.A1(net2764),
.A2(net2824),
.ZN(net2828)
);

OR4_X1 c2712(
.A1(net2827),
.A2(net2806),
.A3(net1868),
.A4(net11165),
.ZN(net2829)
);

NAND2_X2 c2713(
.A1(net2719),
.A2(net2828),
.ZN(net2830)
);

CLKGATETST_X4 c2714(
.E(net1821),
.SE(net2829),
.CK(clk),
.GCK(net2831)
);

AND3_X2 c2715(
.A1(net837),
.A2(net1886),
.A3(net2807),
.ZN(net2832)
);

NOR3_X1 c2716(
.A1(net772),
.A2(net2824),
.A3(net902),
.ZN(net2833)
);

NAND2_X4 c2717(
.A1(net1677),
.A2(net2815),
.ZN(net2834)
);

OR3_X2 c2718(
.A1(net2792),
.A2(net1885),
.A3(net2695),
.ZN(net2835)
);

INV_X1 c2719(
.A(net10139),
.ZN(net2836)
);

AND2_X2 c2720(
.A1(net2745),
.A2(net2826),
.ZN(net2837)
);

XOR2_X1 c2721(
.A(net1574),
.B(net2776),
.Z(net2838)
);

SDFFR_X1 c2722(
.D(net2832),
.RN(net2834),
.SE(net2821),
.SI(net877),
.CK(clk),
.Q(net2840),
.QN(net2839)
);

NOR2_X1 c2723(
.A1(net2544),
.A2(net2783),
.ZN(net2841)
);

OR2_X2 c2724(
.A1(net2841),
.A2(net2558),
.ZN(net2842)
);

DFFRS_X2 c2725(
.D(net2842),
.RN(net2834),
.SN(net2839),
.CK(clk),
.Q(net2844),
.QN(net2843)
);

OAI221_X2 c2726(
.A(net2797),
.B1(net914),
.B2(net2837),
.C1(net2843),
.C2(net2821),
.ZN(net2845)
);

INV_X2 c2727(
.A(net9643),
.ZN(net2846)
);

OAI21_X2 c2728(
.A(net2816),
.B1(net2802),
.B2(net1677),
.ZN(net2847)
);

NOR2_X4 c2729(
.A1(net2843),
.A2(net10601),
.ZN(net2848)
);

NOR2_X2 c2730(
.A1(net2788),
.A2(net2847),
.ZN(net2849)
);

OAI21_X1 c2731(
.A(net1727),
.B1(net2844),
.B2(net2835),
.ZN(net2850)
);

XOR2_X2 c2732(
.A(net1627),
.B(net10601),
.Z(net2851)
);

SDFF_X1 c2733(
.D(net2829),
.SE(net1857),
.SI(net2851),
.CK(clk),
.Q(net2853),
.QN(net2852)
);

OAI22_X1 c2734(
.A1(net1814),
.A2(net2819),
.B1(net2834),
.B2(net2851),
.ZN(net2854)
);

AOI21_X2 c2735(
.A(net2824),
.B1(net2837),
.B2(net2848),
.ZN(net2855)
);

AOI21_X1 c2736(
.A(net2855),
.B1(net2846),
.B2(net2852),
.ZN(net2856)
);

AOI21_X4 c2737(
.A(net2856),
.B1(net2850),
.B2(net2716),
.ZN(net2857)
);

OAI222_X4 c2738(
.A1(net1784),
.A2(net2856),
.B1(net2851),
.B2(net851),
.C1(net2834),
.C2(net10400),
.ZN(net2858)
);

INV_X8 c2739(
.A(net1971),
.ZN(net2859)
);

INV_X16 c2740(
.A(net1946),
.ZN(net2860)
);

INV_X32 c2741(
.A(net951),
.ZN(net2861)
);

CLKGATETST_X8 c2742(
.E(in24),
.SE(net1010),
.CK(clk),
.GCK(net2862)
);

INV_X4 c2743(
.A(net2861),
.ZN(net2863)
);

INV_X1 c2744(
.A(net1906),
.ZN(net2864)
);

INV_X2 c2745(
.A(net2860),
.ZN(net2865)
);

INV_X8 c2746(
.A(net2859),
.ZN(net2866)
);

XNOR2_X1 c2747(
.A(net948),
.B(net11158),
.ZN(net2867)
);

OR2_X4 c2748(
.A1(net956),
.A2(net2861),
.ZN(net2868)
);

OR2_X1 c2749(
.A1(net1900),
.A2(in7),
.ZN(net2869)
);

XNOR2_X2 c2750(
.A(net1932),
.B(net1966),
.ZN(net2870)
);

INV_X16 c2751(
.A(net14),
.ZN(net2871)
);

INV_X32 c2752(
.A(net957),
.ZN(net2872)
);

AND2_X4 c2753(
.A1(net951),
.A2(net1954),
.ZN(net2873)
);

AND3_X1 c2754(
.A1(net2866),
.A2(net2867),
.A3(net2872),
.ZN(net2874)
);

AND2_X1 c2755(
.A1(net2869),
.A2(net1909),
.ZN(net2875)
);

INV_X4 c2756(
.A(net2869),
.ZN(net2876)
);

INV_X1 c2757(
.A(net1922),
.ZN(net2877)
);

NAND2_X1 c2758(
.A1(net2872),
.A2(net11159),
.ZN(net2878)
);

NAND2_X2 c2759(
.A1(net2878),
.A2(net2860),
.ZN(net2879)
);

INV_X2 c2760(
.A(net993),
.ZN(net2880)
);

NAND3_X1 c2761(
.A1(net2877),
.A2(net1906),
.A3(net988),
.ZN(net2881)
);

INV_X8 c2762(
.A(net1954),
.ZN(net2882)
);

INV_X16 c2763(
.A(net1952),
.ZN(net2883)
);

NOR3_X4 c2764(
.A1(net2873),
.A2(net2880),
.A3(net33),
.ZN(net2884)
);

NAND2_X4 c2765(
.A1(net1971),
.A2(net2878),
.ZN(net2885)
);

INV_X32 c2766(
.A(net9555),
.ZN(net2886)
);

DFFR_X1 c2767(
.D(net2881),
.RN(net1912),
.CK(clk),
.Q(net2888),
.QN(net2887)
);

INV_X4 c2768(
.A(net9556),
.ZN(net2889)
);

NOR3_X2 c2769(
.A1(net2889),
.A2(net2875),
.A3(in24),
.ZN(net2890)
);

INV_X1 c2770(
.A(net1906),
.ZN(net2891)
);

AND2_X2 c2771(
.A1(net2872),
.A2(net1942),
.ZN(net2892)
);

AND3_X4 c2772(
.A1(net2890),
.A2(net2876),
.A3(net2882),
.ZN(net2893)
);

XOR2_X1 c2773(
.A(net2868),
.B(net2862),
.Z(net2894)
);

INV_X2 c2774(
.A(net2867),
.ZN(net2895)
);

NOR2_X1 c2775(
.A1(net1906),
.A2(net10524),
.ZN(net2896)
);

OR2_X2 c2776(
.A1(net2894),
.A2(net976),
.ZN(net2897)
);

INV_X8 c2777(
.A(net2886),
.ZN(net2898)
);

NOR2_X4 c2778(
.A1(net1967),
.A2(net1922),
.ZN(net2899)
);

INV_X16 c2779(
.A(net993),
.ZN(net2900)
);

NOR2_X2 c2780(
.A1(net2876),
.A2(net2865),
.ZN(net2901)
);

XOR2_X2 c2781(
.A(net2864),
.B(net2875),
.Z(net2902)
);

INV_X32 c2782(
.A(net2870),
.ZN(net2903)
);

INV_X4 c2783(
.A(net2878),
.ZN(net2904)
);

XNOR2_X1 c2784(
.A(net2883),
.B(net2886),
.ZN(net2905)
);

OR2_X4 c2785(
.A1(net2901),
.A2(net2889),
.ZN(net2906)
);

OR2_X1 c2786(
.A1(net2906),
.A2(net10489),
.ZN(net2907)
);

XNOR2_X2 c2787(
.A(net1909),
.B(net10489),
.ZN(net2908)
);

INV_X1 c2788(
.A(net2874),
.ZN(net2909)
);

AND2_X4 c2789(
.A1(net2908),
.A2(net2902),
.ZN(net2910)
);

INV_X2 c2790(
.A(net2907),
.ZN(net2911)
);

SDFF_X2 c2791(
.D(net2895),
.SE(net2885),
.SI(net2887),
.CK(clk),
.Q(net2913),
.QN(net2912)
);

AND2_X1 c2792(
.A1(net2903),
.A2(net2892),
.ZN(net2914)
);

NAND3_X2 c2793(
.A1(net2896),
.A2(net2886),
.A3(net2889),
.ZN(net2915)
);

DFFR_X2 c2794(
.D(net2904),
.RN(net2888),
.CK(clk),
.Q(net2917),
.QN(net2916)
);

DFFRS_X1 c2795(
.D(net2913),
.RN(net2903),
.SN(net2914),
.CK(clk),
.Q(net2919),
.QN(net2918)
);

NAND2_X1 c2796(
.A1(net1896),
.A2(net2911),
.ZN(net2920)
);

DFFRS_X2 c2797(
.D(net2875),
.RN(net2909),
.SN(net2868),
.CK(clk),
.Q(net2922),
.QN(net2921)
);

NAND2_X2 c2798(
.A1(net2892),
.A2(net2881),
.ZN(net2923)
);

SDFF_X1 c2799(
.D(net2906),
.SE(net2919),
.SI(net2914),
.CK(clk),
.Q(net2925),
.QN(net2924)
);

DFFS_X1 c2800(
.D(net2915),
.SN(net2923),
.CK(clk),
.Q(net2927),
.QN(net2926)
);

NAND2_X4 c2801(
.A1(net2902),
.A2(net948),
.ZN(net2928)
);

SDFF_X2 c2802(
.D(net2888),
.SE(net2909),
.SI(net2912),
.CK(clk),
.Q(net2930),
.QN(net2929)
);

OR3_X1 c2803(
.A1(net2899),
.A2(net2926),
.A3(net2886),
.ZN(net2931)
);

MUX2_X1 c2804(
.A(net2911),
.B(net2866),
.S(net2924),
.Z(net2932)
);

OAI21_X4 c2805(
.A(net2893),
.B1(net2900),
.B2(net2873),
.ZN(net2933)
);

MUX2_X2 c2806(
.A(net2880),
.B(net2925),
.S(net2929),
.Z(net2934)
);

AND2_X2 c2807(
.A1(net2877),
.A2(net2870),
.ZN(net2935)
);

AND4_X2 c2808(
.A1(net2925),
.A2(net2931),
.A3(net2871),
.A4(net1891),
.ZN(net2936)
);

DFFRS_X1 c2809(
.D(net2909),
.RN(net2931),
.SN(net2933),
.CK(clk),
.Q(net2938),
.QN(net2937)
);

XOR2_X1 c2810(
.A(net2891),
.B(net2933),
.Z(net2939)
);

NOR2_X1 c2811(
.A1(net2931),
.A2(net1954),
.ZN(net2940)
);

NAND3_X4 c2812(
.A1(net2930),
.A2(net2937),
.A3(net2934),
.ZN(net2941)
);

OR2_X2 c2813(
.A1(net2933),
.A2(net2935),
.ZN(net2942)
);

NOR2_X4 c2814(
.A1(net2890),
.A2(net2934),
.ZN(net2943)
);

DFFS_X2 c2815(
.D(net1010),
.SN(net1950),
.CK(clk),
.Q(net2945),
.QN(net2944)
);

NOR2_X2 c2816(
.A1(net2934),
.A2(net2940),
.ZN(net2946)
);

DFFRS_X2 c2817(
.D(net1946),
.RN(net2915),
.SN(net2914),
.CK(clk),
.Q(net2948),
.QN(net2947)
);

XOR2_X2 c2818(
.A(net2938),
.B(net2940),
.Z(net2949)
);

AOI221_X4 c2819(
.A(net2895),
.B1(net2886),
.B2(net2933),
.C1(net2920),
.C2(net2943),
.ZN(net2950)
);

SDFFRS_X1 c2820(
.D(net2949),
.RN(net2933),
.SE(net2944),
.SI(net2943),
.SN(net2936),
.CK(clk),
.Q(net2952),
.QN(net2951)
);

XNOR2_X1 c2821(
.A(net2949),
.B(net10489),
.ZN(net2953)
);

OR2_X4 c2822(
.A1(net2871),
.A2(net2047),
.ZN(net2954)
);

INV_X8 c2823(
.A(net1025),
.ZN(net2955)
);

INV_X16 c2824(
.A(net2928),
.ZN(net2956)
);

CLKGATETST_X1 c2825(
.E(net1093),
.SE(net1988),
.CK(clk),
.GCK(net2957)
);

INV_X32 c2826(
.A(net1053),
.ZN(net2958)
);

INV_X4 c2827(
.A(net2945),
.ZN(net2959)
);

OR2_X1 c2828(
.A1(net1942),
.A2(net2897),
.ZN(net2960)
);

INV_X1 c2829(
.A(net1999),
.ZN(net2961)
);

INV_X2 c2830(
.A(net1038),
.ZN(net2962)
);

INV_X8 c2831(
.A(net9572),
.ZN(net2963)
);

INV_X16 c2832(
.A(net2952),
.ZN(net2964)
);

INV_X32 c2833(
.A(net10717),
.ZN(net2965)
);

INV_X4 c2834(
.A(net2917),
.ZN(net2966)
);

INV_X1 c2835(
.A(net10470),
.ZN(net2967)
);

INV_X2 c2836(
.A(net1992),
.ZN(net2968)
);

INV_X8 c2837(
.A(net2900),
.ZN(net2969)
);

INV_X16 c2838(
.A(net2958),
.ZN(net2970)
);

INV_X32 c2839(
.A(net2968),
.ZN(net2971)
);

INV_X4 c2840(
.A(net2967),
.ZN(net2972)
);

XNOR2_X2 c2841(
.A(net2941),
.B(net2956),
.ZN(net2973)
);

INV_X1 c2842(
.A(net2948),
.ZN(net2974)
);

INV_X2 c2843(
.A(net9571),
.ZN(net2975)
);

INV_X8 c2844(
.A(net29),
.ZN(net2976)
);

INV_X16 c2845(
.A(net2970),
.ZN(net2977)
);

AND2_X4 c2846(
.A1(net2897),
.A2(net2970),
.ZN(net2978)
);

AND2_X1 c2847(
.A1(net2961),
.A2(net979),
.ZN(net2979)
);

INV_X32 c2848(
.A(net2927),
.ZN(net2980)
);

NAND2_X1 c2849(
.A1(net2041),
.A2(net2970),
.ZN(net2981)
);

OR3_X4 c2850(
.A1(net2027),
.A2(net2976),
.A3(net2947),
.ZN(net2982)
);

AND3_X2 c2851(
.A1(net2865),
.A2(net2957),
.A3(net2976),
.ZN(net2983)
);

NOR3_X1 c2852(
.A1(net2971),
.A2(net2064),
.A3(net1985),
.ZN(net2984)
);

NAND2_X2 c2853(
.A1(net2980),
.A2(net1927),
.ZN(net2985)
);

NAND2_X4 c2854(
.A1(net2967),
.A2(net2038),
.ZN(net2986)
);

INV_X4 c2855(
.A(net2976),
.ZN(net2987)
);

AND2_X2 c2856(
.A1(net2062),
.A2(net2920),
.ZN(net2988)
);

INV_X1 c2857(
.A(net2057),
.ZN(net2989)
);

INV_X2 c2858(
.A(net2969),
.ZN(net2990)
);

INV_X8 c2859(
.A(net9772),
.ZN(net2991)
);

INV_X16 c2860(
.A(net2962),
.ZN(net2992)
);

OR3_X2 c2861(
.A1(net2987),
.A2(net2970),
.A3(net1908),
.ZN(net2993)
);

INV_X32 c2862(
.A(net9754),
.ZN(net2994)
);

XOR2_X1 c2863(
.A(net2992),
.B(net77),
.Z(net2995)
);

INV_X4 c2864(
.A(net2979),
.ZN(net2996)
);

INV_X1 c2865(
.A(net2995),
.ZN(net2997)
);

INV_X2 c2866(
.A(net2975),
.ZN(net2998)
);

CLKGATETST_X2 c2867(
.E(net2985),
.SE(net2914),
.CK(clk),
.GCK(net2999)
);

CLKGATETST_X4 c2868(
.E(net2981),
.SE(net2046),
.CK(clk),
.GCK(net3000)
);

NOR2_X1 c2869(
.A1(net2996),
.A2(net2991),
.ZN(net3001)
);

OR2_X2 c2870(
.A1(net2974),
.A2(net10500),
.ZN(net3002)
);

NOR2_X4 c2871(
.A1(net2955),
.A2(net2991),
.ZN(net3003)
);

NOR2_X2 c2872(
.A1(net2989),
.A2(net3000),
.ZN(net3004)
);

INV_X8 c2873(
.A(net2997),
.ZN(net3005)
);

INV_X16 c2874(
.A(net9745),
.ZN(net3006)
);

XOR2_X2 c2875(
.A(net2984),
.B(net2974),
.Z(net3007)
);

INV_X32 c2876(
.A(net1932),
.ZN(net3008)
);

INV_X4 c2877(
.A(net3005),
.ZN(net3009)
);

XNOR2_X1 c2878(
.A(net2966),
.B(net2996),
.ZN(net3010)
);

SDFFR_X2 c2879(
.D(net3002),
.RN(net1102),
.SE(net2015),
.SI(net2993),
.CK(clk),
.Q(net3012),
.QN(net3011)
);

OR2_X4 c2880(
.A1(net2963),
.A2(net2916),
.ZN(net3013)
);

OR2_X1 c2881(
.A1(net3004),
.A2(net2991),
.ZN(net3014)
);

XNOR2_X2 c2882(
.A(net974),
.B(net2036),
.ZN(net3015)
);

INV_X1 c2883(
.A(net9972),
.ZN(net3016)
);

AND2_X4 c2884(
.A1(net3008),
.A2(net3012),
.ZN(net3017)
);

AND2_X1 c2885(
.A1(net2956),
.A2(net3017),
.ZN(net3018)
);

OAI21_X2 c2886(
.A(net3018),
.B1(net3006),
.B2(net2047),
.ZN(net3019)
);

NAND2_X1 c2887(
.A1(net2994),
.A2(net3017),
.ZN(net3020)
);

OAI21_X1 c2888(
.A(net2954),
.B1(net2986),
.B2(net2991),
.ZN(net3021)
);

NAND2_X2 c2889(
.A1(net1951),
.A2(net3020),
.ZN(net3022)
);

AOI21_X2 c2890(
.A(net3021),
.B1(net2990),
.B2(net2862),
.ZN(net3023)
);

NAND2_X4 c2891(
.A1(net3006),
.A2(net3022),
.ZN(net3024)
);

CLKGATETST_X8 c2892(
.E(net2957),
.SE(net2051),
.CK(clk),
.GCK(net3025)
);

AND2_X2 c2893(
.A1(net2015),
.A2(net3014),
.ZN(net3026)
);

AOI21_X1 c2894(
.A(net3019),
.B1(net2001),
.B2(net3020),
.ZN(net3027)
);

XOR2_X1 c2895(
.A(net2991),
.B(net10628),
.Z(net3028)
);

SDFF_X1 c2896(
.D(net2010),
.SE(net3024),
.SI(net2918),
.CK(clk),
.Q(net3030),
.QN(net3029)
);

NOR2_X1 c2897(
.A1(net3027),
.A2(net2983),
.ZN(net3031)
);

OR2_X2 c2898(
.A1(net3030),
.A2(net3025),
.ZN(net3032)
);

AOI21_X4 c2899(
.A(net2005),
.B1(net3025),
.B2(net3032),
.ZN(net3033)
);

AND4_X1 c2900(
.A1(net3033),
.A2(net2977),
.A3(net3025),
.A4(net3032),
.ZN(net3034)
);

NOR2_X4 c2901(
.A1(net3029),
.A2(net10540),
.ZN(net3035)
);

OAI222_X2 c2902(
.A1(net3032),
.A2(net3025),
.B1(net3000),
.B2(net3024),
.C1(net3016),
.C2(net2959),
.ZN(net3036)
);

AOI222_X1 c2903(
.A1(net3028),
.A2(net3011),
.B1(net2972),
.B2(net3026),
.C1(net1968),
.C2(net3036),
.ZN(net3037)
);

AND3_X1 c2904(
.A1(net3010),
.A2(net3032),
.A3(net3036),
.ZN(net3038)
);

NOR2_X2 c2905(
.A1(net2999),
.A2(net3036),
.ZN(net3039)
);

AOI22_X4 c2906(
.A1(net2138),
.A2(net2953),
.B1(net2147),
.B2(net33),
.ZN(net3040)
);

INV_X2 c2907(
.A(net2069),
.ZN(net3041)
);

INV_X8 c2908(
.A(net2082),
.ZN(net3042)
);

INV_X16 c2909(
.A(net9661),
.ZN(net3043)
);

XOR2_X2 c2910(
.A(net3009),
.B(net2860),
.Z(net3044)
);

INV_X32 c2911(
.A(net9661),
.ZN(net3045)
);

INV_X4 c2912(
.A(net3042),
.ZN(net3046)
);

XNOR2_X1 c2913(
.A(net3041),
.B(net2090),
.ZN(net3047)
);

NAND3_X1 c2914(
.A1(net2132),
.A2(net1139),
.A3(net2974),
.ZN(net3048)
);

INV_X1 c2915(
.A(net2094),
.ZN(net3049)
);

INV_X2 c2916(
.A(net2022),
.ZN(net3050)
);

OR2_X4 c2917(
.A1(net3050),
.A2(net1177),
.ZN(net3051)
);

OR2_X1 c2918(
.A1(net3049),
.A2(net2022),
.ZN(net3052)
);

XNOR2_X2 c2919(
.A(net3046),
.B(net3020),
.ZN(net3053)
);

INV_X8 c2920(
.A(net10743),
.ZN(net3054)
);

INV_X16 c2921(
.A(net10985),
.ZN(net3055)
);

INV_X32 c2922(
.A(net3053),
.ZN(net3056)
);

AND2_X4 c2923(
.A1(net2139),
.A2(net2056),
.ZN(net3057)
);

INV_X4 c2924(
.A(net2047),
.ZN(net3058)
);

INV_X1 c2925(
.A(net2151),
.ZN(net3059)
);

INV_X2 c2926(
.A(net11041),
.ZN(net3060)
);

AND2_X1 c2927(
.A1(net3047),
.A2(net3056),
.ZN(net3061)
);

NAND2_X1 c2928(
.A1(net3024),
.A2(net2139),
.ZN(net3062)
);

INV_X8 c2929(
.A(net10898),
.ZN(net3063)
);

INV_X16 c2930(
.A(net3052),
.ZN(net3064)
);

INV_X32 c2931(
.A(net3062),
.ZN(net3065)
);

INV_X4 c2932(
.A(net3055),
.ZN(net3066)
);

INV_X1 c2933(
.A(net3063),
.ZN(net3067)
);

NAND2_X2 c2934(
.A1(net3067),
.A2(net3026),
.ZN(net3068)
);

INV_X2 c2935(
.A(net3061),
.ZN(net3069)
);

NAND2_X4 c2936(
.A1(net1139),
.A2(net2151),
.ZN(net3070)
);

INV_X8 c2937(
.A(net11084),
.ZN(net3071)
);

AND2_X2 c2938(
.A1(net2019),
.A2(net1968),
.ZN(net3072)
);

INV_X16 c2939(
.A(net10536),
.ZN(net3073)
);

XOR2_X1 c2940(
.A(net1153),
.B(net3064),
.Z(net3074)
);

INV_X32 c2941(
.A(net3054),
.ZN(net3075)
);

NOR2_X1 c2942(
.A1(net2863),
.A2(net10950),
.ZN(net3076)
);

OR2_X2 c2943(
.A1(net3073),
.A2(net2999),
.ZN(net3077)
);

INV_X4 c2944(
.A(net1968),
.ZN(net3078)
);

INV_X1 c2945(
.A(net9700),
.ZN(net3079)
);

NOR2_X4 c2946(
.A1(net3075),
.A2(net3072),
.ZN(net3080)
);

NOR2_X2 c2947(
.A1(net3043),
.A2(net2147),
.ZN(net3081)
);

XOR2_X2 c2948(
.A(net3020),
.B(net3080),
.Z(net3082)
);

XNOR2_X1 c2949(
.A(net2953),
.B(net3081),
.ZN(net3083)
);

INV_X2 c2950(
.A(net3082),
.ZN(net3084)
);

INV_X8 c2951(
.A(net3003),
.ZN(net3085)
);

OR2_X4 c2952(
.A1(net2914),
.A2(net185),
.ZN(net3086)
);

INV_X16 c2953(
.A(net10868),
.ZN(net3087)
);

INV_X32 c2954(
.A(net10806),
.ZN(net3088)
);

INV_X4 c2955(
.A(net10770),
.ZN(net3089)
);

NOR3_X4 c2956(
.A1(net3079),
.A2(net3078),
.A3(net3080),
.ZN(net3090)
);

OR2_X1 c2957(
.A1(net3090),
.A2(net3089),
.ZN(net3091)
);

XNOR2_X2 c2958(
.A(net3080),
.B(net3073),
.ZN(net3092)
);

NOR3_X2 c2959(
.A1(net3087),
.A2(net3065),
.A3(net3026),
.ZN(net3093)
);

AND2_X4 c2960(
.A1(net3089),
.A2(net3056),
.ZN(net3094)
);

INV_X1 c2961(
.A(net1085),
.ZN(net3095)
);

AND2_X1 c2962(
.A1(net3088),
.A2(net3079),
.ZN(net3096)
);

NAND2_X1 c2963(
.A1(net3058),
.A2(net3065),
.ZN(net3097)
);

NAND2_X2 c2964(
.A1(net3077),
.A2(net3081),
.ZN(net3098)
);

NAND2_X4 c2965(
.A1(net1034),
.A2(net3081),
.ZN(net3099)
);

AND2_X2 c2966(
.A1(net3083),
.A2(net3077),
.ZN(net3100)
);

INV_X2 c2967(
.A(net10851),
.ZN(net3101)
);

INV_X8 c2968(
.A(net9971),
.ZN(net3102)
);

AND3_X4 c2969(
.A1(net3057),
.A2(net3024),
.A3(net3060),
.ZN(net3103)
);

NAND3_X2 c2970(
.A1(net2974),
.A2(net3102),
.A3(net2978),
.ZN(net3104)
);

XOR2_X1 c2971(
.A(net1129),
.B(net2129),
.Z(net3105)
);

AOI221_X2 c2972(
.A(net3105),
.B1(net2151),
.B2(net2953),
.C1(net2112),
.C2(net3081),
.ZN(net3106)
);

NOR2_X1 c2973(
.A1(net3065),
.A2(net3106),
.ZN(net3107)
);

INV_X16 c2974(
.A(net3100),
.ZN(net3108)
);

OR2_X2 c2975(
.A1(net3092),
.A2(net3102),
.ZN(net3109)
);

OAI22_X4 c2976(
.A1(net183),
.A2(net3106),
.B1(net3108),
.B2(net2147),
.ZN(net3110)
);

NOR2_X4 c2977(
.A1(net3099),
.A2(net3072),
.ZN(net3111)
);

NOR2_X2 c2978(
.A1(net3093),
.A2(net3107),
.ZN(net3112)
);

INV_X32 c2979(
.A(net10976),
.ZN(net3113)
);

SDFF_X2 c2980(
.D(net3026),
.SE(net3091),
.SI(net3108),
.CK(clk),
.Q(net3115),
.QN(net3114)
);

OR3_X1 c2981(
.A1(net3097),
.A2(net3101),
.A3(net3114),
.ZN(net3116)
);

MUX2_X1 c2982(
.A(net3103),
.B(net1891),
.S(net3097),
.Z(net3117)
);

AOI221_X1 c2983(
.A(net3068),
.B1(net3085),
.B2(net3094),
.C1(net3080),
.C2(net3060),
.ZN(net3118)
);

OAI221_X1 c2984(
.A(net3059),
.B1(net3085),
.B2(net3113),
.C1(net3035),
.C2(net3060),
.ZN(net3119)
);

OAI21_X4 c2985(
.A(net3095),
.B1(net3102),
.B2(net3089),
.ZN(net3120)
);

DFFRS_X1 c2986(
.D(net3112),
.RN(net3080),
.SN(net10501),
.CK(clk),
.Q(net3122),
.QN(net3121)
);

MUX2_X2 c2987(
.A(net3111),
.B(net3100),
.S(net3122),
.Z(net3123)
);

XOR2_X2 c2988(
.A(net2231),
.B(net2137),
.Z(net3124)
);

XNOR2_X1 c2989(
.A(net3066),
.B(net2195),
.ZN(net3125)
);

INV_X4 c2990(
.A(net3022),
.ZN(net3126)
);

INV_X1 c2991(
.A(net2165),
.ZN(net3127)
);

OR2_X4 c2992(
.A1(net2060),
.A2(net2206),
.ZN(net3128)
);

OR2_X1 c2993(
.A1(net265),
.A2(net1212),
.ZN(net3129)
);

XNOR2_X2 c2994(
.A(net3127),
.B(net2157),
.ZN(net3130)
);

INV_X2 c2995(
.A(net3096),
.ZN(net3131)
);

INV_X8 c2996(
.A(net3094),
.ZN(net3132)
);

AND2_X4 c2997(
.A1(net1270),
.A2(net10949),
.ZN(net3133)
);

INV_X16 c2998(
.A(net10137),
.ZN(net3134)
);

INV_X32 c2999(
.A(net11003),
.ZN(net3135)
);

NAND3_X4 c3000(
.A1(net3132),
.A2(net3094),
.A3(net3121),
.ZN(net3136)
);

AND2_X1 c3001(
.A1(net2137),
.A2(net3022),
.ZN(net3137)
);

OR3_X4 c3002(
.A1(net3124),
.A2(net1212),
.A3(net11012),
.ZN(net3138)
);

NAND2_X1 c3003(
.A1(net1898),
.A2(net3115),
.ZN(net3139)
);

NAND2_X2 c3004(
.A1(net2160),
.A2(net77),
.ZN(net3140)
);

NAND2_X4 c3005(
.A1(net1022),
.A2(net3123),
.ZN(net3141)
);

AND2_X2 c3006(
.A1(net3137),
.A2(net3134),
.ZN(net3142)
);

INV_X4 c3007(
.A(net11003),
.ZN(net3143)
);

XOR2_X1 c3008(
.A(net2164),
.B(net1203),
.Z(net3144)
);

INV_X1 c3009(
.A(net3128),
.ZN(net3145)
);

NOR2_X1 c3010(
.A1(net3098),
.A2(net1995),
.ZN(net3146)
);

OR2_X2 c3011(
.A1(net2206),
.A2(net10973),
.ZN(net3147)
);

NOR2_X4 c3012(
.A1(net2223),
.A2(net2165),
.ZN(net3148)
);

NOR2_X2 c3013(
.A1(net3148),
.A2(net1270),
.ZN(net3149)
);

INV_X2 c3014(
.A(net10202),
.ZN(net3150)
);

DFFR_X1 c3015(
.D(net3109),
.RN(net3150),
.CK(clk),
.Q(net3152),
.QN(net3151)
);

INV_X8 c3016(
.A(net10360),
.ZN(net3153)
);

XOR2_X2 c3017(
.A(net2206),
.B(net3114),
.Z(net3154)
);

INV_X16 c3018(
.A(net3135),
.ZN(net3155)
);

INV_X32 c3019(
.A(net11015),
.ZN(net3156)
);

AND3_X2 c3020(
.A1(net987),
.A2(net3110),
.A3(net3119),
.ZN(net3157)
);

DFFRS_X2 c3021(
.D(net3106),
.RN(net2209),
.SN(net10875),
.CK(clk),
.Q(net3159),
.QN(net3158)
);

XNOR2_X1 c3022(
.A(net1179),
.B(net278),
.ZN(net3160)
);

INV_X4 c3023(
.A(net9863),
.ZN(net3161)
);

INV_X1 c3024(
.A(net10840),
.ZN(net3162)
);

OR2_X4 c3025(
.A1(net3133),
.A2(net10973),
.ZN(net3163)
);

INV_X2 c3026(
.A(net10974),
.ZN(net3164)
);

OAI221_X4 c3027(
.A(net3155),
.B1(net3154),
.B2(net3114),
.C1(net2959),
.C2(net2160),
.ZN(net3165)
);

OR2_X1 c3028(
.A1(net2157),
.A2(net3165),
.ZN(net3166)
);

XNOR2_X2 c3029(
.A(net3140),
.B(net3162),
.ZN(net3167)
);

AND2_X4 c3030(
.A1(net3156),
.A2(net3035),
.ZN(net3168)
);

AND2_X1 c3031(
.A1(net2860),
.A2(net3108),
.ZN(net3169)
);

SDFFRS_X2 c3032(
.D(net3142),
.RN(net276),
.SE(net3169),
.SI(net3153),
.SN(net11012),
.CK(clk),
.Q(net3171),
.QN(net3170)
);

INV_X8 c3033(
.A(net185),
.ZN(net3172)
);

NAND2_X1 c3034(
.A1(net2242),
.A2(net3168),
.ZN(net3173)
);

NAND2_X2 c3035(
.A1(net3154),
.A2(net3150),
.ZN(net3174)
);

NAND2_X4 c3036(
.A1(net3035),
.A2(net3170),
.ZN(net3175)
);

NOR3_X1 c3037(
.A1(net3164),
.A2(net2112),
.A3(net1988),
.ZN(net3176)
);

AND2_X2 c3038(
.A1(net3165),
.A2(net3158),
.ZN(net3177)
);

OR3_X2 c3039(
.A1(net3173),
.A2(net2206),
.A3(net3175),
.ZN(net3178)
);

XOR2_X1 c3040(
.A(net3172),
.B(net3171),
.Z(net3179)
);

NOR2_X1 c3041(
.A1(net3146),
.A2(net3152),
.ZN(net3180)
);

OAI21_X2 c3042(
.A(net3176),
.B1(net3169),
.B2(net3153),
.ZN(net3181)
);

OR2_X2 c3043(
.A1(net3125),
.A2(net1235),
.ZN(net3182)
);

NOR2_X4 c3044(
.A1(net3078),
.A2(net3172),
.ZN(net3183)
);

NOR2_X2 c3045(
.A1(net3167),
.A2(net3123),
.ZN(net3184)
);

XOR2_X2 c3046(
.A(net3174),
.B(net3164),
.Z(net3185)
);

OAI21_X1 c3047(
.A(net3182),
.B1(net3158),
.B2(net10920),
.ZN(net3186)
);

AOI21_X2 c3048(
.A(net2001),
.B1(net3165),
.B2(net3098),
.ZN(net3187)
);

AOI21_X1 c3049(
.A(net1235),
.B1(net3183),
.B2(net3153),
.ZN(net3188)
);

XNOR2_X1 c3050(
.A(net3147),
.B(net3187),
.ZN(net3189)
);

INV_X16 c3051(
.A(net10821),
.ZN(net3190)
);

AOI21_X4 c3052(
.A(net3186),
.B1(net2038),
.B2(net3190),
.ZN(net3191)
);

SDFFRS_X1 c3053(
.D(net3162),
.RN(net3169),
.SE(net3022),
.SI(net2160),
.SN(net3081),
.CK(clk),
.Q(net3193),
.QN(net3192)
);

SDFF_X1 c3054(
.D(net3179),
.SE(net3193),
.SI(net3189),
.CK(clk),
.Q(net3195),
.QN(net3194)
);

AND3_X1 c3055(
.A1(net3139),
.A2(net3172),
.A3(net3125),
.ZN(net3196)
);

OR2_X4 c3056(
.A1(net3185),
.A2(net3168),
.ZN(net3197)
);

OAI221_X2 c3057(
.A(net3196),
.B1(net3182),
.B2(net3180),
.C1(net3134),
.C2(net3194),
.ZN(net3198)
);

OR2_X1 c3058(
.A1(net3180),
.A2(net10920),
.ZN(net3199)
);

NAND3_X1 c3059(
.A1(net3191),
.A2(net3129),
.A3(net3035),
.ZN(net3200)
);

SDFF_X2 c3060(
.D(net3188),
.SE(net3199),
.SI(net2860),
.CK(clk),
.Q(net3202),
.QN(net3201)
);

SDFFRS_X2 c3061(
.D(net3150),
.RN(net3156),
.SE(net1235),
.SI(net3192),
.SN(net3169),
.CK(clk),
.Q(net3204),
.QN(net3203)
);

NOR3_X4 c3062(
.A1(net3183),
.A2(net3122),
.A3(net3175),
.ZN(net3205)
);

AOI222_X4 c3063(
.A1(net3202),
.A2(net3190),
.B1(net3188),
.B2(net3194),
.C1(net3007),
.C2(net3153),
.ZN(net3206)
);

NOR3_X2 c3064(
.A1(net3171),
.A2(net3202),
.A3(net3189),
.ZN(net3207)
);

AND3_X4 c3065(
.A1(net3177),
.A2(net3094),
.A3(net3183),
.ZN(net3208)
);

DFFR_X2 c3066(
.D(net3206),
.RN(net3189),
.CK(clk),
.Q(net3210),
.QN(net3209)
);

INV_X32 c3067(
.A(net10978),
.ZN(net3211)
);

OAI33_X1 c3068(
.A1(net3166),
.A2(net3204),
.A3(net1891),
.B1(net3208),
.B2(net3211),
.B3(net3201),
.ZN(net3212)
);

XNOR2_X2 c3069(
.A(net3131),
.B(net3211),
.ZN(net3213)
);

AOI222_X2 c3070(
.A1(net3198),
.A2(net3120),
.B1(net3209),
.B2(net3211),
.C1(net3150),
.C2(net11028),
.ZN(net3214)
);

INV_X4 c3071(
.A(net2299),
.ZN(net3215)
);

INV_X1 c3072(
.A(net11125),
.ZN(net3216)
);

INV_X2 c3073(
.A(net10821),
.ZN(net3217)
);

INV_X8 c3074(
.A(net2208),
.ZN(net3218)
);

INV_X16 c3075(
.A(net3076),
.ZN(net3219)
);

AND2_X4 c3076(
.A1(net2273),
.A2(net3192),
.ZN(net3220)
);

INV_X32 c3077(
.A(net2147),
.ZN(net3221)
);

NAND3_X2 c3078(
.A1(net365),
.A2(net1995),
.A3(net2203),
.ZN(net3222)
);

AND2_X1 c3079(
.A1(net345),
.A2(net2293),
.ZN(net3223)
);

INV_X4 c3080(
.A(net2294),
.ZN(net3224)
);

NAND2_X1 c3081(
.A1(net2320),
.A2(net2222),
.ZN(net3225)
);

NAND2_X2 c3082(
.A1(net2313),
.A2(net1995),
.ZN(net3226)
);

INV_X1 c3083(
.A(net1332),
.ZN(net3227)
);

INV_X2 c3084(
.A(net9557),
.ZN(net3228)
);

NAND2_X4 c3085(
.A1(net2305),
.A2(net3194),
.ZN(net3229)
);

AND2_X2 c3086(
.A1(net3193),
.A2(net3129),
.ZN(net3230)
);

XOR2_X1 c3087(
.A(net3223),
.B(net2203),
.Z(net3231)
);

INV_X8 c3088(
.A(net3218),
.ZN(net3232)
);

INV_X16 c3089(
.A(net3224),
.ZN(net3233)
);

INV_X32 c3090(
.A(net9557),
.ZN(net3234)
);

INV_X4 c3091(
.A(net3219),
.ZN(net3235)
);

OR3_X1 c3092(
.A1(net3195),
.A2(net3228),
.A3(net10979),
.ZN(net3236)
);

INV_X1 c3093(
.A(net2038),
.ZN(net3237)
);

NOR2_X1 c3094(
.A1(net2302),
.A2(net11121),
.ZN(net3238)
);

INV_X2 c3095(
.A(net10945),
.ZN(net3239)
);

INV_X8 c3096(
.A(net3165),
.ZN(net3240)
);

OR2_X2 c3097(
.A1(net2159),
.A2(net3217),
.ZN(net3241)
);

MUX2_X1 c3098(
.A(net3227),
.B(net3078),
.S(net2038),
.Z(net3242)
);

INV_X16 c3099(
.A(net10296),
.ZN(net3243)
);

NOR2_X4 c3100(
.A1(net3130),
.A2(net2203),
.ZN(net3244)
);

INV_X32 c3101(
.A(net3239),
.ZN(net3245)
);

OAI21_X4 c3102(
.A(net3226),
.B1(net2290),
.B2(net3144),
.ZN(net3246)
);

SDFFS_X1 c3103(
.D(net3237),
.SE(net2294),
.SI(net3144),
.SN(net11161),
.CK(clk),
.Q(net3248),
.QN(net3247)
);

INV_X4 c3104(
.A(net9730),
.ZN(net3249)
);

MUX2_X2 c3105(
.A(net3221),
.B(net2159),
.S(net2299),
.Z(net3250)
);

NAND3_X4 c3106(
.A1(net2884),
.A2(net2244),
.A3(net10999),
.ZN(net3251)
);

OR3_X4 c3107(
.A1(net1252),
.A2(net3238),
.A3(net3243),
.ZN(net3252)
);

AND3_X2 c3108(
.A1(net3252),
.A2(net2299),
.A3(net3239),
.ZN(net3253)
);

NOR2_X2 c3109(
.A1(net2313),
.A2(net10896),
.ZN(net3254)
);

INV_X1 c3110(
.A(net3123),
.ZN(net3255)
);

INV_X2 c3111(
.A(net9709),
.ZN(net3256)
);

DFFS_X1 c3112(
.D(net3197),
.SN(net3219),
.CK(clk),
.Q(net3258),
.QN(net3257)
);

INV_X8 c3113(
.A(net1995),
.ZN(net3259)
);

INV_X16 c3114(
.A(net3234),
.ZN(net3260)
);

XOR2_X2 c3115(
.A(net3256),
.B(net2245),
.Z(net3261)
);

XNOR2_X1 c3116(
.A(net3240),
.B(net3243),
.ZN(net3262)
);

DFFS_X2 c3117(
.D(net3250),
.SN(net3189),
.CK(clk),
.Q(net3264),
.QN(net3263)
);

INV_X32 c3118(
.A(net3231),
.ZN(net3265)
);

OR2_X4 c3119(
.A1(net3265),
.A2(net3259),
.ZN(net3266)
);

OR2_X1 c3120(
.A1(net3238),
.A2(net3266),
.ZN(net3267)
);

NOR3_X1 c3121(
.A1(net2307),
.A2(net1200),
.A3(net3231),
.ZN(net3268)
);

AOI22_X2 c3122(
.A1(net3267),
.A2(net3180),
.B1(net3218),
.B2(net3260),
.ZN(net3269)
);

XNOR2_X2 c3123(
.A(net3235),
.B(net1279),
.ZN(net3270)
);

CLKGATETST_X1 c3124(
.E(net3241),
.SE(net3269),
.CK(clk),
.GCK(net3271)
);

INV_X4 c3125(
.A(net2257),
.ZN(net3272)
);

OR3_X2 c3126(
.A1(net3236),
.A2(net2300),
.A3(net3265),
.ZN(net3273)
);

OAI21_X2 c3127(
.A(net1319),
.B1(net3239),
.B2(net3260),
.ZN(net3274)
);

INV_X1 c3128(
.A(net10853),
.ZN(net3275)
);

OAI21_X1 c3129(
.A(net3270),
.B1(net3153),
.B2(net3234),
.ZN(net3276)
);

DFFRS_X1 c3130(
.D(net3251),
.RN(net1230),
.SN(net2305),
.CK(clk),
.Q(net3278),
.QN(net3277)
);

AND2_X4 c3131(
.A1(net3217),
.A2(net3259),
.ZN(net3279)
);

AND2_X1 c3132(
.A1(net3230),
.A2(net3231),
.ZN(net3280)
);

AOI21_X2 c3133(
.A(net3242),
.B1(net3153),
.B2(net3271),
.ZN(net3281)
);

AOI21_X1 c3134(
.A(net3259),
.B1(net3275),
.B2(net3251),
.ZN(net3282)
);

NAND2_X1 c3135(
.A1(net3275),
.A2(net1252),
.ZN(net3283)
);

NAND2_X2 c3136(
.A1(net3253),
.A2(net3249),
.ZN(net3284)
);

NAND2_X4 c3137(
.A1(net2275),
.A2(net10896),
.ZN(net3285)
);

AOI21_X4 c3138(
.A(net3283),
.B1(net3279),
.B2(net2317),
.ZN(net3286)
);

DFFRS_X2 c3139(
.D(net3255),
.RN(net2248),
.SN(net3223),
.CK(clk),
.Q(net3288),
.QN(net3287)
);

AND2_X2 c3140(
.A1(net3268),
.A2(net3249),
.ZN(net3289)
);

XOR2_X1 c3141(
.A(net3272),
.B(net10955),
.Z(net3290)
);

NOR2_X1 c3142(
.A1(net3274),
.A2(net3123),
.ZN(net3291)
);

OR2_X2 c3143(
.A1(net3260),
.A2(net3280),
.ZN(net3292)
);

AND3_X1 c3144(
.A1(net3290),
.A2(net3287),
.A3(net3274),
.ZN(net3293)
);

NAND3_X1 c3145(
.A1(net3293),
.A2(net3263),
.A3(net3247),
.ZN(net3294)
);

NOR2_X4 c3146(
.A1(net3254),
.A2(net3180),
.ZN(net3295)
);

SDFF_X1 c3147(
.D(net3295),
.SE(net3294),
.SI(net3203),
.CK(clk),
.Q(net3297),
.QN(net3296)
);

NOR3_X4 c3148(
.A1(net3294),
.A2(net3271),
.A3(net3223),
.ZN(net3298)
);

NOR3_X2 c3149(
.A1(net3233),
.A2(net3218),
.A3(net3292),
.ZN(net3299)
);

AND3_X4 c3150(
.A1(net3288),
.A2(net3297),
.A3(net3254),
.ZN(net3300)
);

NOR2_X2 c3151(
.A1(net3280),
.A2(net3299),
.ZN(net3301)
);

OAI222_X1 c3152(
.A1(net3301),
.A2(net3281),
.B1(net3300),
.B2(net3260),
.C1(net3271),
.C2(net3292),
.ZN(net3302)
);

NAND4_X4 c3153(
.A1(net3299),
.A2(net3288),
.A3(net3283),
.A4(net3292),
.ZN(net3303)
);

INV_X2 c3154(
.A(net11134),
.ZN(net3304)
);

INV_X8 c3155(
.A(net2203),
.ZN(net3305)
);

XOR2_X2 c3156(
.A(net1208),
.B(net3081),
.Z(net3306)
);

INV_X16 c3157(
.A(net10931),
.ZN(net3307)
);

INV_X32 c3158(
.A(net10821),
.ZN(net3308)
);

XNOR2_X1 c3159(
.A(net337),
.B(net3271),
.ZN(net3309)
);

INV_X4 c3160(
.A(net10926),
.ZN(net3310)
);

NAND3_X2 c3161(
.A1(net2375),
.A2(net3283),
.A3(net3309),
.ZN(net3311)
);

INV_X1 c3162(
.A(net10234),
.ZN(net3312)
);

INV_X2 c3163(
.A(net3311),
.ZN(net3313)
);

OR2_X4 c3164(
.A1(net2355),
.A2(net2402),
.ZN(net3314)
);

OR2_X1 c3165(
.A1(net421),
.A2(net2314),
.ZN(net3315)
);

INV_X8 c3166(
.A(net2314),
.ZN(net3316)
);

XNOR2_X2 c3167(
.A(net2377),
.B(net3307),
.ZN(net3317)
);

AND2_X4 c3168(
.A1(net2407),
.A2(net3307),
.ZN(net3318)
);

AND2_X1 c3169(
.A1(net3314),
.A2(net1342),
.ZN(net3319)
);

INV_X16 c3170(
.A(net3317),
.ZN(net3320)
);

INV_X32 c3171(
.A(net3308),
.ZN(net3321)
);

OR3_X1 c3172(
.A1(net1444),
.A2(net3314),
.A3(net3129),
.ZN(net3322)
);

INV_X4 c3173(
.A(net9609),
.ZN(net3323)
);

INV_X1 c3174(
.A(net3245),
.ZN(net3324)
);

INV_X2 c3175(
.A(net3321),
.ZN(net3325)
);

INV_X8 c3176(
.A(net2405),
.ZN(net3326)
);

MUX2_X1 c3177(
.A(net3129),
.B(net2411),
.S(net2385),
.Z(net3327)
);

NAND2_X1 c3178(
.A1(net3289),
.A2(net3273),
.ZN(net3328)
);

INV_X16 c3179(
.A(net3309),
.ZN(net3329)
);

INV_X32 c3180(
.A(net2398),
.ZN(net3330)
);

INV_X4 c3181(
.A(net3320),
.ZN(net3331)
);

OAI21_X4 c3182(
.A(net2397),
.B1(net3285),
.B2(net2375),
.ZN(net3332)
);

INV_X1 c3183(
.A(net10107),
.ZN(net3333)
);

INV_X2 c3184(
.A(net11161),
.ZN(net3334)
);

NAND2_X2 c3185(
.A1(net3304),
.A2(net3273),
.ZN(net3335)
);

OAI222_X4 c3186(
.A1(net2312),
.A2(net3305),
.B1(net3296),
.B2(net3334),
.C1(net2317),
.C2(net2352),
.ZN(net3336)
);

MUX2_X2 c3187(
.A(net362),
.B(net2345),
.S(net10989),
.Z(net3337)
);

INV_X8 c3188(
.A(net9886),
.ZN(net3338)
);

INV_X16 c3189(
.A(net9958),
.ZN(net3339)
);

NAND2_X4 c3190(
.A1(net2284),
.A2(net3326),
.ZN(net3340)
);

AND2_X2 c3191(
.A1(net3331),
.A2(net3321),
.ZN(net3341)
);

XOR2_X1 c3192(
.A(net3328),
.B(net2398),
.Z(net3342)
);

INV_X32 c3193(
.A(net9709),
.ZN(net3343)
);

NOR2_X1 c3194(
.A1(net3326),
.A2(net2398),
.ZN(net3344)
);

INV_X4 c3195(
.A(net10977),
.ZN(net3345)
);

OR2_X2 c3196(
.A1(net3335),
.A2(net3334),
.ZN(net3346)
);

NOR2_X4 c3197(
.A1(net3345),
.A2(net3327),
.ZN(net3347)
);

NOR2_X2 c3198(
.A1(net3347),
.A2(net3335),
.ZN(net3348)
);

XOR2_X2 c3199(
.A(net3343),
.B(net2356),
.Z(net3349)
);

INV_X1 c3200(
.A(net3334),
.ZN(net3350)
);

XNOR2_X1 c3201(
.A(net3338),
.B(net421),
.ZN(net3351)
);

OR2_X4 c3202(
.A1(net3327),
.A2(net3334),
.ZN(net3352)
);

OR2_X1 c3203(
.A1(net3340),
.A2(net3333),
.ZN(net3353)
);

INV_X2 c3204(
.A(net10743),
.ZN(net3354)
);

OAI211_X2 c3205(
.A(net3352),
.B(net3310),
.C1(net2354),
.C2(net3348),
.ZN(net3355)
);

INV_X8 c3206(
.A(net10584),
.ZN(net3356)
);

INV_X16 c3207(
.A(net3337),
.ZN(net3357)
);

XNOR2_X2 c3208(
.A(net3339),
.B(net2404),
.ZN(net3358)
);

AND2_X4 c3209(
.A1(net3346),
.A2(net1334),
.ZN(net3359)
);

OR4_X2 c3210(
.A1(net3144),
.A2(net3352),
.A3(net3178),
.A4(net3260),
.ZN(net3360)
);

INV_X32 c3211(
.A(net3353),
.ZN(net3361)
);

AND2_X1 c3212(
.A1(net1382),
.A2(net3340),
.ZN(net3362)
);

INV_X4 c3213(
.A(net3349),
.ZN(net3363)
);

AOI221_X4 c3214(
.A(net3354),
.B1(net3359),
.B2(net3311),
.C1(net3297),
.C2(net3320),
.ZN(net3364)
);

INV_X1 c3215(
.A(net10976),
.ZN(net3365)
);

OAI222_X2 c3216(
.A1(net3363),
.A2(net3365),
.B1(net2398),
.B2(net1382),
.C1(net2209),
.C2(net3292),
.ZN(net3366)
);

NAND3_X4 c3217(
.A1(net2414),
.A2(net10551),
.A3(net10977),
.ZN(net3367)
);

NAND2_X1 c3218(
.A1(net421),
.A2(net10989),
.ZN(net3368)
);

INV_X2 c3219(
.A(net3332),
.ZN(net3369)
);

INV_X8 c3220(
.A(net10108),
.ZN(net3370)
);

INV_X16 c3221(
.A(net3273),
.ZN(net3371)
);

OR3_X4 c3222(
.A1(net3370),
.A2(net3328),
.A3(net3321),
.ZN(net3372)
);

NAND2_X2 c3223(
.A1(net3372),
.A2(net10875),
.ZN(net3373)
);

NAND2_X4 c3224(
.A1(net3357),
.A2(net11128),
.ZN(net3374)
);

INV_X32 c3225(
.A(net9609),
.ZN(net3375)
);

AND2_X2 c3226(
.A1(net3298),
.A2(net3337),
.ZN(net3376)
);

XOR2_X1 c3227(
.A(net3372),
.B(net3371),
.Z(net3377)
);

INV_X4 c3228(
.A(net3312),
.ZN(net3378)
);

NOR2_X1 c3229(
.A1(net3371),
.A2(net3129),
.ZN(net3379)
);

AND3_X2 c3230(
.A1(net3378),
.A2(net2356),
.A3(net337),
.ZN(net3380)
);

INV_X1 c3231(
.A(net10931),
.ZN(net3381)
);

NOR3_X1 c3232(
.A1(net2411),
.A2(net3380),
.A3(net3260),
.ZN(net3382)
);

INV_X2 c3233(
.A(net10938),
.ZN(net3383)
);

OR3_X2 c3234(
.A1(net3350),
.A2(net3383),
.A3(net3356),
.ZN(net3384)
);

OR2_X2 c3235(
.A1(net3381),
.A2(net3383),
.ZN(net3385)
);

NOR2_X4 c3236(
.A1(net3385),
.A2(net10999),
.ZN(net3386)
);

INV_X8 c3237(
.A(net3325),
.ZN(net3387)
);

INV_X16 c3238(
.A(net3125),
.ZN(net3388)
);

NOR2_X2 c3239(
.A1(net3271),
.A2(net2402),
.ZN(net3389)
);

XOR2_X2 c3240(
.A(net2479),
.B(net2455),
.Z(net3390)
);

XNOR2_X1 c3241(
.A(net1355),
.B(net3388),
.ZN(net3391)
);

INV_X32 c3242(
.A(net1494),
.ZN(net3392)
);

INV_X4 c3243(
.A(net1367),
.ZN(net3393)
);

OR2_X4 c3244(
.A1(net3389),
.A2(net1455),
.ZN(net3394)
);

INV_X1 c3245(
.A(net3387),
.ZN(net3395)
);

OR2_X1 c3246(
.A1(net3232),
.A2(net2345),
.ZN(net3396)
);

INV_X2 c3247(
.A(net10212),
.ZN(net3397)
);

OAI21_X2 c3248(
.A(net3313),
.B1(net2497),
.B2(net3291),
.ZN(net3398)
);

XNOR2_X2 c3249(
.A(net3297),
.B(net3356),
.ZN(net3399)
);

AND2_X4 c3250(
.A1(net3395),
.A2(net3216),
.ZN(net3400)
);

INV_X8 c3251(
.A(net2470),
.ZN(net3401)
);

SDFF_X2 c3252(
.D(net3326),
.SE(net3374),
.SI(net3305),
.CK(clk),
.Q(net3403),
.QN(net3402)
);

AND2_X1 c3253(
.A1(net2356),
.A2(net1471),
.ZN(net3404)
);

INV_X16 c3254(
.A(net2240),
.ZN(net3405)
);

INV_X32 c3255(
.A(net10814),
.ZN(net3406)
);

INV_X4 c3256(
.A(net9640),
.ZN(net3407)
);

INV_X1 c3257(
.A(net10955),
.ZN(net3408)
);

NAND2_X1 c3258(
.A1(net3323),
.A2(net11167),
.ZN(net3409)
);

NAND2_X2 c3259(
.A1(net3400),
.A2(net3399),
.ZN(net3410)
);

INV_X2 c3260(
.A(net10916),
.ZN(net3411)
);

INV_X8 c3261(
.A(net10442),
.ZN(net3412)
);

NAND2_X4 c3262(
.A1(net3412),
.A2(net3405),
.ZN(net3413)
);

INV_X16 c3263(
.A(net3389),
.ZN(net3414)
);

AND2_X2 c3264(
.A1(net3329),
.A2(net11166),
.ZN(net3415)
);

INV_X32 c3265(
.A(net3413),
.ZN(net3416)
);

XOR2_X1 c3266(
.A(net2509),
.B(net1507),
.Z(net3417)
);

NOR2_X1 c3267(
.A1(net2290),
.A2(net3379),
.ZN(net3418)
);

OR2_X2 c3268(
.A1(net3271),
.A2(net3405),
.ZN(net3419)
);

INV_X4 c3269(
.A(net2458),
.ZN(net3420)
);

NOR2_X4 c3270(
.A1(net3390),
.A2(net1392),
.ZN(net3421)
);

INV_X1 c3271(
.A(net10336),
.ZN(net3422)
);

NOR2_X2 c3272(
.A1(net3416),
.A2(net3415),
.ZN(net3423)
);

XOR2_X2 c3273(
.A(net3388),
.B(net2506),
.Z(net3424)
);

XNOR2_X1 c3274(
.A(net339),
.B(net3389),
.ZN(net3425)
);

OR2_X4 c3275(
.A1(net3276),
.A2(net3399),
.ZN(net3426)
);

OR2_X1 c3276(
.A1(net3407),
.A2(net2481),
.ZN(net3427)
);

XNOR2_X2 c3277(
.A(net3423),
.B(net2498),
.ZN(net3428)
);

INV_X2 c3278(
.A(net10002),
.ZN(net3429)
);

OAI21_X1 c3279(
.A(net3418),
.B1(net2454),
.B2(net3344),
.ZN(net3430)
);

AND2_X4 c3280(
.A1(net3392),
.A2(net10552),
.ZN(net3431)
);

INV_X8 c3281(
.A(net2402),
.ZN(net3432)
);

AOI21_X2 c3282(
.A(net3419),
.B1(net2239),
.B2(net3421),
.ZN(net3433)
);

AND2_X1 c3283(
.A1(net3432),
.A2(net2509),
.ZN(net3434)
);

INV_X16 c3284(
.A(net9639),
.ZN(net3435)
);

AOI21_X1 c3285(
.A(net3379),
.B1(net2470),
.B2(net3428),
.ZN(net3436)
);

AOI21_X4 c3286(
.A(net3426),
.B1(net3399),
.B2(net530),
.ZN(net3437)
);

AND3_X1 c3287(
.A1(net3436),
.A2(net1455),
.A3(net1367),
.ZN(net3438)
);

SDFFS_X2 c3288(
.D(net3437),
.SE(net3404),
.SI(net3369),
.SN(net3296),
.CK(clk),
.Q(net3440),
.QN(net3439)
);

NAND3_X1 c3289(
.A1(net530),
.A2(net3440),
.A3(net3428),
.ZN(net3441)
);

NAND2_X1 c3290(
.A1(net1455),
.A2(net3388),
.ZN(net3442)
);

NAND2_X2 c3291(
.A1(net2490),
.A2(net11048),
.ZN(net3443)
);

INV_X32 c3292(
.A(net10342),
.ZN(net3444)
);

INV_X4 c3293(
.A(net10192),
.ZN(net3445)
);

NOR3_X4 c3294(
.A1(net3434),
.A2(net3404),
.A3(net3411),
.ZN(net3446)
);

NAND2_X4 c3295(
.A1(net3401),
.A2(net1494),
.ZN(net3447)
);

INV_X1 c3296(
.A(net3431),
.ZN(net3448)
);

AND2_X2 c3297(
.A1(net3410),
.A2(net1484),
.ZN(net3449)
);

XOR2_X1 c3298(
.A(net2470),
.B(net10959),
.Z(net3450)
);

INV_X2 c3299(
.A(net10222),
.ZN(net3451)
);

NOR2_X1 c3300(
.A1(net3451),
.A2(net3449),
.ZN(net3452)
);

AOI211_X1 c3301(
.A(net1459),
.B(net3369),
.C1(net3405),
.C2(net3449),
.ZN(net3453)
);

OR2_X2 c3302(
.A1(net3435),
.A2(net3452),
.ZN(net3454)
);

DFFRS_X1 c3303(
.D(net3356),
.RN(net3438),
.SN(net3421),
.CK(clk),
.Q(net3456),
.QN(net3455)
);

NOR2_X4 c3304(
.A1(net3423),
.A2(net10757),
.ZN(net3457)
);

NOR3_X2 c3305(
.A1(net3440),
.A2(net3435),
.A3(net3216),
.ZN(net3458)
);

NOR2_X2 c3306(
.A1(net2345),
.A2(net3428),
.ZN(net3459)
);

INV_X8 c3307(
.A(net10998),
.ZN(net3460)
);

AOI222_X1 c3308(
.A1(net3438),
.A2(net3365),
.B1(net3459),
.B2(net3422),
.C1(net3324),
.C2(net2121),
.ZN(net3461)
);

AND3_X4 c3309(
.A1(net3424),
.A2(net3436),
.A3(net2433),
.ZN(net3462)
);

NAND3_X2 c3310(
.A1(net3452),
.A2(net3400),
.A3(net3460),
.ZN(net3463)
);

OR3_X1 c3311(
.A1(net3457),
.A2(net2345),
.A3(net11167),
.ZN(net3464)
);

XOR2_X2 c3312(
.A(net3414),
.B(net3439),
.Z(net3465)
);

NAND4_X2 c3313(
.A1(net3445),
.A2(net3324),
.A3(net3463),
.A4(net3460),
.ZN(net3466)
);

MUX2_X1 c3314(
.A(net3455),
.B(net3449),
.S(net10992),
.Z(net3467)
);

INV_X16 c3315(
.A(net9970),
.ZN(net3468)
);

OAI21_X4 c3316(
.A(net3468),
.B1(net3452),
.B2(net11170),
.ZN(net3469)
);

AOI222_X4 c3317(
.A1(net3464),
.A2(net3463),
.B1(net3467),
.B2(net1334),
.C1(net3369),
.C2(net3421),
.ZN(net3470)
);

MUX2_X2 c3318(
.A(net3422),
.B(net3415),
.S(net10551),
.Z(net3471)
);

NAND3_X4 c3319(
.A1(net2404),
.A2(net2402),
.A3(net3468),
.ZN(net3472)
);

INV_X32 c3320(
.A(net9541),
.ZN(net3473)
);

INV_X4 c3321(
.A(net2565),
.ZN(net3474)
);

XNOR2_X1 c3322(
.A(net2573),
.B(net2346),
.ZN(net3475)
);

INV_X1 c3323(
.A(net2497),
.ZN(net3476)
);

OR2_X4 c3324(
.A1(net2300),
.A2(net3467),
.ZN(net3477)
);

OR2_X1 c3325(
.A1(net2487),
.A2(net3324),
.ZN(net3478)
);

INV_X2 c3326(
.A(net2567),
.ZN(net3479)
);

INV_X8 c3327(
.A(net11030),
.ZN(net3480)
);

INV_X16 c3328(
.A(net618),
.ZN(net3481)
);

INV_X32 c3329(
.A(net9951),
.ZN(net3482)
);

XNOR2_X2 c3330(
.A(net2420),
.B(net2343),
.ZN(net3483)
);

INV_X4 c3331(
.A(net9897),
.ZN(net3484)
);

INV_X1 c3332(
.A(net2533),
.ZN(net3485)
);

INV_X2 c3333(
.A(net3483),
.ZN(net3486)
);

CLKGATETST_X2 c3334(
.E(net2566),
.SE(net3324),
.CK(clk),
.GCK(net3487)
);

AND2_X4 c3335(
.A1(net3420),
.A2(net2565),
.ZN(net3488)
);

INV_X8 c3336(
.A(net3474),
.ZN(net3489)
);

INV_X16 c3337(
.A(net3489),
.ZN(net3490)
);

AND2_X1 c3338(
.A1(net3488),
.A2(net3422),
.ZN(net3491)
);

NAND2_X1 c3339(
.A1(net2121),
.A2(net1587),
.ZN(net3492)
);

INV_X32 c3340(
.A(net9766),
.ZN(net3493)
);

OR3_X4 c3341(
.A1(net3473),
.A2(net3481),
.A3(net3478),
.ZN(net3494)
);

INV_X4 c3342(
.A(net3459),
.ZN(net3495)
);

NAND2_X2 c3343(
.A1(net3415),
.A2(net3460),
.ZN(net3496)
);

DFFRS_X2 c3344(
.D(net2574),
.RN(net2419),
.SN(net3291),
.CK(clk),
.Q(net3498),
.QN(net3497)
);

NAND2_X4 c3345(
.A1(net3487),
.A2(net3493),
.ZN(net3499)
);

INV_X1 c3346(
.A(net9766),
.ZN(net3500)
);

AND2_X2 c3347(
.A1(net3481),
.A2(net3423),
.ZN(net3501)
);

AND3_X2 c3348(
.A1(net2578),
.A2(net3481),
.A3(net2496),
.ZN(net3502)
);

XOR2_X1 c3349(
.A(net3400),
.B(net3487),
.Z(net3503)
);

INV_X2 c3350(
.A(net3496),
.ZN(net3504)
);

INV_X8 c3351(
.A(net9829),
.ZN(net3505)
);

NOR2_X1 c3352(
.A1(net2554),
.A2(net2573),
.ZN(net3506)
);

OR2_X2 c3353(
.A1(net1587),
.A2(net3504),
.ZN(net3507)
);

INV_X16 c3354(
.A(net9996),
.ZN(net3508)
);

INV_X32 c3355(
.A(net2550),
.ZN(net3509)
);

INV_X4 c3356(
.A(net3506),
.ZN(net3510)
);

INV_X1 c3357(
.A(net10155),
.ZN(net3511)
);

NOR2_X4 c3358(
.A1(net3509),
.A2(net3423),
.ZN(net3512)
);

NOR2_X2 c3359(
.A1(net3500),
.A2(net3511),
.ZN(net3513)
);

INV_X2 c3360(
.A(net3456),
.ZN(net3514)
);

XOR2_X2 c3361(
.A(net1384),
.B(net3486),
.Z(net3515)
);

XNOR2_X1 c3362(
.A(net2561),
.B(net3511),
.ZN(net3516)
);

OR2_X4 c3363(
.A1(net3504),
.A2(net3386),
.ZN(net3517)
);

OR2_X1 c3364(
.A1(net3502),
.A2(net3514),
.ZN(net3518)
);

XNOR2_X2 c3365(
.A(net3476),
.B(net3507),
.ZN(net3519)
);

AND2_X4 c3366(
.A1(net3510),
.A2(net3478),
.ZN(net3520)
);

INV_X8 c3367(
.A(net3511),
.ZN(net3521)
);

AND2_X1 c3368(
.A1(net3484),
.A2(net2521),
.ZN(net3522)
);

OAI33_X1 c3369(
.A1(net3382),
.A2(net3514),
.A3(net2593),
.B1(net3404),
.B2(net2521),
.B3(net1493),
.ZN(net3523)
);

INV_X16 c3370(
.A(net11108),
.ZN(net3524)
);

NOR3_X1 c3371(
.A1(net3487),
.A2(net1617),
.A3(net3511),
.ZN(net3525)
);

INV_X32 c3372(
.A(net11101),
.ZN(net3526)
);

NAND2_X1 c3373(
.A1(net3520),
.A2(net3511),
.ZN(net3527)
);

INV_X4 c3374(
.A(net10017),
.ZN(net3528)
);

INV_X1 c3375(
.A(net3503),
.ZN(net3529)
);

INV_X2 c3376(
.A(net3512),
.ZN(net3530)
);

AOI221_X2 c3377(
.A(net1484),
.B1(net3514),
.B2(net3524),
.C1(net2553),
.C2(net2593),
.ZN(net3531)
);

OR3_X2 c3378(
.A1(net3478),
.A2(net3530),
.A3(net2884),
.ZN(net3532)
);

OAI21_X2 c3379(
.A(net2423),
.B1(net3403),
.B2(net3530),
.ZN(net3533)
);

NAND2_X2 c3380(
.A1(net3528),
.A2(net3511),
.ZN(net3534)
);

NAND2_X4 c3381(
.A1(net3508),
.A2(net3514),
.ZN(net3535)
);

OAI21_X1 c3382(
.A(net3423),
.B1(net3518),
.B2(net3514),
.ZN(net3536)
);

INV_X8 c3383(
.A(net10992),
.ZN(net3537)
);

AND2_X2 c3384(
.A1(net3393),
.A2(net2565),
.ZN(net3538)
);

XOR2_X1 c3385(
.A(net3531),
.B(net3530),
.Z(net3539)
);

NOR2_X1 c3386(
.A1(net3514),
.A2(net3528),
.ZN(net3540)
);

AOI21_X2 c3387(
.A(net3524),
.B1(net3494),
.B2(net2496),
.ZN(net3541)
);

OR2_X2 c3388(
.A1(net3537),
.A2(net3474),
.ZN(net3542)
);

AOI21_X1 c3389(
.A(net3526),
.B1(net3495),
.B2(net3504),
.ZN(net3543)
);

INV_X16 c3390(
.A(net9541),
.ZN(net3544)
);

NOR2_X4 c3391(
.A1(net3534),
.A2(net3544),
.ZN(net3545)
);

NOR2_X2 c3392(
.A1(net3507),
.A2(net3534),
.ZN(net3546)
);

AOI21_X4 c3393(
.A(net3516),
.B1(net3545),
.B2(net3546),
.ZN(net3547)
);

XOR2_X2 c3394(
.A(net3539),
.B(net3546),
.Z(net3548)
);

AND3_X1 c3395(
.A1(net3529),
.A2(net3530),
.A3(net3544),
.ZN(net3549)
);

SDFF_X1 c3396(
.D(net3530),
.SE(net3527),
.SI(net3549),
.CK(clk),
.Q(net3551),
.QN(net3550)
);

XNOR2_X1 c3397(
.A(net3541),
.B(net10378),
.ZN(net3552)
);

NAND3_X1 c3398(
.A1(net2596),
.A2(net1291),
.A3(net3550),
.ZN(net3553)
);

NOR3_X4 c3399(
.A1(net3553),
.A2(net3545),
.A3(net3530),
.ZN(net3554)
);

NOR3_X2 c3400(
.A1(net2494),
.A2(net3540),
.A3(net3554),
.ZN(net3555)
);

OR2_X4 c3401(
.A1(net3551),
.A2(net10378),
.ZN(net3556)
);

AND3_X4 c3402(
.A1(net3556),
.A2(net3544),
.A3(net10671),
.ZN(net3557)
);

OR2_X1 c3403(
.A1(net2612),
.A2(net684),
.ZN(net3558)
);

XNOR2_X2 c3404(
.A(net3480),
.B(net3525),
.ZN(net3559)
);

AND2_X4 c3405(
.A1(net1334),
.A2(net2585),
.ZN(net3560)
);

AND2_X1 c3406(
.A1(net1589),
.A2(net2553),
.ZN(net3561)
);

NAND2_X1 c3407(
.A1(net499),
.A2(net3518),
.ZN(net3562)
);

INV_X32 c3408(
.A(net10870),
.ZN(net3563)
);

INV_X4 c3409(
.A(net10730),
.ZN(net3564)
);

INV_X1 c3410(
.A(net3485),
.ZN(net3565)
);

INV_X2 c3411(
.A(net3443),
.ZN(net3566)
);

CLKGATETST_X4 c3412(
.E(net3449),
.SE(net2569),
.CK(clk),
.GCK(net3567)
);

INV_X8 c3413(
.A(net10870),
.ZN(net3568)
);

INV_X16 c3414(
.A(net3547),
.ZN(net3569)
);

NAND2_X2 c3415(
.A1(net3490),
.A2(net2612),
.ZN(net3570)
);

NAND2_X4 c3416(
.A1(net3549),
.A2(net3494),
.ZN(net3571)
);

INV_X32 c3417(
.A(net3392),
.ZN(net3572)
);

NAND3_X2 c3418(
.A1(net3305),
.A2(net3515),
.A3(net2612),
.ZN(net3573)
);

INV_X4 c3419(
.A(net10169),
.ZN(net3574)
);

AND2_X2 c3420(
.A1(net3501),
.A2(net3542),
.ZN(net3575)
);

INV_X1 c3421(
.A(net11039),
.ZN(net3576)
);

INV_X2 c3422(
.A(net3486),
.ZN(net3577)
);

XOR2_X1 c3423(
.A(net3567),
.B(net3486),
.Z(net3578)
);

SDFF_X2 c3424(
.D(net1505),
.SE(net3449),
.SI(net645),
.CK(clk),
.Q(net3580),
.QN(net3579)
);

NOR2_X1 c3425(
.A1(net3444),
.A2(net3579),
.ZN(net3581)
);

OR2_X2 c3426(
.A1(net2447),
.A2(net2674),
.ZN(net3582)
);

NOR2_X4 c3427(
.A1(net746),
.A2(net2553),
.ZN(net3583)
);

NOR2_X2 c3428(
.A1(net3542),
.A2(net3549),
.ZN(net3584)
);

XOR2_X2 c3429(
.A(net1625),
.B(net3449),
.Z(net3585)
);

XNOR2_X1 c3430(
.A(net2585),
.B(net3575),
.ZN(net3586)
);

INV_X8 c3431(
.A(net10870),
.ZN(net3587)
);

OR3_X1 c3432(
.A1(net3573),
.A2(net3583),
.A3(net1707),
.ZN(net3588)
);

OR2_X4 c3433(
.A1(net3482),
.A2(net2521),
.ZN(net3589)
);

OR2_X1 c3434(
.A1(net2303),
.A2(net3580),
.ZN(net3590)
);

INV_X16 c3435(
.A(net10994),
.ZN(net3591)
);

INV_X32 c3436(
.A(net10884),
.ZN(net3592)
);

XNOR2_X2 c3437(
.A(net3585),
.B(net2585),
.ZN(net3593)
);

INV_X4 c3438(
.A(net3572),
.ZN(net3594)
);

AND2_X4 c3439(
.A1(net1502),
.A2(net3576),
.ZN(net3595)
);

INV_X1 c3440(
.A(net10238),
.ZN(net3596)
);

AND2_X1 c3441(
.A1(net3564),
.A2(net2612),
.ZN(net3597)
);

INV_X2 c3442(
.A(net10771),
.ZN(net3598)
);

NAND2_X1 c3443(
.A1(net3577),
.A2(net2624),
.ZN(net3599)
);

NAND2_X2 c3444(
.A1(net3581),
.A2(net3586),
.ZN(net3600)
);

INV_X8 c3445(
.A(net9803),
.ZN(net3601)
);

NAND2_X4 c3446(
.A1(net2639),
.A2(net3582),
.ZN(net3602)
);

INV_X16 c3447(
.A(net10963),
.ZN(net3603)
);

MUX2_X1 c3448(
.A(net3596),
.B(net2121),
.S(net3587),
.Z(net3604)
);

AND2_X2 c3449(
.A1(net3574),
.A2(net3593),
.ZN(net3605)
);

XOR2_X1 c3450(
.A(net3563),
.B(net3494),
.Z(net3606)
);

NOR2_X1 c3451(
.A1(net3594),
.A2(net10902),
.ZN(net3607)
);

INV_X32 c3452(
.A(net11120),
.ZN(net3608)
);

OR2_X2 c3453(
.A1(net3599),
.A2(net10902),
.ZN(net3609)
);

NOR2_X4 c3454(
.A1(net3525),
.A2(net3560),
.ZN(net3610)
);

NOR2_X2 c3455(
.A1(net3587),
.A2(net3607),
.ZN(net3611)
);

XOR2_X2 c3456(
.A(net3518),
.B(net2597),
.Z(net3612)
);

XNOR2_X1 c3457(
.A(net2334),
.B(net3562),
.ZN(net3613)
);

OR2_X4 c3458(
.A1(net3579),
.A2(net10858),
.ZN(net3614)
);

OAI21_X4 c3459(
.A(net3499),
.B1(net3614),
.B2(net3587),
.ZN(net3615)
);

OR2_X1 c3460(
.A1(net3604),
.A2(net3486),
.ZN(net3616)
);

XNOR2_X2 c3461(
.A(net3607),
.B(net3578),
.ZN(net3617)
);

AND2_X4 c3462(
.A1(net3608),
.A2(net3578),
.ZN(net3618)
);

AND2_X1 c3463(
.A1(net3559),
.A2(net3618),
.ZN(net3619)
);

NAND2_X1 c3464(
.A1(net3523),
.A2(net3619),
.ZN(net3620)
);

MUX2_X2 c3465(
.A(net3606),
.B(net2665),
.S(net3615),
.Z(net3621)
);

AOI222_X2 c3466(
.A1(net3590),
.A2(net3475),
.B1(net3562),
.B2(net3615),
.C1(net2612),
.C2(net3565),
.ZN(net3622)
);

AOI221_X1 c3467(
.A(net3621),
.B1(net1681),
.B2(net3583),
.C1(net3581),
.C2(net3615),
.ZN(net3623)
);

NAND2_X2 c3468(
.A1(net3592),
.A2(net1667),
.ZN(net3624)
);

INV_X4 c3469(
.A(net10884),
.ZN(net3625)
);

INV_X1 c3470(
.A(net10817),
.ZN(net3626)
);

NAND3_X4 c3471(
.A1(net3323),
.A2(net3617),
.A3(net3567),
.ZN(net3627)
);

INV_X2 c3472(
.A(net9882),
.ZN(net3628)
);

NAND2_X4 c3473(
.A1(net3628),
.A2(net682),
.ZN(net3629)
);

AND2_X2 c3474(
.A1(net3629),
.A2(net10882),
.ZN(net3630)
);

XOR2_X1 c3475(
.A(net3546),
.B(net3565),
.Z(net3631)
);

NOR2_X1 c3476(
.A1(net3607),
.A2(net10882),
.ZN(net3632)
);

OR2_X2 c3477(
.A1(net2620),
.A2(net3632),
.ZN(net3633)
);

OR3_X4 c3478(
.A1(net3633),
.A2(net3581),
.A3(net3619),
.ZN(net3634)
);

AND3_X2 c3479(
.A1(net3633),
.A2(net3567),
.A3(net10858),
.ZN(net3635)
);

OAI221_X1 c3480(
.A(net3632),
.B1(net3547),
.B2(net3615),
.C1(net3565),
.C2(net1579),
.ZN(net3636)
);

NOR2_X4 c3481(
.A1(net3631),
.A2(net3560),
.ZN(net3637)
);

NOR2_X2 c3482(
.A1(net3627),
.A2(net3631),
.ZN(net3638)
);

XOR2_X2 c3483(
.A(net2478),
.B(net3627),
.Z(net3639)
);

SDFFRS_X1 c3484(
.D(net3638),
.RN(net3627),
.SE(net3633),
.SI(net3402),
.SN(net3615),
.CK(clk),
.Q(net3641),
.QN(net3640)
);

OR4_X4 c3485(
.A1(net2626),
.A2(net3633),
.A3(net3641),
.A4(net3615),
.ZN(net3642)
);

INV_X8 c3486(
.A(net831),
.ZN(net3643)
);

INV_X16 c3487(
.A(net10912),
.ZN(net3644)
);

XNOR2_X1 c3488(
.A(net2728),
.B(net2710),
.ZN(net3645)
);

INV_X32 c3489(
.A(net11173),
.ZN(net3646)
);

OR2_X4 c3490(
.A1(net2705),
.A2(net2766),
.ZN(net3647)
);

OR2_X1 c3491(
.A1(net489),
.A2(net2741),
.ZN(net3648)
);

INV_X4 c3492(
.A(net9542),
.ZN(net3649)
);

XNOR2_X2 c3493(
.A(net3582),
.B(net2765),
.ZN(net3650)
);

AND2_X4 c3494(
.A1(net1759),
.A2(net762),
.ZN(net3651)
);

INV_X1 c3495(
.A(net11009),
.ZN(net3652)
);

NOR3_X1 c3496(
.A1(net1655),
.A2(net3624),
.A3(net3615),
.ZN(net3653)
);

AND2_X1 c3497(
.A1(net2693),
.A2(net3653),
.ZN(net3654)
);

INV_X2 c3498(
.A(net10409),
.ZN(net3655)
);

NAND2_X1 c3499(
.A1(net2711),
.A2(net3492),
.ZN(net3656)
);

INV_X8 c3500(
.A(net1671),
.ZN(net3657)
);

OAI22_X2 c3501(
.A1(net777),
.A2(net2677),
.B1(net3653),
.B2(net10793),
.ZN(net3658)
);

INV_X16 c3502(
.A(net2755),
.ZN(net3659)
);

OR3_X2 c3503(
.A1(net2761),
.A2(net3657),
.A3(net2715),
.ZN(net3660)
);

INV_X32 c3504(
.A(net9543),
.ZN(net3661)
);

OAI21_X2 c3505(
.A(net460),
.B1(net3491),
.B2(net2715),
.ZN(net3662)
);

DFFRS_X1 c3506(
.D(net3591),
.RN(net2761),
.SN(net3657),
.CK(clk),
.Q(net3664),
.QN(net3663)
);

NAND2_X2 c3507(
.A1(net3652),
.A2(net3578),
.ZN(net3665)
);

OAI211_X4 c3508(
.A(net3643),
.B(net2686),
.C1(net3663),
.C2(net3615),
.ZN(net3666)
);

OAI21_X1 c3509(
.A(net2714),
.B1(net3644),
.B2(net10395),
.ZN(net3667)
);

NAND2_X4 c3510(
.A1(net3324),
.A2(net1720),
.ZN(net3668)
);

AND2_X2 c3511(
.A1(net3580),
.A2(net828),
.ZN(net3669)
);

INV_X4 c3512(
.A(net11044),
.ZN(net3670)
);

AOI21_X2 c3513(
.A(net1759),
.B1(net3661),
.B2(net10959),
.ZN(net3671)
);

INV_X1 c3514(
.A(net10356),
.ZN(net3672)
);

XOR2_X1 c3515(
.A(net2765),
.B(net2725),
.Z(net3673)
);

INV_X2 c3516(
.A(net10295),
.ZN(net3674)
);

NOR2_X1 c3517(
.A1(net2670),
.A2(net3657),
.ZN(net3675)
);

OR2_X2 c3518(
.A1(net3655),
.A2(net827),
.ZN(net3676)
);

NOR2_X4 c3519(
.A1(net1666),
.A2(net3674),
.ZN(net3677)
);

NOR2_X2 c3520(
.A1(net3661),
.A2(net3674),
.ZN(net3678)
);

XOR2_X2 c3521(
.A(net3669),
.B(net1768),
.Z(net3679)
);

INV_X8 c3522(
.A(net3671),
.ZN(net3680)
);

XNOR2_X1 c3523(
.A(net3680),
.B(net3672),
.ZN(net3681)
);

OR2_X4 c3524(
.A1(net3515),
.A2(net3653),
.ZN(net3682)
);

OR2_X1 c3525(
.A1(net2647),
.A2(net3680),
.ZN(net3683)
);

AOI21_X1 c3526(
.A(net1753),
.B1(net2728),
.B2(net10972),
.ZN(net3684)
);

XNOR2_X2 c3527(
.A(net2725),
.B(net2677),
.ZN(net3685)
);

AND2_X4 c3528(
.A1(net2708),
.A2(net3676),
.ZN(net3686)
);

AOI21_X4 c3529(
.A(net3681),
.B1(net3670),
.B2(net3667),
.ZN(net3687)
);

INV_X16 c3530(
.A(net10808),
.ZN(net3688)
);

AND2_X1 c3531(
.A1(net3645),
.A2(net2677),
.ZN(net3689)
);

AND3_X1 c3532(
.A1(net2694),
.A2(net3681),
.A3(net3657),
.ZN(net3690)
);

NAND2_X1 c3533(
.A1(net3687),
.A2(net3646),
.ZN(net3691)
);

NAND2_X2 c3534(
.A1(net3674),
.A2(net11172),
.ZN(net3692)
);

NAND2_X4 c3535(
.A1(net823),
.A2(net2759),
.ZN(net3693)
);

AND2_X2 c3536(
.A1(net3679),
.A2(net3565),
.ZN(net3694)
);

INV_X32 c3537(
.A(net11034),
.ZN(net3695)
);

XOR2_X1 c3538(
.A(net3654),
.B(net3681),
.Z(net3696)
);

INV_X4 c3539(
.A(net10323),
.ZN(net3697)
);

CLKGATETST_X8 c3540(
.E(net3658),
.SE(net3681),
.CK(clk),
.GCK(net3698)
);

NOR2_X1 c3541(
.A1(net3693),
.A2(net2425),
.ZN(net3699)
);

OR2_X2 c3542(
.A1(net3665),
.A2(net3676),
.ZN(net3700)
);

NOR2_X4 c3543(
.A1(net3675),
.A2(net1655),
.ZN(net3701)
);

NAND3_X1 c3544(
.A1(net3683),
.A2(net3684),
.A3(net2569),
.ZN(net3702)
);

OAI222_X1 c3545(
.A1(net3692),
.A2(net3683),
.B1(net682),
.B2(net2670),
.C1(net3682),
.C2(net3672),
.ZN(net3703)
);

NOR2_X2 c3546(
.A1(net3701),
.A2(net3699),
.ZN(net3704)
);

DFFR_X1 c3547(
.D(net3668),
.RN(net2569),
.CK(clk),
.Q(net3706),
.QN(net3705)
);

XOR2_X2 c3548(
.A(net3662),
.B(net3661),
.Z(net3707)
);

NOR3_X4 c3549(
.A1(net3697),
.A2(net3705),
.A3(net3684),
.ZN(net3708)
);

XNOR2_X1 c3550(
.A(net3704),
.B(net2425),
.ZN(net3709)
);

OAI222_X4 c3551(
.A1(net3666),
.A2(net3704),
.B1(net3681),
.B2(net3691),
.C1(net3698),
.C2(net11173),
.ZN(net3710)
);

OR2_X4 c3552(
.A1(net3682),
.A2(net3666),
.ZN(net3711)
);

NOR3_X2 c3553(
.A1(net734),
.A2(net2499),
.A3(net3694),
.ZN(net3712)
);

INV_X1 c3554(
.A(net3657),
.ZN(net3713)
);

OAI221_X4 c3555(
.A(net2681),
.B1(net3707),
.B2(net3687),
.C1(net3672),
.C2(net1720),
.ZN(net3714)
);

DFFRS_X2 c3556(
.D(net3711),
.RN(net3658),
.SN(net3447),
.CK(clk),
.Q(net3716),
.QN(net3715)
);

OR2_X1 c3557(
.A1(net3578),
.A2(net3674),
.ZN(net3717)
);

AND3_X4 c3558(
.A1(net3706),
.A2(net3671),
.A3(net10654),
.ZN(net3718)
);

OAI211_X1 c3559(
.A(net3709),
.B(net3682),
.C1(net3673),
.C2(net3715),
.ZN(net3719)
);

OAI221_X2 c3560(
.A(net2731),
.B1(net3698),
.B2(net2715),
.C1(net3672),
.C2(net11037),
.ZN(net3720)
);

NAND3_X2 c3561(
.A1(net3717),
.A2(net1709),
.A3(net2677),
.ZN(net3721)
);

INV_X2 c3562(
.A(net10210),
.ZN(net3722)
);

AOI221_X4 c3563(
.A(net3649),
.B1(net3680),
.B2(net3722),
.C1(net3672),
.C2(net1666),
.ZN(net3723)
);

OR3_X1 c3564(
.A1(net1623),
.A2(net3716),
.A3(net1783),
.ZN(net3724)
);

MUX2_X1 c3565(
.A(net3720),
.B(net3722),
.S(net11025),
.Z(net3725)
);

SDFFR_X1 c3566(
.D(net3684),
.RN(net2472),
.SE(net2685),
.SI(net3663),
.CK(clk),
.Q(net3727),
.QN(net3726)
);

NOR4_X4 c3567(
.A1(net3725),
.A2(net3726),
.A3(net3653),
.A4(net11025),
.ZN(net3728)
);

AOI221_X2 c3568(
.A(net3673),
.B1(net3727),
.B2(net2759),
.C1(net3722),
.C2(net10858),
.ZN(net3729)
);

NOR4_X2 c3569(
.A1(net3492),
.A2(net1868),
.A3(net3615),
.A4(net1833),
.ZN(net3730)
);

XNOR2_X2 c3570(
.A(net895),
.B(net3618),
.ZN(net3731)
);

AND2_X4 c3571(
.A1(net1869),
.A2(net762),
.ZN(net3732)
);

AND2_X1 c3572(
.A1(net1850),
.A2(net2848),
.ZN(net3733)
);

NAND2_X1 c3573(
.A1(net2813),
.A2(net2809),
.ZN(net3734)
);

INV_X8 c3574(
.A(net9552),
.ZN(net3735)
);

NAND2_X2 c3575(
.A1(net2848),
.A2(net1779),
.ZN(net3736)
);

INV_X16 c3576(
.A(net9688),
.ZN(net3737)
);

OAI21_X4 c3577(
.A(net865),
.B1(net2733),
.B2(net1846),
.ZN(net3738)
);

DFFR_X2 c3578(
.D(net2769),
.RN(net3653),
.CK(clk),
.Q(net3740),
.QN(net3739)
);

NAND2_X4 c3579(
.A1(net1801),
.A2(net2814),
.ZN(net3741)
);

AND2_X2 c3580(
.A1(net2771),
.A2(net3664),
.ZN(net3742)
);

XOR2_X1 c3581(
.A(net905),
.B(net11120),
.Z(net3743)
);

MUX2_X2 c3582(
.A(net3664),
.B(net3742),
.S(net3739),
.Z(net3744)
);

NOR2_X1 c3583(
.A1(net2767),
.A2(net10856),
.ZN(net3745)
);

OR2_X2 c3584(
.A1(net3745),
.A2(net3641),
.ZN(net3746)
);

NOR2_X4 c3585(
.A1(net2831),
.A2(net2714),
.ZN(net3747)
);

NOR2_X2 c3586(
.A1(net1805),
.A2(net1779),
.ZN(net3748)
);

SDFF_X1 c3587(
.D(net902),
.SE(net2710),
.SI(net2809),
.CK(clk),
.Q(net3750),
.QN(net3749)
);

XOR2_X2 c3588(
.A(net3732),
.B(net1846),
.Z(net3751)
);

NAND3_X4 c3589(
.A1(net2800),
.A2(net1779),
.A3(net2821),
.ZN(net3752)
);

XNOR2_X1 c3590(
.A(net1615),
.B(net10678),
.ZN(net3753)
);

INV_X32 c3591(
.A(net10170),
.ZN(net3754)
);

DFFS_X1 c3592(
.D(net2853),
.SN(net3746),
.CK(clk),
.Q(net3756),
.QN(net3755)
);

OR2_X4 c3593(
.A1(net2836),
.A2(net3647),
.ZN(net3757)
);

OR3_X4 c3594(
.A1(net3730),
.A2(net2820),
.A3(net1869),
.ZN(net3758)
);

OR2_X1 c3595(
.A1(net3648),
.A2(net2680),
.ZN(net3759)
);

XNOR2_X2 c3596(
.A(net1862),
.B(net3747),
.ZN(net3760)
);

AND2_X4 c3597(
.A1(net3735),
.A2(net10606),
.ZN(net3761)
);

AND2_X1 c3598(
.A1(net2796),
.A2(net1827),
.ZN(net3762)
);

AND3_X2 c3599(
.A1(net3760),
.A2(net3730),
.A3(net865),
.ZN(net3763)
);

NOR3_X1 c3600(
.A1(net3761),
.A2(net3760),
.A3(net2808),
.ZN(net3764)
);

NAND2_X1 c3601(
.A1(net2793),
.A2(net2821),
.ZN(net3765)
);

NAND2_X2 c3602(
.A1(net2741),
.A2(net1857),
.ZN(net3766)
);

OR3_X2 c3603(
.A1(net1834),
.A2(net2715),
.A3(net10510),
.ZN(net3767)
);

NAND2_X4 c3604(
.A1(net3566),
.A2(net2557),
.ZN(net3768)
);

INV_X4 c3605(
.A(net10247),
.ZN(net3769)
);

AND2_X2 c3606(
.A1(net2714),
.A2(net3736),
.ZN(net3770)
);

XOR2_X1 c3607(
.A(net2715),
.B(net867),
.Z(net3771)
);

SDFF_X2 c3608(
.D(net3763),
.SE(net3733),
.SI(net3492),
.CK(clk),
.Q(net3773),
.QN(net3772)
);

NOR2_X1 c3609(
.A1(net3735),
.A2(net3751),
.ZN(net3774)
);

OAI21_X2 c3610(
.A(net3754),
.B1(net3760),
.B2(net877),
.ZN(net3775)
);

DFFRS_X1 c3611(
.D(net3740),
.RN(net2769),
.SN(net2710),
.CK(clk),
.Q(net3777),
.QN(net3776)
);

OR2_X2 c3612(
.A1(net3759),
.A2(net10856),
.ZN(net3778)
);

OAI21_X1 c3613(
.A(net3644),
.B1(net3760),
.B2(net3768),
.ZN(net3779)
);

AOI21_X2 c3614(
.A(net3770),
.B1(net3772),
.B2(net2799),
.ZN(net3780)
);

NOR2_X4 c3615(
.A1(net2840),
.A2(net11120),
.ZN(net3781)
);

INV_X1 c3616(
.A(net10138),
.ZN(net3782)
);

NOR2_X2 c3617(
.A1(net3688),
.A2(net2820),
.ZN(net3783)
);

AOI21_X1 c3618(
.A(net2799),
.B1(net2779),
.B2(net3760),
.ZN(net3784)
);

AOI21_X4 c3619(
.A(net2793),
.B1(net3755),
.B2(net10695),
.ZN(net3785)
);

XOR2_X2 c3620(
.A(net1846),
.B(net2789),
.Z(net3786)
);

XNOR2_X1 c3621(
.A(net877),
.B(net3716),
.ZN(net3787)
);

OR2_X4 c3622(
.A1(net2780),
.A2(net3782),
.ZN(net3788)
);

OR2_X1 c3623(
.A1(net3753),
.A2(net3783),
.ZN(net3789)
);

AND3_X1 c3624(
.A1(net1841),
.A2(net3751),
.A3(net3749),
.ZN(net3790)
);

DFFS_X2 c3625(
.D(net3790),
.SN(net1827),
.CK(clk),
.Q(net3792),
.QN(net3791)
);

XNOR2_X2 c3626(
.A(net3653),
.B(net3782),
.ZN(net3793)
);

NAND3_X1 c3627(
.A1(net2710),
.A2(net3785),
.A3(net3782),
.ZN(net3794)
);

AND2_X4 c3628(
.A1(net1708),
.A2(net3793),
.ZN(net3795)
);

AND2_X1 c3629(
.A1(net1681),
.A2(net2813),
.ZN(net3796)
);

AOI211_X4 c3630(
.A(net3765),
.B(net3788),
.C1(net3777),
.C2(net3492),
.ZN(net3797)
);

CLKGATETST_X1 c3631(
.E(net3779),
.SE(net3789),
.CK(clk),
.GCK(net3798)
);

NAND2_X1 c3632(
.A1(net762),
.A2(net2857),
.ZN(net3799)
);

OAI222_X2 c3633(
.A1(net1853),
.A2(net3799),
.B1(net3776),
.B2(net851),
.C1(net2808),
.C2(net2851),
.ZN(net3800)
);

SDFFR_X2 c3634(
.D(net3793),
.RN(net3783),
.SE(net3790),
.SI(net3653),
.CK(clk),
.Q(net3802),
.QN(net3801)
);

NOR4_X1 c3635(
.A1(net3775),
.A2(net3566),
.A3(net2680),
.A4(net3797),
.ZN(net3803)
);

SDFFS_X1 c3636(
.D(net3748),
.SE(net3801),
.SI(net3789),
.SN(net1801),
.CK(clk),
.Q(net3805),
.QN(net3804)
);

AOI211_X2 c3637(
.A(net2827),
.B(net3771),
.C1(net2804),
.C2(net1861),
.ZN(net3806)
);

NAND2_X2 c3638(
.A1(net3799),
.A2(net10731),
.ZN(net3807)
);

NOR3_X4 c3639(
.A1(net3743),
.A2(net3767),
.A3(net3783),
.ZN(net3808)
);

SDFFS_X2 c3640(
.D(net3793),
.SE(net3797),
.SI(net2809),
.SN(net10674),
.CK(clk),
.Q(net3810),
.QN(net3809)
);

INV_X2 c3641(
.A(net9551),
.ZN(net3811)
);

NOR3_X2 c3642(
.A1(net3731),
.A2(net2838),
.A3(net3759),
.ZN(net3812)
);

SDFFR_X1 c3643(
.D(net3795),
.RN(net3805),
.SE(net2821),
.SI(net3776),
.CK(clk),
.Q(net3814),
.QN(net3813)
);

AOI22_X1 c3644(
.A1(net2770),
.A2(net3786),
.B1(net3782),
.B2(net10673),
.ZN(net3815)
);

AND3_X4 c3645(
.A1(net3647),
.A2(net3796),
.A3(net3768),
.ZN(net3816)
);

SDFFR_X2 c3646(
.D(net3767),
.RN(net3787),
.SE(net3813),
.SI(net1846),
.CK(clk),
.Q(net3818),
.QN(net3817)
);

AND4_X4 c3647(
.A1(net3751),
.A2(net3810),
.A3(net3804),
.A4(net3619),
.ZN(net3819)
);

DFFRS_X2 c3648(
.D(net2817),
.RN(net3756),
.SN(net2831),
.CK(clk),
.Q(net3821),
.QN(net3820)
);

SDFF_X1 c3649(
.D(net3815),
.SE(net3819),
.SI(net3809),
.CK(clk),
.Q(net3823),
.QN(net3822)
);

NAND4_X1 c3650(
.A1(net3799),
.A2(net3814),
.A3(net3819),
.A4(net3782),
.ZN(net3824)
);

NAND3_X2 c3651(
.A1(net887),
.A2(net708),
.A3(net10766),
.ZN(net3825)
);

INV_X8 c3652(
.A(net9649),
.ZN(net3826)
);

INV_X16 c3653(
.A(net988),
.ZN(net3827)
);

INV_X32 c3654(
.A(net9649),
.ZN(net3828)
);

INV_X4 c3655(
.A(net2862),
.ZN(net3829)
);

INV_X1 c3656(
.A(net1931),
.ZN(net3830)
);

CLKGATETST_X2 c3657(
.E(net999),
.SE(net2932),
.CK(clk),
.GCK(net3831)
);

NAND2_X4 c3658(
.A1(net3826),
.A2(net3827),
.ZN(net3832)
);

AND2_X2 c3659(
.A1(net1903),
.A2(net2882),
.ZN(net3833)
);

INV_X2 c3660(
.A(net2932),
.ZN(net3834)
);

INV_X8 c3661(
.A(net3829),
.ZN(net3835)
);

XOR2_X1 c3662(
.A(net3835),
.B(net1008),
.Z(net3836)
);

NOR2_X1 c3663(
.A1(net942),
.A2(net3835),
.ZN(net3837)
);

INV_X16 c3664(
.A(net2868),
.ZN(net3838)
);

OR2_X2 c3665(
.A1(net1958),
.A2(net2942),
.ZN(net3839)
);

INV_X32 c3666(
.A(net29),
.ZN(net3840)
);

INV_X4 c3667(
.A(net3826),
.ZN(net3841)
);

NOR2_X4 c3668(
.A1(net3832),
.A2(net3838),
.ZN(net3842)
);

INV_X1 c3669(
.A(net3840),
.ZN(net3843)
);

INV_X2 c3670(
.A(net3827),
.ZN(net3844)
);

NOR2_X2 c3671(
.A1(net1977),
.A2(net3832),
.ZN(net3845)
);

INV_X8 c3672(
.A(net9773),
.ZN(net3846)
);

INV_X16 c3673(
.A(net9774),
.ZN(net3847)
);

INV_X32 c3674(
.A(net979),
.ZN(net3848)
);

INV_X4 c3675(
.A(net3846),
.ZN(net3849)
);

XOR2_X2 c3676(
.A(net3844),
.B(net3838),
.Z(net3850)
);

CLKGATETST_X4 c3677(
.E(net3842),
.SE(net3834),
.CK(clk),
.GCK(net3851)
);

XNOR2_X1 c3678(
.A(net3851),
.B(net2882),
.ZN(net3852)
);

INV_X1 c3679(
.A(net3841),
.ZN(net3853)
);

INV_X2 c3680(
.A(net1931),
.ZN(net3854)
);

CLKGATETST_X8 c3681(
.E(net2946),
.SE(net3841),
.CK(clk),
.GCK(net3855)
);

OR2_X4 c3682(
.A1(net3852),
.A2(net1961),
.ZN(net3856)
);

INV_X8 c3683(
.A(net9804),
.ZN(net3857)
);

INV_X16 c3684(
.A(net2910),
.ZN(net3858)
);

DFFR_X1 c3685(
.D(net3857),
.RN(net3850),
.CK(clk),
.Q(net3860),
.QN(net3859)
);

INV_X32 c3686(
.A(net1959),
.ZN(net3861)
);

DFFR_X2 c3687(
.D(net2864),
.RN(net3845),
.CK(clk),
.Q(net3863),
.QN(net3862)
);

INV_X4 c3688(
.A(net9815),
.ZN(net3864)
);

INV_X1 c3689(
.A(net3853),
.ZN(net3865)
);

DFFS_X1 c3690(
.D(net3835),
.SN(net3842),
.CK(clk),
.Q(net3867),
.QN(net3866)
);

INV_X2 c3691(
.A(net3867),
.ZN(net3868)
);

INV_X8 c3692(
.A(net3863),
.ZN(net3869)
);

INV_X16 c3693(
.A(net3869),
.ZN(net3870)
);

OR2_X1 c3694(
.A1(net930),
.A2(net3840),
.ZN(net3871)
);

INV_X32 c3695(
.A(net9814),
.ZN(net3872)
);

INV_X4 c3696(
.A(net3847),
.ZN(net3873)
);

INV_X1 c3697(
.A(net3849),
.ZN(net3874)
);

INV_X2 c3698(
.A(net10485),
.ZN(net3875)
);

XNOR2_X2 c3699(
.A(net1952),
.B(net3854),
.ZN(net3876)
);

AND2_X4 c3700(
.A1(net3873),
.A2(net2868),
.ZN(net3877)
);

INV_X8 c3701(
.A(net3867),
.ZN(net3878)
);

OR3_X1 c3702(
.A1(net2882),
.A2(net3862),
.A3(net3848),
.ZN(net3879)
);

AND2_X1 c3703(
.A1(net3840),
.A2(net3858),
.ZN(net3880)
);

SDFF_X2 c3704(
.D(net2922),
.SE(net3876),
.SI(net3853),
.CK(clk),
.Q(net3882),
.QN(net3881)
);

INV_X16 c3705(
.A(net3875),
.ZN(net3883)
);

INV_X32 c3706(
.A(net3871),
.ZN(net3884)
);

INV_X4 c3707(
.A(net3836),
.ZN(net3885)
);

NAND2_X1 c3708(
.A1(net3874),
.A2(net3870),
.ZN(net3886)
);

INV_X1 c3709(
.A(net10485),
.ZN(net3887)
);

AOI222_X1 c3710(
.A1(net3870),
.A2(net3873),
.B1(net3852),
.B2(net3857),
.C1(net3848),
.C2(net2868),
.ZN(net3888)
);

NAND2_X2 c3711(
.A1(net3870),
.A2(net3853),
.ZN(net3889)
);

AOI222_X4 c3712(
.A1(net3838),
.A2(net3869),
.B1(net3831),
.B2(net2882),
.C1(net3850),
.C2(net3848),
.ZN(net3890)
);

INV_X2 c3713(
.A(net3868),
.ZN(net3891)
);

NAND2_X4 c3714(
.A1(net3883),
.A2(net3861),
.ZN(net3892)
);

INV_X8 c3715(
.A(net9856),
.ZN(net3893)
);

INV_X16 c3716(
.A(net3889),
.ZN(net3894)
);

MUX2_X1 c3717(
.A(net3893),
.B(net3858),
.S(net3864),
.Z(net3895)
);

AND2_X2 c3718(
.A1(net3887),
.A2(net3866),
.ZN(net3896)
);

INV_X32 c3719(
.A(net9804),
.ZN(net3897)
);

XOR2_X1 c3720(
.A(net3888),
.B(net2882),
.Z(net3898)
);

NOR2_X1 c3721(
.A1(net3830),
.A2(net3874),
.ZN(net3899)
);

OR2_X2 c3722(
.A1(net2939),
.A2(net3850),
.ZN(net3900)
);

OAI21_X4 c3723(
.A(net3876),
.B1(net2910),
.B2(net2921),
.ZN(net3901)
);

NOR2_X4 c3724(
.A1(net3879),
.A2(net3864),
.ZN(net3902)
);

DFFS_X2 c3725(
.D(net3871),
.SN(net3884),
.CK(clk),
.Q(net3904),
.QN(net3903)
);

INV_X4 c3726(
.A(net3885),
.ZN(net3905)
);

INV_X1 c3727(
.A(net3882),
.ZN(net3906)
);

NOR2_X2 c3728(
.A1(net3840),
.A2(net10676),
.ZN(net3907)
);

MUX2_X2 c3729(
.A(net3891),
.B(net3865),
.S(net2898),
.Z(net3908)
);

XOR2_X2 c3730(
.A(net3895),
.B(net3898),
.Z(net3909)
);

XNOR2_X1 c3731(
.A(net3897),
.B(net3905),
.ZN(net3910)
);

NAND3_X4 c3732(
.A1(net3910),
.A2(net3888),
.A3(net3881),
.ZN(net3911)
);

OR2_X4 c3733(
.A1(net3902),
.A2(net10675),
.ZN(net3912)
);

OR2_X1 c3734(
.A1(net3909),
.A2(net3899),
.ZN(net3913)
);

INV_X2 c3735(
.A(net3014),
.ZN(net3914)
);

XNOR2_X2 c3736(
.A(net3037),
.B(net3884),
.ZN(net3915)
);

INV_X8 c3737(
.A(net2037),
.ZN(net3916)
);

AND2_X4 c3738(
.A1(net3017),
.A2(net2037),
.ZN(net3917)
);

INV_X16 c3739(
.A(net2983),
.ZN(net3918)
);

INV_X32 c3740(
.A(net10173),
.ZN(net3919)
);

OR3_X4 c3741(
.A1(net3012),
.A2(net2920),
.A3(net3016),
.ZN(net3920)
);

AND2_X1 c3742(
.A1(net2023),
.A2(net930),
.ZN(net3921)
);

AND3_X2 c3743(
.A1(net3896),
.A2(net3017),
.A3(net2023),
.ZN(net3922)
);

INV_X4 c3744(
.A(net3907),
.ZN(net3923)
);

INV_X1 c3745(
.A(net9618),
.ZN(net3924)
);

CLKGATETST_X1 c3746(
.E(net3861),
.SE(net1912),
.CK(clk),
.GCK(net3925)
);

CLKGATETST_X2 c3747(
.E(net3922),
.SE(net2998),
.CK(clk),
.GCK(net3926)
);

NAND2_X1 c3748(
.A1(net2986),
.A2(net3861),
.ZN(net3927)
);

NAND2_X2 c3749(
.A1(net3923),
.A2(net2943),
.ZN(net3928)
);

NAND2_X4 c3750(
.A1(net3872),
.A2(net2936),
.ZN(net3929)
);

AND2_X2 c3751(
.A1(net3916),
.A2(net2983),
.ZN(net3930)
);

INV_X2 c3752(
.A(net11175),
.ZN(net3931)
);

INV_X8 c3753(
.A(net10505),
.ZN(net3932)
);

INV_X16 c3754(
.A(net1102),
.ZN(net3933)
);

NOR3_X1 c3755(
.A1(net1097),
.A2(net2066),
.A3(net2986),
.ZN(net3934)
);

INV_X32 c3756(
.A(net10812),
.ZN(net3935)
);

OR3_X2 c3757(
.A1(net3926),
.A2(net3914),
.A3(net3911),
.ZN(net3936)
);

OAI21_X2 c3758(
.A(net2998),
.B1(net3013),
.B2(net3929),
.ZN(net3937)
);

INV_X4 c3759(
.A(net3902),
.ZN(net3938)
);

XOR2_X1 c3760(
.A(net3914),
.B(net10543),
.Z(net3939)
);

INV_X1 c3761(
.A(net2965),
.ZN(net3940)
);

NOR2_X1 c3762(
.A1(net2045),
.A2(net3929),
.ZN(net3941)
);

INV_X2 c3763(
.A(net3013),
.ZN(net3942)
);

INV_X8 c3764(
.A(net3905),
.ZN(net3943)
);

OR2_X2 c3765(
.A1(net3828),
.A2(net3925),
.ZN(net3944)
);

INV_X16 c3766(
.A(net1985),
.ZN(net3945)
);

INV_X32 c3767(
.A(net3938),
.ZN(net3946)
);

NOR2_X4 c3768(
.A1(net3936),
.A2(net10783),
.ZN(net3947)
);

OAI21_X1 c3769(
.A(net2972),
.B1(net3930),
.B2(net3013),
.ZN(net3948)
);

NOR2_X2 c3770(
.A1(net3937),
.A2(net3947),
.ZN(net3949)
);

XOR2_X2 c3771(
.A(net3940),
.B(net3902),
.Z(net3950)
);

INV_X4 c3772(
.A(net3935),
.ZN(net3951)
);

XNOR2_X1 c3773(
.A(net3000),
.B(net3013),
.ZN(net3952)
);

OR2_X4 c3774(
.A1(net3947),
.A2(net3952),
.ZN(net3953)
);

INV_X1 c3775(
.A(net3944),
.ZN(net3954)
);

OR2_X1 c3776(
.A1(net3951),
.A2(net3831),
.ZN(net3955)
);

INV_X2 c3777(
.A(net11124),
.ZN(net3956)
);

OR4_X1 c3778(
.A1(net3952),
.A2(net3892),
.A3(net2918),
.A4(net3911),
.ZN(net3957)
);

XNOR2_X2 c3779(
.A(net1008),
.B(net3937),
.ZN(net3958)
);

AOI21_X2 c3780(
.A(net1912),
.B1(net3829),
.B2(net1920),
.ZN(net3959)
);

INV_X8 c3781(
.A(net3955),
.ZN(net3960)
);

INV_X16 c3782(
.A(net3950),
.ZN(net3961)
);

CLKGATETST_X4 c3783(
.E(net3922),
.SE(net2965),
.CK(clk),
.GCK(net3962)
);

INV_X32 c3784(
.A(net9618),
.ZN(net3963)
);

AND2_X4 c3785(
.A1(net2936),
.A2(net10582),
.ZN(net3964)
);

AND2_X1 c3786(
.A1(net77),
.A2(net3957),
.ZN(net3965)
);

INV_X4 c3787(
.A(net10288),
.ZN(net3966)
);

INV_X1 c3788(
.A(net3924),
.ZN(net3967)
);

INV_X2 c3789(
.A(net3966),
.ZN(net3968)
);

NAND2_X1 c3790(
.A1(net3954),
.A2(net3947),
.ZN(net3969)
);

SDFFS_X1 c3791(
.D(net1903),
.SE(net3964),
.SI(net2983),
.SN(net3925),
.CK(clk),
.Q(net3971),
.QN(net3970)
);

NAND2_X2 c3792(
.A1(net3963),
.A2(net10505),
.ZN(net3972)
);

AOI21_X1 c3793(
.A(net2964),
.B1(net3970),
.B2(net2965),
.ZN(net3973)
);

NAND2_X4 c3794(
.A1(net2862),
.A2(net3848),
.ZN(net3974)
);

AOI21_X4 c3795(
.A(net3958),
.B1(net3967),
.B2(net11174),
.ZN(net3975)
);

SDFFS_X2 c3796(
.D(net3964),
.SE(net3966),
.SI(net3957),
.SN(net3850),
.CK(clk),
.Q(net3977),
.QN(net3976)
);

INV_X8 c3797(
.A(net10373),
.ZN(net3978)
);

AND2_X2 c3798(
.A1(net3914),
.A2(net3947),
.ZN(net3979)
);

AND3_X1 c3799(
.A1(net3932),
.A2(net3962),
.A3(net3930),
.ZN(net3980)
);

XOR2_X1 c3800(
.A(net3933),
.B(net3944),
.Z(net3981)
);

OAI33_X1 c3801(
.A1(net3968),
.A2(net3944),
.A3(net3934),
.B1(net3942),
.B2(net2046),
.B3(net3036),
.ZN(net3982)
);

INV_X16 c3802(
.A(net10171),
.ZN(net3983)
);

NAND3_X1 c3803(
.A1(net3942),
.A2(net3011),
.A3(net10582),
.ZN(net3984)
);

CLKGATETST_X8 c3804(
.E(net3949),
.SE(net3955),
.CK(clk),
.GCK(net3985)
);

NOR2_X1 c3805(
.A1(net3972),
.A2(net3926),
.ZN(net3986)
);

OR2_X2 c3806(
.A1(net3983),
.A2(net3976),
.ZN(net3987)
);

NOR2_X4 c3807(
.A1(net2982),
.A2(net3014),
.ZN(net3988)
);

NOR2_X2 c3808(
.A1(net3975),
.A2(net3919),
.ZN(net3989)
);

INV_X32 c3809(
.A(net10633),
.ZN(net3990)
);

XOR2_X2 c3810(
.A(net988),
.B(net3942),
.Z(net3991)
);

XNOR2_X1 c3811(
.A(net3991),
.B(net3924),
.ZN(net3992)
);

NOR3_X4 c3812(
.A1(net3987),
.A2(net3985),
.A3(net3957),
.ZN(net3993)
);

NOR3_X2 c3813(
.A1(net3973),
.A2(net3905),
.A3(net3989),
.ZN(net3994)
);

AND3_X4 c3814(
.A1(net3978),
.A2(net3989),
.A3(net3993),
.ZN(net3995)
);

NAND3_X2 c3815(
.A1(net3031),
.A2(net3993),
.A3(net10525),
.ZN(net3996)
);

OR2_X4 c3816(
.A1(net3939),
.A2(net10846),
.ZN(net3997)
);

OR3_X1 c3817(
.A1(net3985),
.A2(net3962),
.A3(net10846),
.ZN(net3998)
);

INV_X4 c3818(
.A(net9772),
.ZN(net3999)
);

OR2_X1 c3819(
.A1(net3089),
.A2(net2129),
.ZN(net4000)
);

XNOR2_X2 c3820(
.A(net3032),
.B(net3113),
.ZN(net4001)
);

AND2_X4 c3821(
.A1(net1157),
.A2(net2121),
.ZN(net4002)
);

AND2_X1 c3822(
.A1(net3071),
.A2(net3993),
.ZN(net4003)
);

NAND2_X1 c3823(
.A1(net3016),
.A2(net10950),
.ZN(net4004)
);

NAND2_X2 c3824(
.A1(net1158),
.A2(net3036),
.ZN(net4005)
);

NAND2_X4 c3825(
.A1(net3088),
.A2(net1125),
.ZN(net4006)
);

INV_X1 c3826(
.A(net3906),
.ZN(net4007)
);

AND2_X2 c3827(
.A1(net1176),
.A2(net3985),
.ZN(net4008)
);

INV_X2 c3828(
.A(net3993),
.ZN(net4009)
);

XOR2_X1 c3829(
.A(net1125),
.B(net3956),
.Z(net4010)
);

NOR2_X1 c3830(
.A1(net4010),
.A2(net2959),
.ZN(net4011)
);

OR2_X2 c3831(
.A1(net2056),
.A2(net2112),
.ZN(net4012)
);

INV_X8 c3832(
.A(net10458),
.ZN(net4013)
);

INV_X16 c3833(
.A(net9628),
.ZN(net4014)
);

INV_X32 c3834(
.A(net4012),
.ZN(net4015)
);

INV_X4 c3835(
.A(net10128),
.ZN(net4016)
);

NOR2_X4 c3836(
.A1(net3986),
.A2(net3989),
.ZN(net4017)
);

INV_X1 c3837(
.A(net11084),
.ZN(net4018)
);

NOR2_X2 c3838(
.A1(net3957),
.A2(net2959),
.ZN(net4019)
);

XOR2_X2 c3839(
.A(net4004),
.B(net3894),
.Z(net4020)
);

INV_X2 c3840(
.A(net10904),
.ZN(net4021)
);

INV_X8 c3841(
.A(net9628),
.ZN(net4022)
);

XNOR2_X1 c3842(
.A(net1898),
.B(net10542),
.ZN(net4023)
);

DFFR_X1 c3843(
.D(net3985),
.RN(net3989),
.CK(clk),
.Q(net4025),
.QN(net4024)
);

INV_X16 c3844(
.A(net9786),
.ZN(net4026)
);

OR2_X4 c3845(
.A1(net4023),
.A2(net11049),
.ZN(net4027)
);

OR2_X1 c3846(
.A1(net4021),
.A2(net3856),
.ZN(net4028)
);

INV_X32 c3847(
.A(net10851),
.ZN(net4029)
);

XNOR2_X2 c3848(
.A(net3045),
.B(net4025),
.ZN(net4030)
);

DFFR_X2 c3849(
.D(net4028),
.RN(net3117),
.CK(clk),
.Q(net4032),
.QN(net4031)
);

MUX2_X1 c3850(
.A(net3911),
.B(net3894),
.S(net3919),
.Z(net4033)
);

AND2_X4 c3851(
.A1(net4027),
.A2(net4015),
.ZN(net4034)
);

DFFRS_X1 c3852(
.D(net2046),
.RN(net3848),
.SN(net3036),
.CK(clk),
.Q(net4036),
.QN(net4035)
);

OAI21_X4 c3853(
.A(net4029),
.B1(net4033),
.B2(net4023),
.ZN(net4037)
);

INV_X4 c3854(
.A(net4000),
.ZN(net4038)
);

AND2_X1 c3855(
.A1(net4016),
.A2(net4019),
.ZN(net4039)
);

MUX2_X2 c3856(
.A(net4018),
.B(net4007),
.S(net3936),
.Z(net4040)
);

NAND2_X1 c3857(
.A1(net2090),
.A2(net4002),
.ZN(net4041)
);

NAND2_X2 c3858(
.A1(net4010),
.A2(net4035),
.ZN(net4042)
);

INV_X1 c3859(
.A(net4040),
.ZN(net4043)
);

NAND3_X4 c3860(
.A1(net4013),
.A2(net4020),
.A3(net4022),
.ZN(net4044)
);

OR3_X4 c3861(
.A1(net4014),
.A2(net4002),
.A3(net3931),
.ZN(net4045)
);

NAND2_X4 c3862(
.A1(net3963),
.A2(net3943),
.ZN(net4046)
);

INV_X2 c3863(
.A(net10850),
.ZN(net4047)
);

INV_X8 c3864(
.A(net4018),
.ZN(net4048)
);

INV_X16 c3865(
.A(net10833),
.ZN(net4049)
);

DFFS_X1 c3866(
.D(net4043),
.SN(net2943),
.CK(clk),
.Q(net4051),
.QN(net4050)
);

AND2_X2 c3867(
.A1(net4037),
.A2(net4013),
.ZN(net4052)
);

XOR2_X1 c3868(
.A(net4002),
.B(net4047),
.Z(net4053)
);

NOR2_X1 c3869(
.A1(net3931),
.A2(net11024),
.ZN(net4054)
);

INV_X32 c3870(
.A(net10868),
.ZN(net4055)
);

OR2_X2 c3871(
.A1(net4053),
.A2(net4029),
.ZN(net4056)
);

INV_X4 c3872(
.A(net11012),
.ZN(net4057)
);

INV_X1 c3873(
.A(net11024),
.ZN(net4058)
);

INV_X2 c3874(
.A(net11084),
.ZN(net4059)
);

AND3_X2 c3875(
.A1(net3894),
.A2(net4041),
.A3(net4059),
.ZN(net4060)
);

NOR2_X4 c3876(
.A1(net4046),
.A2(net3894),
.ZN(net4061)
);

NOR3_X1 c3877(
.A1(net4058),
.A2(net3072),
.A3(net4047),
.ZN(net4062)
);

NOR2_X2 c3878(
.A1(net3956),
.A2(net10904),
.ZN(net4063)
);

OR3_X2 c3879(
.A1(net2920),
.A2(net3965),
.A3(net4048),
.ZN(net4064)
);

AOI221_X1 c3880(
.A(net3997),
.B1(net4058),
.B2(net3921),
.C1(net4009),
.C2(net4024),
.ZN(net4065)
);

XOR2_X2 c3881(
.A(net4054),
.B(net3911),
.Z(net4066)
);

OAI21_X2 c3882(
.A(net4066),
.B1(net2112),
.B2(net3088),
.ZN(net4067)
);

OAI21_X1 c3883(
.A(net3074),
.B1(net4013),
.B2(net4048),
.ZN(net4068)
);

INV_X8 c3884(
.A(net10353),
.ZN(net4069)
);

XNOR2_X1 c3885(
.A(net4038),
.B(net4010),
.ZN(net4070)
);

AOI21_X2 c3886(
.A(net4069),
.B1(net4066),
.B2(net1177),
.ZN(net4071)
);

OR2_X4 c3887(
.A1(net4063),
.A2(net4035),
.ZN(net4072)
);

AOI21_X1 c3888(
.A(net4036),
.B1(net3016),
.B2(net4027),
.ZN(net4073)
);

AOI222_X2 c3889(
.A1(net4003),
.A2(net3060),
.B1(net4048),
.B2(net3108),
.C1(net3036),
.C2(net11086),
.ZN(net4074)
);

DFFRS_X2 c3890(
.D(net3977),
.RN(net3117),
.SN(net4049),
.CK(clk),
.Q(net4076),
.QN(net4075)
);

SDFF_X1 c3891(
.D(net4071),
.SE(net4014),
.SI(net4003),
.CK(clk),
.Q(net4078),
.QN(net4077)
);

INV_X16 c3892(
.A(net10259),
.ZN(net4079)
);

AOI21_X4 c3893(
.A(net4034),
.B1(net2920),
.B2(net4073),
.ZN(net4080)
);

OR2_X1 c3894(
.A1(net4079),
.A2(net11086),
.ZN(net4081)
);

OAI221_X1 c3895(
.A(net4049),
.B1(net4048),
.B2(net4028),
.C1(net3999),
.C2(net2121),
.ZN(net4082)
);

AND3_X1 c3896(
.A1(net3052),
.A2(net4081),
.A3(net11177),
.ZN(net4083)
);

OAI221_X4 c3897(
.A(net4033),
.B1(net4073),
.B2(net4081),
.C1(net4024),
.C2(net3925),
.ZN(net4084)
);

OAI22_X1 c3898(
.A1(net4044),
.A2(net4045),
.B1(net3957),
.B2(net11177),
.ZN(net4085)
);

XNOR2_X2 c3899(
.A(net4072),
.B(net11176),
.ZN(net4086)
);

NAND3_X1 c3900(
.A1(net4076),
.A2(net4086),
.A3(net10609),
.ZN(net4087)
);

AND2_X4 c3901(
.A1(net3106),
.A2(net4087),
.ZN(net4088)
);

AND2_X1 c3902(
.A1(net4061),
.A2(net3970),
.ZN(net4089)
);

INV_X32 c3903(
.A(net10841),
.ZN(net4090)
);

INV_X4 c3904(
.A(net10205),
.ZN(net4091)
);

NAND2_X1 c3905(
.A1(net2112),
.A2(net3210),
.ZN(net4092)
);

INV_X1 c3906(
.A(net4022),
.ZN(net4093)
);

NAND2_X2 c3907(
.A1(net85),
.A2(net2007),
.ZN(net4094)
);

NAND2_X4 c3908(
.A1(net1113),
.A2(net4050),
.ZN(net4095)
);

INV_X2 c3909(
.A(net11118),
.ZN(net4096)
);

AND2_X2 c3910(
.A1(net3115),
.A2(net3132),
.ZN(net4097)
);

XOR2_X1 c3911(
.A(net1927),
.B(net3971),
.Z(net4098)
);

NOR2_X1 c3912(
.A1(net2007),
.A2(net3195),
.ZN(net4099)
);

INV_X8 c3913(
.A(net4089),
.ZN(net4100)
);

INV_X16 c3914(
.A(net10315),
.ZN(net4101)
);

OR2_X2 c3915(
.A1(net3213),
.A2(net3101),
.ZN(net4102)
);

NOR2_X4 c3916(
.A1(net4006),
.A2(net3080),
.ZN(net4103)
);

INV_X32 c3917(
.A(net10978),
.ZN(net4104)
);

NOR2_X2 c3918(
.A1(net3143),
.A2(net3856),
.ZN(net4105)
);

XOR2_X2 c3919(
.A(net3036),
.B(net4019),
.Z(net4106)
);

XNOR2_X1 c3920(
.A(net2066),
.B(net4077),
.ZN(net4107)
);

NOR3_X4 c3921(
.A1(net3108),
.A2(net2066),
.A3(net3936),
.ZN(net4108)
);

NOR3_X2 c3922(
.A1(net4091),
.A2(net3859),
.A3(net2233),
.ZN(net4109)
);

OAI222_X1 c3923(
.A1(net3039),
.A2(net4099),
.B1(net1113),
.B2(net2066),
.C1(net4107),
.C2(net3187),
.ZN(net4110)
);

DFFS_X2 c3924(
.D(net3056),
.SN(net4100),
.CK(clk),
.Q(net4112),
.QN(net4111)
);

OR2_X4 c3925(
.A1(net4094),
.A2(net4104),
.ZN(net4113)
);

OR2_X1 c3926(
.A1(net3168),
.A2(net4107),
.ZN(net4114)
);

XNOR2_X2 c3927(
.A(net3999),
.B(net10521),
.ZN(net4115)
);

AND2_X4 c3928(
.A1(net4112),
.A2(net3859),
.ZN(net4116)
);

AND2_X1 c3929(
.A1(net4101),
.A2(net3935),
.ZN(net4117)
);

NAND2_X1 c3930(
.A1(net4117),
.A2(net11178),
.ZN(net4118)
);

AND3_X4 c3931(
.A1(net4112),
.A2(net2959),
.A3(net4107),
.ZN(net4119)
);

NAND2_X2 c3932(
.A1(net4102),
.A2(net4019),
.ZN(net4120)
);

NAND3_X2 c3933(
.A1(net3971),
.A2(net4118),
.A3(net11179),
.ZN(net4121)
);

OR3_X1 c3934(
.A1(net3119),
.A2(net1988),
.A3(net4121),
.ZN(net4122)
);

INV_X4 c3935(
.A(net10996),
.ZN(net4123)
);

INV_X1 c3936(
.A(net2199),
.ZN(net4124)
);

NAND2_X4 c3937(
.A1(net4088),
.A2(net3115),
.ZN(net4125)
);

AND2_X2 c3938(
.A1(net4116),
.A2(net4115),
.ZN(net4126)
);

XOR2_X1 c3939(
.A(net3007),
.B(net3016),
.Z(net4127)
);

MUX2_X1 c3940(
.A(net4042),
.B(net1203),
.S(net4047),
.Z(net4128)
);

INV_X2 c3941(
.A(net11124),
.ZN(net4129)
);

NOR2_X1 c3942(
.A1(net4124),
.A2(net1093),
.ZN(net4130)
);

OR2_X2 c3943(
.A1(net4105),
.A2(net11179),
.ZN(net4131)
);

INV_X8 c3944(
.A(net10317),
.ZN(net4132)
);

INV_X16 c3945(
.A(net10978),
.ZN(net4133)
);

NOR2_X4 c3946(
.A1(net4132),
.A2(net3159),
.ZN(net4134)
);

NOR2_X2 c3947(
.A1(net4133),
.A2(net4121),
.ZN(net4135)
);

XOR2_X2 c3948(
.A(net4104),
.B(net2166),
.Z(net4136)
);

XNOR2_X1 c3949(
.A(net4126),
.B(net4135),
.ZN(net4137)
);

OR2_X4 c3950(
.A1(net4135),
.A2(net4116),
.ZN(net4138)
);

INV_X32 c3951(
.A(net10907),
.ZN(net4139)
);

OR2_X1 c3952(
.A1(net3152),
.A2(net4123),
.ZN(net4140)
);

XNOR2_X2 c3953(
.A(net4055),
.B(net3992),
.ZN(net4141)
);

SDFF_X2 c3954(
.D(net4138),
.SE(net4107),
.SI(net3169),
.CK(clk),
.Q(net4143),
.QN(net4142)
);

AND2_X4 c3955(
.A1(net3132),
.A2(net4142),
.ZN(net4144)
);

AND2_X1 c3956(
.A1(net3205),
.A2(net11023),
.ZN(net4145)
);

NAND2_X1 c3957(
.A1(net4139),
.A2(net4022),
.ZN(net4146)
);

OAI21_X4 c3958(
.A(net4137),
.B1(net4136),
.B2(net4111),
.ZN(net4147)
);

INV_X4 c3959(
.A(net10812),
.ZN(net4148)
);

INV_X1 c3960(
.A(net10984),
.ZN(net4149)
);

NAND2_X2 c3961(
.A1(net4136),
.A2(net4019),
.ZN(net4150)
);

INV_X2 c3962(
.A(net11015),
.ZN(net4151)
);

NAND2_X4 c3963(
.A1(net4131),
.A2(net3913),
.ZN(net4152)
);

MUX2_X2 c3964(
.A(net4151),
.B(net4090),
.S(net2171),
.Z(net4153)
);

AND2_X2 c3965(
.A1(net3205),
.A2(net4133),
.ZN(net4154)
);

XOR2_X1 c3966(
.A(net3016),
.B(net4149),
.Z(net4155)
);

NAND3_X4 c3967(
.A1(net4144),
.A2(net4116),
.A3(net4154),
.ZN(net4156)
);

OR3_X4 c3968(
.A1(net4129),
.A2(net4138),
.A3(net4133),
.ZN(net4157)
);

NOR2_X1 c3969(
.A1(net4123),
.A2(net4146),
.ZN(net4158)
);

OR2_X2 c3970(
.A1(net4004),
.A2(net4137),
.ZN(net4159)
);

NOR2_X4 c3971(
.A1(net4025),
.A2(net10608),
.ZN(net4160)
);

INV_X8 c3972(
.A(net10997),
.ZN(net4161)
);

AND3_X2 c3973(
.A1(net4157),
.A2(net2121),
.A3(net4160),
.ZN(net4162)
);

NOR3_X1 c3974(
.A1(net4092),
.A2(net1251),
.A3(net4154),
.ZN(net4163)
);

OAI222_X4 c3975(
.A1(net4097),
.A2(net2229),
.B1(net4137),
.B2(net4099),
.C1(net4098),
.C2(net4107),
.ZN(net4164)
);

NOR2_X2 c3976(
.A1(net4125),
.A2(net4137),
.ZN(net4165)
);

OR3_X2 c3977(
.A1(net4162),
.A2(net4080),
.A3(net4150),
.ZN(net4166)
);

INV_X16 c3978(
.A(net10996),
.ZN(net4167)
);

OAI21_X2 c3979(
.A(net4124),
.B1(net4167),
.B2(net10915),
.ZN(net4168)
);

INV_X32 c3980(
.A(net9911),
.ZN(net4169)
);

OAI21_X1 c3981(
.A(net276),
.B1(net4157),
.B2(net4154),
.ZN(net4170)
);

INV_X4 c3982(
.A(net11118),
.ZN(net4171)
);

AOI21_X2 c3983(
.A(net4149),
.B1(net4161),
.B2(net10680),
.ZN(net4172)
);

XOR2_X2 c3984(
.A(net3159),
.B(net3936),
.Z(net4173)
);

INV_X1 c3985(
.A(net3300),
.ZN(net4174)
);

INV_X2 c3986(
.A(net10831),
.ZN(net4175)
);

OAI221_X2 c3987(
.A(net4143),
.B1(net4174),
.B2(net4050),
.C1(net4100),
.C2(net1200),
.ZN(net4176)
);

INV_X8 c3988(
.A(net10341),
.ZN(net4177)
);

XNOR2_X1 c3989(
.A(net2110),
.B(net3992),
.ZN(net4178)
);

AOI21_X1 c3990(
.A(net3281),
.B1(net3857),
.B2(net3279),
.ZN(net4179)
);

OR2_X4 c3991(
.A1(net4086),
.A2(net2245),
.ZN(net4180)
);

INV_X16 c3992(
.A(net9980),
.ZN(net4181)
);

OR2_X1 c3993(
.A1(net4158),
.A2(net3208),
.ZN(net4182)
);

INV_X32 c3994(
.A(net3284),
.ZN(net4183)
);

XNOR2_X2 c3995(
.A(net4078),
.B(net4175),
.ZN(net4184)
);

INV_X4 c3996(
.A(net4183),
.ZN(net4185)
);

AND2_X4 c3997(
.A1(net4173),
.A2(net3999),
.ZN(net4186)
);

AND2_X1 c3998(
.A1(net3243),
.A2(net1279),
.ZN(net4187)
);

AOI21_X4 c3999(
.A(net4178),
.B1(net3266),
.B2(net4173),
.ZN(net4188)
);

INV_X1 c4000(
.A(net3195),
.ZN(net4189)
);

INV_X2 c4001(
.A(net10526),
.ZN(net4190)
);

INV_X8 c4002(
.A(net11038),
.ZN(net4191)
);

INV_X16 c4003(
.A(net4115),
.ZN(net4192)
);

INV_X32 c4004(
.A(net2263),
.ZN(net4193)
);

NAND2_X1 c4005(
.A1(net1322),
.A2(net2284),
.ZN(net4194)
);

NAND2_X2 c4006(
.A1(net3936),
.A2(net4150),
.ZN(net4195)
);

INV_X4 c4007(
.A(net4020),
.ZN(net4196)
);

AND3_X1 c4008(
.A1(net4187),
.A2(net3300),
.A3(net10479),
.ZN(net4197)
);

NAND2_X4 c4009(
.A1(net3220),
.A2(net2121),
.ZN(net4198)
);

AND2_X2 c4010(
.A1(net4081),
.A2(net10732),
.ZN(net4199)
);

INV_X1 c4011(
.A(net3244),
.ZN(net4200)
);

INV_X2 c4012(
.A(net11038),
.ZN(net4201)
);

NAND3_X1 c4013(
.A1(net3992),
.A2(net3264),
.A3(net4194),
.ZN(net4202)
);

INV_X8 c4014(
.A(net10684),
.ZN(net4203)
);

XOR2_X1 c4015(
.A(net4200),
.B(net3281),
.Z(net4204)
);

NOR2_X1 c4016(
.A1(net4090),
.A2(net3277),
.ZN(net4205)
);

INV_X16 c4017(
.A(net10853),
.ZN(net4206)
);

NOR3_X4 c4018(
.A1(net4149),
.A2(net2245),
.A3(net10936),
.ZN(net4207)
);

INV_X32 c4019(
.A(net3264),
.ZN(net4208)
);

OR2_X2 c4020(
.A1(net4181),
.A2(net4194),
.ZN(net4209)
);

INV_X4 c4021(
.A(net4206),
.ZN(net4210)
);

NOR2_X4 c4022(
.A1(net3060),
.A2(net10915),
.ZN(net4211)
);

NOR3_X2 c4023(
.A1(net3279),
.A2(net4210),
.A3(net3216),
.ZN(net4212)
);

INV_X1 c4024(
.A(net10027),
.ZN(net4213)
);

NOR2_X2 c4025(
.A1(net3998),
.A2(net4200),
.ZN(net4214)
);

XOR2_X2 c4026(
.A(net4193),
.B(net4205),
.Z(net4215)
);

INV_X2 c4027(
.A(net4215),
.ZN(net4216)
);

INV_X8 c4028(
.A(net11024),
.ZN(net4217)
);

XNOR2_X1 c4029(
.A(net3261),
.B(net3257),
.ZN(net4218)
);

OR2_X4 c4030(
.A1(net4192),
.A2(net4175),
.ZN(net4219)
);

OR2_X1 c4031(
.A1(net4211),
.A2(net4214),
.ZN(net4220)
);

INV_X16 c4032(
.A(net10281),
.ZN(net4221)
);

XNOR2_X2 c4033(
.A(net4169),
.B(net4212),
.ZN(net4222)
);

AND2_X4 c4034(
.A1(net3856),
.A2(net4217),
.ZN(net4223)
);

DFFRS_X1 c4035(
.D(net4186),
.RN(net4098),
.SN(net4194),
.CK(clk),
.Q(net4225),
.QN(net4224)
);

AND2_X1 c4036(
.A1(net4171),
.A2(net4217),
.ZN(net4226)
);

AND3_X4 c4037(
.A1(net4081),
.A2(net4051),
.A3(net4193),
.ZN(net4227)
);

INV_X32 c4038(
.A(net10133),
.ZN(net4228)
);

NAND2_X1 c4039(
.A1(net4208),
.A2(net4096),
.ZN(net4229)
);

DFFRS_X2 c4040(
.D(net4224),
.RN(net4011),
.SN(net10521),
.CK(clk),
.Q(net4231),
.QN(net4230)
);

NAND3_X2 c4041(
.A1(net4187),
.A2(net2317),
.A3(net4224),
.ZN(net4232)
);

NAND2_X2 c4042(
.A1(net4218),
.A2(net4219),
.ZN(net4233)
);

NAND2_X4 c4043(
.A1(net4210),
.A2(net4222),
.ZN(net4234)
);

AND2_X2 c4044(
.A1(net4019),
.A2(net4212),
.ZN(net4235)
);

CLKGATETST_X1 c4045(
.E(net4194),
.SE(net4235),
.CK(clk),
.GCK(net4236)
);

OR3_X1 c4046(
.A1(net4236),
.A2(net4200),
.A3(net11013),
.ZN(net4237)
);

INV_X4 c4047(
.A(net9979),
.ZN(net4238)
);

AND4_X2 c4048(
.A1(net4238),
.A2(net4233),
.A3(net4213),
.A4(net4217),
.ZN(net4239)
);

MUX2_X1 c4049(
.A(net4239),
.B(net4203),
.S(net4237),
.Z(net4240)
);

OAI21_X4 c4050(
.A(net4180),
.B1(net4236),
.B2(net11013),
.ZN(net4241)
);

XOR2_X1 c4051(
.A(net3195),
.B(net10936),
.Z(net4242)
);

NOR2_X1 c4052(
.A1(net3215),
.A2(net2263),
.ZN(net4243)
);

MUX2_X2 c4053(
.A(net4155),
.B(net4235),
.S(net4194),
.Z(net4244)
);

OR2_X2 c4054(
.A1(net3118),
.A2(net4203),
.ZN(net4245)
);

SDFF_X1 c4055(
.D(net4107),
.SE(net4245),
.SI(net4236),
.CK(clk),
.Q(net4247),
.QN(net4246)
);

NAND3_X4 c4056(
.A1(net3266),
.A2(net4237),
.A3(net4213),
.ZN(net4248)
);

OR3_X4 c4057(
.A1(net4234),
.A2(net4231),
.A3(net4213),
.ZN(net4249)
);

SDFFR_X1 c4058(
.D(net4236),
.RN(net4134),
.SE(net4108),
.SI(net10569),
.CK(clk),
.Q(net4251),
.QN(net4250)
);

AND3_X2 c4059(
.A1(net4249),
.A2(net4217),
.A3(net4242),
.ZN(net4252)
);

NOR3_X1 c4060(
.A1(net4228),
.A2(net3122),
.A3(net4250),
.ZN(net4253)
);

OR3_X2 c4061(
.A1(net4247),
.A2(net4252),
.A3(net4108),
.ZN(net4254)
);

OAI21_X2 c4062(
.A(net4229),
.B1(net4219),
.B2(net4252),
.ZN(net4255)
);

SDFF_X2 c4063(
.D(net4252),
.SE(net4248),
.SI(net4242),
.CK(clk),
.Q(net4257),
.QN(net4256)
);

OAI222_X2 c4064(
.A1(net4253),
.A2(net4108),
.B1(net4246),
.B2(net4245),
.C1(net4203),
.C2(net4185),
.ZN(net4258)
);

OAI21_X1 c4065(
.A(net4197),
.B1(net4230),
.B2(net10732),
.ZN(net4259)
);

DFFRS_X1 c4066(
.D(net4108),
.RN(net4210),
.SN(net11074),
.CK(clk),
.Q(net4261),
.QN(net4260)
);

AOI222_X1 c4067(
.A1(net4326),
.A2(net3307),
.B1(net3364),
.B2(net4344),
.C1(net3292),
.C2(net2248),
.ZN(net4262)
);

NOR2_X4 c4068(
.A1(net4324),
.A2(net4344),
.ZN(net4263)
);

NOR2_X2 c4069(
.A1(net4343),
.A2(net4342),
.ZN(net4264)
);

XOR2_X2 c4070(
.A(net4319),
.B(net4300),
.Z(net4265)
);

DFFRS_X2 c4071(
.D(net4315),
.RN(net3364),
.SN(net3359),
.CK(clk),
.Q(net4267),
.QN(net4266)
);

AND4_X1 c4072(
.A1(net2233),
.A2(net4342),
.A3(net4302),
.A4(net4098),
.ZN(net4268)
);

AOI21_X2 c4073(
.A(net4248),
.B1(net4265),
.B2(net4293),
.ZN(net4269)
);

XNOR2_X1 c4074(
.A(net4346),
.B(net4300),
.ZN(net4270)
);

OR2_X4 c4075(
.A1(net4339),
.A2(net4310),
.ZN(net4271)
);

OR2_X1 c4076(
.A1(net4265),
.A2(net3333),
.ZN(net4272)
);

AOI21_X1 c4077(
.A(net4348),
.B1(net4272),
.B2(net4271),
.ZN(net4273)
);

AOI21_X4 c4078(
.A(net4337),
.B1(net4226),
.B2(net11004),
.ZN(net4274)
);

XNOR2_X2 c4079(
.A(net4323),
.B(net4189),
.ZN(net4275)
);

AND2_X4 c4080(
.A1(net4297),
.A2(net4233),
.ZN(net4276)
);

AND2_X1 c4081(
.A1(net4268),
.A2(net4344),
.ZN(net4277)
);

NAND2_X1 c4082(
.A1(net4264),
.A2(net4339),
.ZN(net4278)
);

NAND2_X2 c4083(
.A1(net4310),
.A2(net4272),
.ZN(net4279)
);

INV_X1 c4084(
.A(net4294),
.ZN(net4280)
);

CLKGATETST_X2 c4085(
.E(net4277),
.SE(net3348),
.CK(clk),
.GCK(net4281)
);

AND3_X1 c4086(
.A1(net3359),
.A2(net4268),
.A3(net4241),
.ZN(net4282)
);

NAND3_X1 c4087(
.A1(net4281),
.A2(net4294),
.A3(net4334),
.ZN(net4283)
);

NOR3_X4 c4088(
.A1(net4327),
.A2(net4317),
.A3(net4279),
.ZN(net4284)
);

INV_X2 c4089(
.A(net4308),
.ZN(net4285)
);

NAND2_X4 c4090(
.A1(net4274),
.A2(net3283),
.ZN(net4286)
);

AOI222_X4 c4091(
.A1(net4227),
.A2(net4266),
.B1(net3358),
.B2(net4237),
.C1(net4212),
.C2(net3376),
.ZN(net4287)
);

NOR3_X2 c4092(
.A1(net2349),
.A2(net4281),
.A3(net4286),
.ZN(net4288)
);

AND3_X4 c4093(
.A1(net4283),
.A2(net4309),
.A3(net11004),
.ZN(net4289)
);

NAND3_X2 c4094(
.A1(net4278),
.A2(net4283),
.A3(net4287),
.ZN(net4290)
);

OR3_X1 c4095(
.A1(net4278),
.A2(net4198),
.A3(net10989),
.ZN(net4291)
);

AND2_X2 c4096(
.A1(net4272),
.A2(net10989),
.ZN(net4292)
);

SDFF_X1 c4097(
.D(net3969),
.SE(net3375),
.SI(net10480),
.CK(clk),
.Q(net4294),
.QN(net4293)
);

XOR2_X1 c4098(
.A(net1898),
.B(net4237),
.Z(net4295)
);

NOR2_X1 c4099(
.A1(net4051),
.A2(net4212),
.ZN(net4296)
);

INV_X8 c4100(
.A(net4296),
.ZN(net4297)
);

INV_X16 c4101(
.A(net10781),
.ZN(net4298)
);

INV_X32 c4102(
.A(net2248),
.ZN(net4299)
);

INV_X4 c4103(
.A(net9611),
.ZN(net4300)
);

INV_X1 c4104(
.A(net9611),
.ZN(net4301)
);

INV_X2 c4105(
.A(net11078),
.ZN(net4302)
);

OR2_X2 c4106(
.A1(net3334),
.A2(net1236),
.ZN(net4303)
);

INV_X8 c4107(
.A(net3375),
.ZN(net4304)
);

INV_X16 c4108(
.A(net9722),
.ZN(net4305)
);

INV_X32 c4109(
.A(net10830),
.ZN(net4306)
);

NOR2_X4 c4110(
.A1(net4199),
.A2(net4212),
.ZN(net4307)
);

INV_X4 c4111(
.A(net4226),
.ZN(net4308)
);

NOR2_X2 c4112(
.A1(net3341),
.A2(net3357),
.ZN(net4309)
);

XOR2_X2 c4113(
.A(net4257),
.B(net1392),
.Z(net4310)
);

XNOR2_X1 c4114(
.A(net3384),
.B(net4298),
.ZN(net4311)
);

MUX2_X1 c4115(
.A(net3285),
.B(net4225),
.S(net3925),
.Z(net4312)
);

OR2_X4 c4116(
.A1(net4309),
.A2(net4256),
.ZN(net4313)
);

INV_X1 c4117(
.A(net3307),
.ZN(net4314)
);

OR2_X1 c4118(
.A1(net4221),
.A2(net4185),
.ZN(net4315)
);

INV_X2 c4119(
.A(net2348),
.ZN(net4316)
);

CLKGATETST_X4 c4120(
.E(net4315),
.SE(net4240),
.CK(clk),
.GCK(net4317)
);

OAI21_X4 c4121(
.A(net362),
.B1(net4308),
.B2(net4025),
.ZN(net4318)
);

XNOR2_X2 c4122(
.A(net4317),
.B(net4098),
.ZN(net4319)
);

MUX2_X2 c4123(
.A(net4243),
.B(net4315),
.S(net3384),
.Z(net4320)
);

NAND3_X4 c4124(
.A1(net3283),
.A2(net4219),
.A3(net2348),
.ZN(net4321)
);

AND2_X4 c4125(
.A1(net4308),
.A2(net2348),
.ZN(net4322)
);

INV_X8 c4126(
.A(net10191),
.ZN(net4323)
);

AOI22_X4 c4127(
.A1(net4306),
.A2(net3384),
.B1(net4321),
.B2(net2295),
.ZN(net4324)
);

AND2_X1 c4128(
.A1(net4299),
.A2(net3285),
.ZN(net4325)
);

NAND2_X1 c4129(
.A1(net4324),
.A2(net2376),
.ZN(net4326)
);

NAND2_X2 c4130(
.A1(net4219),
.A2(net4257),
.ZN(net4327)
);

INV_X16 c4131(
.A(net4322),
.ZN(net4328)
);

INV_X32 c4132(
.A(net4300),
.ZN(net4329)
);

NAND2_X4 c4133(
.A1(net3925),
.A2(net3341),
.ZN(net4330)
);

AND2_X2 c4134(
.A1(net4225),
.A2(net4316),
.ZN(net4331)
);

XOR2_X1 c4135(
.A(net4322),
.B(net4314),
.Z(net4332)
);

INV_X4 c4136(
.A(net10312),
.ZN(net4333)
);

NOR2_X1 c4137(
.A1(net1446),
.A2(net4319),
.ZN(net4334)
);

INV_X1 c4138(
.A(net10985),
.ZN(net4335)
);

INV_X2 c4139(
.A(net10831),
.ZN(net4336)
);

SDFF_X2 c4140(
.D(net4295),
.SE(net3306),
.SI(net2295),
.CK(clk),
.Q(net4338),
.QN(net4337)
);

INV_X8 c4141(
.A(net3333),
.ZN(net4339)
);

INV_X16 c4142(
.A(net9900),
.ZN(net4340)
);

DFFRS_X1 c4143(
.D(net1414),
.RN(net4332),
.SN(net3322),
.CK(clk),
.Q(net4342),
.QN(net4341)
);

OR2_X2 c4144(
.A1(net4212),
.A2(net4307),
.ZN(net4343)
);

NOR2_X4 c4145(
.A1(net4332),
.A2(net10691),
.ZN(net4344)
);

NOR2_X2 c4146(
.A1(net3316),
.A2(net2295),
.ZN(net4345)
);

XOR2_X2 c4147(
.A(net4307),
.B(net3210),
.Z(net4346)
);

XNOR2_X1 c4148(
.A(net4335),
.B(net460),
.ZN(net4347)
);

INV_X32 c4149(
.A(net10230),
.ZN(net4348)
);

INV_X4 c4150(
.A(net10157),
.ZN(net4349)
);

OR3_X4 c4151(
.A1(net4032),
.A2(net3358),
.A3(net10617),
.ZN(net4350)
);

INV_X1 c4152(
.A(net10905),
.ZN(net4351)
);

OR2_X4 c4153(
.A1(net3462),
.A2(net3471),
.ZN(net4352)
);

OR2_X1 c4154(
.A1(net3406),
.A2(net4347),
.ZN(net4353)
);

INV_X2 c4155(
.A(net4242),
.ZN(net4354)
);

XNOR2_X2 c4156(
.A(net3450),
.B(net4332),
.ZN(net4355)
);

AND2_X4 c4157(
.A1(net4271),
.A2(net4255),
.ZN(net4356)
);

INV_X8 c4158(
.A(net4316),
.ZN(net4357)
);

AND2_X1 c4159(
.A1(net3365),
.A2(net4270),
.ZN(net4358)
);

INV_X16 c4160(
.A(net4237),
.ZN(net4359)
);

INV_X32 c4161(
.A(net4286),
.ZN(net4360)
);

AND3_X2 c4162(
.A1(net4351),
.A2(net3471),
.A3(net4329),
.ZN(net4361)
);

NAND2_X1 c4163(
.A1(net3472),
.A2(net3348),
.ZN(net4362)
);

INV_X4 c4164(
.A(net10937),
.ZN(net4363)
);

NOR3_X1 c4165(
.A1(net4362),
.A2(net4287),
.A3(net4242),
.ZN(net4364)
);

OR3_X2 c4166(
.A1(net3411),
.A2(net4328),
.A3(net1493),
.ZN(net4365)
);

NAND2_X2 c4167(
.A1(net3408),
.A2(net2490),
.ZN(net4366)
);

NAND2_X4 c4168(
.A1(net4361),
.A2(net4298),
.ZN(net4367)
);

AND2_X2 c4169(
.A1(net4356),
.A2(net2433),
.ZN(net4368)
);

XOR2_X1 c4170(
.A(net4328),
.B(net4362),
.Z(net4369)
);

INV_X1 c4171(
.A(net459),
.ZN(net4370)
);

INV_X2 c4172(
.A(net10213),
.ZN(net4371)
);

NOR2_X1 c4173(
.A1(net4270),
.A2(net4363),
.ZN(net4372)
);

OR2_X2 c4174(
.A1(net4332),
.A2(net4333),
.ZN(net4373)
);

INV_X8 c4175(
.A(net3405),
.ZN(net4374)
);

INV_X16 c4176(
.A(net4305),
.ZN(net4375)
);

INV_X32 c4177(
.A(net10206),
.ZN(net4376)
);

INV_X4 c4178(
.A(net4366),
.ZN(net4377)
);

INV_X1 c4179(
.A(net9889),
.ZN(net4378)
);

INV_X2 c4180(
.A(net4292),
.ZN(net4379)
);

NOR2_X4 c4181(
.A1(net4376),
.A2(net4185),
.ZN(net4380)
);

NOR2_X2 c4182(
.A1(net3358),
.A2(net4185),
.ZN(net4381)
);

XOR2_X2 c4183(
.A(net4373),
.B(net4379),
.Z(net4382)
);

INV_X8 c4184(
.A(net4370),
.ZN(net4383)
);

OAI21_X2 c4185(
.A(net2449),
.B1(net1510),
.B2(net4379),
.ZN(net4384)
);

XNOR2_X1 c4186(
.A(net4354),
.B(net4360),
.ZN(net4385)
);

DFFRS_X2 c4187(
.D(net3427),
.RN(net4362),
.SN(net365),
.CK(clk),
.Q(net4387),
.QN(net4386)
);

INV_X16 c4188(
.A(net4355),
.ZN(net4388)
);

OR2_X4 c4189(
.A1(net2506),
.A2(net3471),
.ZN(net4389)
);

OAI21_X1 c4190(
.A(net3361),
.B1(net4316),
.B2(net3399),
.ZN(net4390)
);

AOI21_X2 c4191(
.A(net4385),
.B1(net3428),
.B2(net3411),
.ZN(net4391)
);

SDFF_X1 c4192(
.D(net2337),
.SE(net4368),
.SI(net4353),
.CK(clk),
.Q(net4393),
.QN(net4392)
);

OR2_X1 c4193(
.A1(net4387),
.A2(net4271),
.ZN(net4394)
);

XNOR2_X2 c4194(
.A(net4390),
.B(net4388),
.ZN(net4395)
);

AND2_X4 c4195(
.A1(net4391),
.A2(net11113),
.ZN(net4396)
);

AOI21_X1 c4196(
.A(net4370),
.B1(net4391),
.B2(net10731),
.ZN(net4397)
);

INV_X32 c4197(
.A(net10305),
.ZN(net4398)
);

INV_X4 c4198(
.A(net9781),
.ZN(net4399)
);

INV_X1 c4199(
.A(net4391),
.ZN(net4400)
);

AOI21_X4 c4200(
.A(net4381),
.B1(net4371),
.B2(net4242),
.ZN(net4401)
);

AND2_X1 c4201(
.A1(net4393),
.A2(net4378),
.ZN(net4402)
);

NAND2_X1 c4202(
.A1(net3460),
.A2(net11121),
.ZN(net4403)
);

INV_X2 c4203(
.A(net10028),
.ZN(net4404)
);

AND3_X1 c4204(
.A1(net4377),
.A2(net4160),
.A3(net4241),
.ZN(net4405)
);

NAND3_X1 c4205(
.A1(net4403),
.A2(net4391),
.A3(net4386),
.ZN(net4406)
);

NAND2_X2 c4206(
.A1(net4404),
.A2(net4385),
.ZN(net4407)
);

NOR3_X4 c4207(
.A1(net4282),
.A2(net4349),
.A3(net3365),
.ZN(net4408)
);

NAND2_X4 c4208(
.A1(net4405),
.A2(net4363),
.ZN(net4409)
);

AND2_X2 c4209(
.A1(net4357),
.A2(net4391),
.ZN(net4410)
);

SDFF_X2 c4210(
.D(net3216),
.SE(net4404),
.SI(net2484),
.CK(clk),
.Q(net4412),
.QN(net4411)
);

XOR2_X1 c4211(
.A(net4380),
.B(net4392),
.Z(net4413)
);

NOR2_X1 c4212(
.A1(net4388),
.A2(net10979),
.ZN(net4414)
);

INV_X8 c4213(
.A(net11115),
.ZN(net4415)
);

INV_X16 c4214(
.A(net10905),
.ZN(net4416)
);

AOI221_X4 c4215(
.A(net1398),
.B1(net4393),
.B2(net4413),
.C1(net3216),
.C2(net2425),
.ZN(net4417)
);

DFFRS_X1 c4216(
.D(net4349),
.RN(net3292),
.SN(net2317),
.CK(clk),
.Q(net4419),
.QN(net4418)
);

OR2_X2 c4217(
.A1(net4398),
.A2(net4399),
.ZN(net4420)
);

NOR3_X2 c4218(
.A1(net4399),
.A2(net4385),
.A3(net4420),
.ZN(net4421)
);

AND3_X4 c4219(
.A1(net4359),
.A2(net4409),
.A3(net4407),
.ZN(net4422)
);

NOR2_X4 c4220(
.A1(net4358),
.A2(net4409),
.ZN(net4423)
);

NOR2_X2 c4221(
.A1(net4406),
.A2(net4423),
.ZN(net4424)
);

NAND3_X2 c4222(
.A1(net4415),
.A2(net4387),
.A3(net4389),
.ZN(net4425)
);

OR3_X1 c4223(
.A1(net3428),
.A2(net4404),
.A3(net4411),
.ZN(net4426)
);

XOR2_X2 c4224(
.A(net4421),
.B(net4426),
.Z(net4427)
);

MUX2_X1 c4225(
.A(net4378),
.B(net4427),
.S(net3216),
.Z(net4428)
);

OAI21_X4 c4226(
.A(net4410),
.B1(net4423),
.B2(net11035),
.ZN(net4429)
);

XNOR2_X1 c4227(
.A(net4427),
.B(net4410),
.ZN(net4430)
);

MUX2_X2 c4228(
.A(net4412),
.B(net4430),
.S(net4425),
.Z(net4431)
);

OR2_X4 c4229(
.A1(net4370),
.A2(net11128),
.ZN(net4432)
);

NAND3_X4 c4230(
.A1(net4431),
.A2(net4427),
.A3(net4420),
.ZN(net4433)
);

DFFRS_X2 c4231(
.D(net4245),
.RN(net4426),
.SN(net4428),
.CK(clk),
.Q(net4435),
.QN(net4434)
);

OR3_X4 c4232(
.A1(net4429),
.A2(net4435),
.A3(net4432),
.ZN(net4436)
);

AND3_X2 c4233(
.A1(net4428),
.A2(net4255),
.A3(net1493),
.ZN(net4437)
);

INV_X32 c4234(
.A(net4407),
.ZN(net4438)
);

NOR3_X1 c4235(
.A1(net4233),
.A2(net3498),
.A3(net3554),
.ZN(net4439)
);

INV_X4 c4236(
.A(net3541),
.ZN(net4440)
);

INV_X1 c4237(
.A(net3460),
.ZN(net4441)
);

OR2_X1 c4238(
.A1(net4394),
.A2(net11180),
.ZN(net4442)
);

XNOR2_X2 c4239(
.A(net4426),
.B(net4424),
.ZN(net4443)
);

AND2_X4 c4240(
.A1(net3497),
.A2(net11171),
.ZN(net4444)
);

OR3_X2 c4241(
.A1(net2515),
.A2(net4395),
.A3(net645),
.ZN(net4445)
);

AND2_X1 c4242(
.A1(net3551),
.A2(net4407),
.ZN(net4446)
);

INV_X2 c4243(
.A(net4446),
.ZN(net4447)
);

OAI21_X2 c4244(
.A(net645),
.B1(net3550),
.B2(net2594),
.ZN(net4448)
);

NAND2_X1 c4245(
.A1(net3409),
.A2(net3497),
.ZN(net4449)
);

INV_X8 c4246(
.A(net11106),
.ZN(net4450)
);

NAND2_X2 c4247(
.A1(net2343),
.A2(net4365),
.ZN(net4451)
);

AOI221_X2 c4248(
.A(net4396),
.B1(net3493),
.B2(net2593),
.C1(net3544),
.C2(net11181),
.ZN(net4452)
);

NAND2_X4 c4249(
.A1(net581),
.A2(net4321),
.ZN(net4453)
);

AND2_X2 c4250(
.A1(net2496),
.A2(net4428),
.ZN(net4454)
);

XOR2_X1 c4251(
.A(net4365),
.B(net3505),
.Z(net4455)
);

INV_X16 c4252(
.A(net3422),
.ZN(net4456)
);

NOR2_X1 c4253(
.A1(net3292),
.A2(net4365),
.ZN(net4457)
);

INV_X32 c4254(
.A(net3517),
.ZN(net4458)
);

OR2_X2 c4255(
.A1(net1493),
.A2(net11180),
.ZN(net4459)
);

SDFFRS_X2 c4256(
.D(net4440),
.RN(net4437),
.SE(net3460),
.SI(net3292),
.SN(net3544),
.CK(clk),
.Q(net4461),
.QN(net4460)
);

NOR2_X4 c4257(
.A1(net4450),
.A2(net3548),
.ZN(net4462)
);

NOR2_X2 c4258(
.A1(net2531),
.A2(net3544),
.ZN(net4463)
);

OAI22_X4 c4259(
.A1(net1626),
.A2(net3535),
.B1(net3344),
.B2(net2557),
.ZN(net4464)
);

INV_X4 c4260(
.A(net4444),
.ZN(net4465)
);

XOR2_X2 c4261(
.A(net4447),
.B(net4438),
.Z(net4466)
);

INV_X1 c4262(
.A(net10126),
.ZN(net4467)
);

INV_X2 c4263(
.A(net4423),
.ZN(net4468)
);

INV_X8 c4264(
.A(net4314),
.ZN(net4469)
);

XNOR2_X1 c4265(
.A(net4401),
.B(net4442),
.ZN(net4470)
);

OR2_X4 c4266(
.A1(net4453),
.A2(net4241),
.ZN(net4471)
);

INV_X16 c4267(
.A(net2499),
.ZN(net4472)
);

INV_X32 c4268(
.A(net10099),
.ZN(net4473)
);

OR2_X1 c4269(
.A1(net4473),
.A2(net11049),
.ZN(net4474)
);

XNOR2_X2 c4270(
.A(net4466),
.B(net3517),
.ZN(net4475)
);

INV_X4 c4271(
.A(net10233),
.ZN(net4476)
);

AND2_X4 c4272(
.A1(net4389),
.A2(net4420),
.ZN(net4477)
);

AND2_X1 c4273(
.A1(net4459),
.A2(net4477),
.ZN(net4478)
);

NAND2_X1 c4274(
.A1(net3493),
.A2(net4477),
.ZN(net4479)
);

NAND2_X2 c4275(
.A1(net3477),
.A2(net4466),
.ZN(net4480)
);

NAND2_X4 c4276(
.A1(net4472),
.A2(net4463),
.ZN(net4481)
);

AND2_X2 c4277(
.A1(net4438),
.A2(net337),
.ZN(net4482)
);

INV_X1 c4278(
.A(net4448),
.ZN(net4483)
);

INV_X2 c4279(
.A(net4473),
.ZN(net4484)
);

SDFFR_X2 c4280(
.D(net4475),
.RN(net278),
.SE(net4438),
.SI(net3544),
.CK(clk),
.Q(net4486),
.QN(net4485)
);

INV_X8 c4281(
.A(net4465),
.ZN(net4487)
);

INV_X16 c4282(
.A(net11085),
.ZN(net4488)
);

XOR2_X1 c4283(
.A(net4458),
.B(net11049),
.Z(net4489)
);

NOR2_X1 c4284(
.A1(net4489),
.A2(net2346),
.ZN(net4490)
);

INV_X32 c4285(
.A(net10857),
.ZN(net4491)
);

OAI21_X1 c4286(
.A(net4442),
.B1(net4402),
.B2(net4389),
.ZN(net4492)
);

INV_X4 c4287(
.A(net4469),
.ZN(net4493)
);

OR2_X2 c4288(
.A1(net1510),
.A2(net4466),
.ZN(net4494)
);

INV_X1 c4289(
.A(net4468),
.ZN(net4495)
);

INV_X2 c4290(
.A(net10992),
.ZN(net4496)
);

AOI22_X2 c4291(
.A1(net4434),
.A2(net4478),
.B1(net4494),
.B2(net11113),
.ZN(net4497)
);

INV_X8 c4292(
.A(net10945),
.ZN(net4498)
);

NOR2_X4 c4293(
.A1(net4496),
.A2(net4379),
.ZN(net4499)
);

NOR2_X2 c4294(
.A1(net4483),
.A2(net4098),
.ZN(net4500)
);

AOI221_X1 c4295(
.A(net4490),
.B1(net3292),
.B2(net4498),
.C1(net3536),
.C2(net3544),
.ZN(net4501)
);

XOR2_X2 c4296(
.A(net4442),
.B(net10512),
.Z(net4502)
);

NAND4_X4 c4297(
.A1(net4488),
.A2(net3541),
.A3(net4424),
.A4(net3402),
.ZN(net4503)
);

AOI21_X2 c4298(
.A(net4493),
.B1(net3552),
.B2(net3369),
.ZN(net4504)
);

INV_X16 c4299(
.A(net10125),
.ZN(net4505)
);

INV_X32 c4300(
.A(net10270),
.ZN(net4506)
);

INV_X4 c4301(
.A(net11106),
.ZN(net4507)
);

SDFFS_X1 c4302(
.D(net4445),
.SE(net4495),
.SI(net4498),
.SN(net4476),
.CK(clk),
.Q(net4509),
.QN(net4508)
);

XNOR2_X1 c4303(
.A(net4486),
.B(net10672),
.ZN(net4510)
);

INV_X1 c4304(
.A(net11085),
.ZN(net4511)
);

AOI21_X1 c4305(
.A(net4452),
.B1(net4511),
.B2(net3292),
.ZN(net4512)
);

OAI211_X2 c4306(
.A(net4512),
.B(net4461),
.C1(net4476),
.C2(net4463),
.ZN(net4513)
);

INV_X2 c4307(
.A(net10256),
.ZN(net4514)
);

AOI21_X4 c4308(
.A(net4514),
.B1(net4511),
.B2(net4486),
.ZN(net4515)
);

OR2_X4 c4309(
.A1(net4482),
.A2(net11029),
.ZN(net4516)
);

OAI221_X1 c4310(
.A(net4498),
.B1(net4502),
.B2(net4473),
.C1(net4205),
.C2(net4479),
.ZN(net4517)
);

OR2_X1 c4311(
.A1(net4511),
.A2(net10798),
.ZN(net4518)
);

INV_X8 c4312(
.A(net10067),
.ZN(net4519)
);

XNOR2_X2 c4313(
.A(net4516),
.B(net4518),
.ZN(net4520)
);

OR4_X2 c4314(
.A1(net4519),
.A2(net4518),
.A3(net4502),
.A4(net4478),
.ZN(net4521)
);

AND2_X4 c4315(
.A1(net4498),
.A2(net11066),
.ZN(net4522)
);

CLKGATETST_X8 c4316(
.E(net1706),
.SE(net3640),
.CK(clk),
.GCK(net4523)
);

AND2_X1 c4317(
.A1(net4400),
.A2(net4463),
.ZN(net4524)
);

AND3_X1 c4318(
.A1(net3609),
.A2(net645),
.A3(net4463),
.ZN(net4525)
);

INV_X16 c4319(
.A(net3081),
.ZN(net4526)
);

INV_X32 c4320(
.A(net9612),
.ZN(net4527)
);

INV_X4 c4321(
.A(net11138),
.ZN(net4528)
);

INV_X1 c4322(
.A(net4505),
.ZN(net4529)
);

NAND3_X1 c4323(
.A1(net3630),
.A2(net4526),
.A3(net4457),
.ZN(net4530)
);

INV_X2 c4324(
.A(net4517),
.ZN(net4531)
);

INV_X8 c4325(
.A(net2644),
.ZN(net4532)
);

INV_X16 c4326(
.A(net11123),
.ZN(net4533)
);

INV_X32 c4327(
.A(net9737),
.ZN(net4534)
);

INV_X4 c4328(
.A(net3601),
.ZN(net4535)
);

NAND2_X1 c4329(
.A1(net4534),
.A2(net10462),
.ZN(net4536)
);

NAND2_X2 c4330(
.A1(net4523),
.A2(net4524),
.ZN(net4537)
);

INV_X1 c4331(
.A(net9737),
.ZN(net4538)
);

INV_X2 c4332(
.A(net11181),
.ZN(net4539)
);

INV_X8 c4333(
.A(net9736),
.ZN(net4540)
);

INV_X16 c4334(
.A(net4535),
.ZN(net4541)
);

INV_X32 c4335(
.A(net9736),
.ZN(net4542)
);

INV_X4 c4336(
.A(net3535),
.ZN(net4543)
);

INV_X1 c4337(
.A(net9728),
.ZN(net4544)
);

INV_X2 c4338(
.A(net11108),
.ZN(net4545)
);

INV_X8 c4339(
.A(net4532),
.ZN(net4546)
);

AOI211_X1 c4340(
.A(net3586),
.B(net4402),
.C1(net4459),
.C2(net4534),
.ZN(net4547)
);

NAND2_X4 c4341(
.A1(net1707),
.A2(net4505),
.ZN(net4548)
);

INV_X16 c4342(
.A(net4424),
.ZN(net4549)
);

INV_X32 c4343(
.A(net2624),
.ZN(net4550)
);

INV_X4 c4344(
.A(net4435),
.ZN(net4551)
);

AND2_X2 c4345(
.A1(net3611),
.A2(net3584),
.ZN(net4552)
);

INV_X1 c4346(
.A(net9690),
.ZN(net4553)
);

XOR2_X1 c4347(
.A(net4534),
.B(net10595),
.Z(net4554)
);

INV_X2 c4348(
.A(net4255),
.ZN(net4555)
);

NOR3_X4 c4349(
.A1(net4536),
.A2(net4476),
.A3(net4459),
.ZN(net4556)
);

NOR3_X2 c4350(
.A1(net684),
.A2(net4544),
.A3(net4437),
.ZN(net4557)
);

AND3_X4 c4351(
.A1(net4545),
.A2(net3584),
.A3(net4555),
.ZN(net4558)
);

INV_X8 c4352(
.A(net9690),
.ZN(net4559)
);

NOR2_X1 c4353(
.A1(net4463),
.A2(net4526),
.ZN(net4560)
);

INV_X16 c4354(
.A(net3589),
.ZN(net4561)
);

INV_X32 c4355(
.A(net10318),
.ZN(net4562)
);

INV_X4 c4356(
.A(net9848),
.ZN(net4563)
);

INV_X1 c4357(
.A(net11040),
.ZN(net4564)
);

OR2_X2 c4358(
.A1(net2661),
.A2(net4556),
.ZN(net4565)
);

NOR2_X4 c4359(
.A1(net4459),
.A2(net4375),
.ZN(net4566)
);

INV_X2 c4360(
.A(net4507),
.ZN(net4567)
);

NOR2_X2 c4361(
.A1(net2346),
.A2(net10747),
.ZN(net4568)
);

XOR2_X2 c4362(
.A(net715),
.B(net2632),
.Z(net4569)
);

XNOR2_X1 c4363(
.A(net4263),
.B(net4569),
.ZN(net4570)
);

INV_X8 c4364(
.A(net4568),
.ZN(net4571)
);

OR2_X4 c4365(
.A1(net4529),
.A2(net4538),
.ZN(net4572)
);

INV_X16 c4366(
.A(net10793),
.ZN(net4573)
);

INV_X32 c4367(
.A(net9881),
.ZN(net4574)
);

INV_X4 c4368(
.A(net10730),
.ZN(net4575)
);

INV_X1 c4369(
.A(net10692),
.ZN(net4576)
);

INV_X2 c4370(
.A(net4570),
.ZN(net4577)
);

INV_X8 c4371(
.A(net4555),
.ZN(net4578)
);

INV_X16 c4372(
.A(net4241),
.ZN(net4579)
);

OR2_X1 c4373(
.A1(net4561),
.A2(net4535),
.ZN(net4580)
);

XNOR2_X2 c4374(
.A(net3505),
.B(net3611),
.ZN(net4581)
);

INV_X32 c4375(
.A(net9612),
.ZN(net4582)
);

INV_X4 c4376(
.A(net4567),
.ZN(net4583)
);

OAI221_X4 c4377(
.A(net4575),
.B1(net2680),
.B2(net4573),
.C1(net4524),
.C2(net4432),
.ZN(net4584)
);

AND2_X4 c4378(
.A1(net4542),
.A2(net3641),
.ZN(net4585)
);

NAND3_X2 c4379(
.A1(net4543),
.A2(net4574),
.A3(net2558),
.ZN(net4586)
);

AND2_X1 c4380(
.A1(net4554),
.A2(net4425),
.ZN(net4587)
);

INV_X1 c4381(
.A(net4581),
.ZN(net4588)
);

OAI33_X1 c4382(
.A1(net4587),
.A2(net4273),
.A3(net4556),
.B1(net4463),
.B2(net3640),
.B3(net4528),
.ZN(net4589)
);

OR3_X1 c4383(
.A1(net4560),
.A2(net4585),
.A3(net4576),
.ZN(net4590)
);

MUX2_X1 c4384(
.A(net4553),
.B(net4575),
.S(net10605),
.Z(net4591)
);

INV_X2 c4385(
.A(net10913),
.ZN(net4592)
);

INV_X8 c4386(
.A(net11079),
.ZN(net4593)
);

NAND2_X1 c4387(
.A1(net4553),
.A2(net4579),
.ZN(net4594)
);

INV_X16 c4388(
.A(net11138),
.ZN(net4595)
);

NAND2_X2 c4389(
.A1(net4583),
.A2(net4594),
.ZN(net4596)
);

NAND2_X4 c4390(
.A1(net4538),
.A2(net4579),
.ZN(net4597)
);

OAI21_X4 c4391(
.A(net4580),
.B1(net4523),
.B2(net11109),
.ZN(net4598)
);

AND2_X2 c4392(
.A1(net4566),
.A2(net10944),
.ZN(net4599)
);

MUX2_X2 c4393(
.A(net1291),
.B(net4561),
.S(net10944),
.Z(net4600)
);

OAI221_X2 c4394(
.A(net4541),
.B1(net4255),
.B2(net4505),
.C1(net4544),
.C2(net3565),
.ZN(net4601)
);

AOI221_X4 c4395(
.A(net2632),
.B1(net4577),
.B2(net4600),
.C1(net4463),
.C2(net11133),
.ZN(net4602)
);

NAND4_X2 c4396(
.A1(net4592),
.A2(net4596),
.A3(net4534),
.A4(net4600),
.ZN(net4603)
);

NAND3_X4 c4397(
.A1(net4576),
.A2(net4587),
.A3(net4600),
.ZN(net4604)
);

AOI222_X2 c4398(
.A1(net4593),
.A2(net4592),
.B1(net4601),
.B2(net4550),
.C1(net4556),
.C2(net4600),
.ZN(net4605)
);

OR3_X4 c4399(
.A1(net3695),
.A2(net4479),
.A3(net3715),
.ZN(net4606)
);

XOR2_X1 c4400(
.A(net4509),
.B(net4273),
.Z(net4607)
);

SDFF_X1 c4401(
.D(net2570),
.SE(net2766),
.SI(net10793),
.CK(clk),
.Q(net4609),
.QN(net4608)
);

INV_X32 c4402(
.A(net4367),
.ZN(net4610)
);

NOR2_X1 c4403(
.A1(net2724),
.A2(net2633),
.ZN(out1)
);

OR2_X2 c4404(
.A1(net2633),
.A2(net1616),
.ZN(net4611)
);

INV_X4 c4405(
.A(net11112),
.ZN(net4612)
);

NOR2_X4 c4406(
.A1(net4611),
.A2(net10444),
.ZN(net4613)
);

NOR2_X2 c4407(
.A1(net4526),
.A2(net4579),
.ZN(net4614)
);

XOR2_X2 c4408(
.A(net4607),
.B(net3575),
.Z(net4615)
);

INV_X1 c4409(
.A(net9990),
.ZN(net4616)
);

INV_X2 c4410(
.A(net1793),
.ZN(net4617)
);

DFFR_X1 c4411(
.D(net3584),
.RN(net3715),
.CK(clk),
.Q(net4619),
.QN(net4618)
);

XNOR2_X1 c4412(
.A(net4571),
.B(net1720),
.ZN(net4620)
);

INV_X8 c4413(
.A(net11055),
.ZN(net4621)
);

OR2_X4 c4414(
.A1(net4586),
.A2(net4479),
.ZN(net4622)
);

OR2_X1 c4415(
.A1(net4621),
.A2(net4616),
.ZN(net4623)
);

XNOR2_X2 c4416(
.A(net3568),
.B(net4601),
.ZN(net4624)
);

AND2_X4 c4417(
.A1(net2766),
.A2(net3491),
.ZN(net4625)
);

AND2_X1 c4418(
.A1(net689),
.A2(net1720),
.ZN(net4626)
);

AND3_X2 c4419(
.A1(net3677),
.A2(net4604),
.A3(net689),
.ZN(net4627)
);

INV_X16 c4420(
.A(net11044),
.ZN(net4628)
);

NAND2_X1 c4421(
.A1(net4522),
.A2(net689),
.ZN(net4629)
);

NOR3_X1 c4422(
.A1(net4622),
.A2(net1616),
.A3(net4260),
.ZN(net4630)
);

NAND2_X2 c4423(
.A1(net3700),
.A2(net814),
.ZN(net4631)
);

NAND2_X4 c4424(
.A1(net4579),
.A2(net4625),
.ZN(net4632)
);

OR3_X2 c4425(
.A1(net682),
.A2(net4611),
.A3(net4617),
.ZN(net4633)
);

INV_X32 c4426(
.A(net9756),
.ZN(net4634)
);

OAI21_X2 c4427(
.A(net4321),
.B1(net1793),
.B2(net4550),
.ZN(net4635)
);

INV_X4 c4428(
.A(net1667),
.ZN(net4636)
);

AND2_X2 c4429(
.A1(net2521),
.A2(net4526),
.ZN(net4637)
);

SDFF_X2 c4430(
.D(net3728),
.SE(net773),
.SI(net1542),
.CK(clk),
.Q(net4639),
.QN(net4638)
);

XOR2_X1 c4431(
.A(net814),
.B(net4629),
.Z(net4640)
);

NOR2_X1 c4432(
.A1(net3494),
.A2(net4636),
.ZN(net4641)
);

OR4_X4 c4433(
.A1(net3686),
.A2(net2680),
.A3(net4608),
.A4(net4508),
.ZN(net4642)
);

OR2_X2 c4434(
.A1(net4625),
.A2(net4633),
.ZN(net4643)
);

NOR2_X4 c4435(
.A1(net798),
.A2(net2759),
.ZN(net4644)
);

NOR2_X2 c4436(
.A1(net2425),
.A2(net4616),
.ZN(net4645)
);

INV_X1 c4437(
.A(net9986),
.ZN(net4646)
);

XOR2_X2 c4438(
.A(net4626),
.B(net3713),
.Z(net4647)
);

INV_X2 c4439(
.A(net11009),
.ZN(net4648)
);

XNOR2_X1 c4440(
.A(net4617),
.B(net3672),
.ZN(net4649)
);

DFFRS_X1 c4441(
.D(net3721),
.RN(net4610),
.SN(net3691),
.CK(clk),
.Q(net4651),
.QN(net4650)
);

OAI22_X2 c4442(
.A1(net4628),
.A2(net2731),
.B1(net4610),
.B2(net4640),
.ZN(net4652)
);

OR2_X4 c4443(
.A1(net1768),
.A2(net4375),
.ZN(net4653)
);

OR2_X1 c4444(
.A1(net4606),
.A2(net4609),
.ZN(net4654)
);

XNOR2_X2 c4445(
.A(net3491),
.B(net4649),
.ZN(net4655)
);

AND2_X4 c4446(
.A1(net4620),
.A2(net10395),
.ZN(net4656)
);

OAI21_X1 c4447(
.A(net2472),
.B1(net2633),
.B2(net4651),
.ZN(net4657)
);

AND2_X1 c4448(
.A1(net4634),
.A2(net4655),
.ZN(net4658)
);

NAND2_X1 c4449(
.A1(net4634),
.A2(net11133),
.ZN(net4659)
);

AOI21_X2 c4450(
.A(net4654),
.B1(net4647),
.B2(net4594),
.ZN(net4660)
);

NAND2_X2 c4451(
.A1(net4630),
.A2(net4653),
.ZN(net4661)
);

AOI21_X1 c4452(
.A(net4658),
.B1(net4659),
.B2(net4616),
.ZN(net4662)
);

INV_X8 c4453(
.A(net9795),
.ZN(net4663)
);

DFFRS_X2 c4454(
.D(net4487),
.RN(net4662),
.SN(net3723),
.CK(clk),
.Q(net4665),
.QN(net4664)
);

AOI21_X4 c4455(
.A(net4613),
.B1(net4664),
.B2(net4617),
.ZN(net4666)
);

NAND2_X4 c4456(
.A1(net2700),
.A2(net4664),
.ZN(net4667)
);

AND3_X1 c4457(
.A1(net4642),
.A2(net4586),
.A3(net4651),
.ZN(net4668)
);

SDFF_X1 c4458(
.D(net4524),
.SE(net4659),
.SI(net4619),
.CK(clk),
.Q(net4670),
.QN(net4669)
);

NAND3_X1 c4459(
.A1(net4637),
.A2(net4616),
.A3(net4653),
.ZN(net4671)
);

AND2_X2 c4460(
.A1(net4641),
.A2(net4671),
.ZN(net4672)
);

NOR3_X4 c4461(
.A1(net2665),
.A2(net4667),
.A3(net4606),
.ZN(net4673)
);

SDFF_X2 c4462(
.D(net4662),
.SE(net1779),
.SI(net4670),
.CK(clk),
.Q(net4675),
.QN(net4674)
);

XOR2_X1 c4463(
.A(net4632),
.B(net4669),
.Z(net4676)
);

DFFRS_X1 c4464(
.D(net4647),
.RN(net4673),
.SN(net4676),
.CK(clk),
.Q(net4678),
.QN(net4677)
);

AOI221_X2 c4465(
.A(net4631),
.B1(net4609),
.B2(net4677),
.C1(net3565),
.C2(net4620),
.ZN(net4679)
);

NOR3_X2 c4466(
.A1(net4645),
.A2(net4673),
.A3(net4677),
.ZN(net4680)
);

AND3_X4 c4467(
.A1(net4657),
.A2(net2696),
.A3(net1720),
.ZN(net4681)
);

NAND3_X2 c4468(
.A1(net4644),
.A2(net4674),
.A3(net4668),
.ZN(net4682)
);

OR3_X1 c4469(
.A1(net4670),
.A2(net4675),
.A3(net4679),
.ZN(net4683)
);

NOR2_X1 c4470(
.A1(net4679),
.A2(net4646),
.ZN(net4684)
);

MUX2_X1 c4471(
.A(net4684),
.B(net4683),
.S(net3677),
.Z(net4685)
);

INV_X16 c4472(
.A(net11112),
.ZN(net4686)
);

OAI21_X4 c4473(
.A(net2731),
.B1(net4614),
.B2(net4659),
.ZN(net4687)
);

MUX2_X2 c4474(
.A(net4682),
.B(net4620),
.S(net4634),
.Z(net4688)
);

OR2_X2 c4475(
.A1(net4686),
.A2(net4639),
.ZN(net4689)
);

NOR2_X4 c4476(
.A1(net4375),
.A2(net4663),
.ZN(net4690)
);

NAND3_X4 c4477(
.A1(net3694),
.A2(net4676),
.A3(net4655),
.ZN(net4691)
);

SDFFS_X2 c4478(
.D(net4585),
.SE(net4674),
.SI(net4691),
.SN(net10756),
.CK(clk),
.Q(net4693),
.QN(net4692)
);

OR3_X4 c4479(
.A1(net4666),
.A2(net4693),
.A3(net10693),
.ZN(net4694)
);

OAI211_X4 c4480(
.A(net4690),
.B(net4694),
.C1(net4691),
.C2(net4601),
.ZN(net4695)
);

OAI211_X1 c4481(
.A(net4688),
.B(net4679),
.C1(net4691),
.C2(net10797),
.ZN(net4696)
);

NOR2_X2 c4482(
.A1(net3619),
.A2(net2782),
.ZN(net4697)
);

XOR2_X2 c4483(
.A(net3615),
.B(net807),
.Z(net4698)
);

XNOR2_X1 c4484(
.A(net3646),
.B(net3802),
.ZN(net4699)
);

OR2_X4 c4485(
.A1(net708),
.A2(net1816),
.ZN(net4700)
);

AND3_X2 c4486(
.A1(net4564),
.A2(net851),
.A3(net4692),
.ZN(net4701)
);

OR2_X1 c4487(
.A1(net2680),
.A2(net3797),
.ZN(net4702)
);

NOR3_X1 c4488(
.A1(net3757),
.A2(net3797),
.A3(net4668),
.ZN(net4703)
);

XNOR2_X2 c4489(
.A(net4652),
.B(net2849),
.ZN(net4704)
);

OR3_X2 c4490(
.A1(net3773),
.A2(net3757),
.A3(net4528),
.ZN(net4705)
);

DFFRS_X2 c4491(
.D(net2789),
.RN(net3803),
.SN(net3699),
.CK(clk),
.Q(net4707),
.QN(net4706)
);

OAI21_X2 c4492(
.A(net3803),
.B1(net4693),
.B2(net2809),
.ZN(net4708)
);

INV_X32 c4493(
.A(net9602),
.ZN(net4709)
);

OAI21_X1 c4494(
.A(net3620),
.B1(net2838),
.B2(net3646),
.ZN(net4710)
);

AND2_X4 c4495(
.A1(net851),
.A2(net3729),
.ZN(net4711)
);

AND2_X1 c4496(
.A1(net2815),
.A2(net2837),
.ZN(net4712)
);

NAND2_X1 c4497(
.A1(net3747),
.A2(net2815),
.ZN(net4713)
);

AOI21_X2 c4498(
.A(net4462),
.B1(net3774),
.B2(net10594),
.ZN(net4714)
);

AOI21_X1 c4499(
.A(net3805),
.B1(net3788),
.B2(net867),
.ZN(net4715)
);

AOI21_X4 c4500(
.A(net3676),
.B1(net4711),
.B2(net4652),
.ZN(net4716)
);

NAND2_X2 c4501(
.A1(net4643),
.A2(net3768),
.ZN(net4717)
);

NAND2_X4 c4502(
.A1(net4528),
.A2(net10822),
.ZN(net4718)
);

INV_X4 c4503(
.A(net10301),
.ZN(net4719)
);

AND3_X1 c4504(
.A1(net3750),
.A2(net3676),
.A3(net3794),
.ZN(net4720)
);

NAND3_X1 c4505(
.A1(net2777),
.A2(net3821),
.A3(net3737),
.ZN(net4721)
);

DFFR_X2 c4506(
.D(net4602),
.RN(net3699),
.CK(clk),
.Q(net4723),
.QN(net4722)
);

NOR3_X4 c4507(
.A1(net2837),
.A2(out1),
.A3(net4329),
.ZN(net4724)
);

NOR4_X4 c4508(
.A1(net4709),
.A2(net1779),
.A3(net773),
.A4(net3809),
.ZN(net4725)
);

NOR3_X2 c4509(
.A1(net773),
.A2(net4706),
.A3(net3737),
.ZN(net4726)
);

SDFF_X1 c4510(
.D(net3742),
.SE(net3741),
.SI(net4528),
.CK(clk),
.Q(net4728),
.QN(net4727)
);

AND3_X4 c4511(
.A1(net3798),
.A2(net3817),
.A3(net3782),
.ZN(net4729)
);

AND2_X2 c4512(
.A1(net905),
.A2(net3792),
.ZN(net4730)
);

SDFF_X2 c4513(
.D(net2834),
.SE(net4699),
.SI(net2849),
.CK(clk),
.Q(net4732),
.QN(net4731)
);

NAND3_X2 c4514(
.A1(net3729),
.A2(net4711),
.A3(net773),
.ZN(net4733)
);

NOR4_X2 c4515(
.A1(net4668),
.A2(net4713),
.A3(net3825),
.A4(net4731),
.ZN(net4734)
);

OR3_X1 c4516(
.A1(net3807),
.A2(net2808),
.A3(net3646),
.ZN(net4735)
);

XOR2_X1 c4517(
.A(net3716),
.B(net4732),
.Z(net4736)
);

NOR2_X1 c4518(
.A1(net4721),
.A2(net4698),
.ZN(net4737)
);

OR2_X2 c4519(
.A1(net4726),
.A2(net10648),
.ZN(net4738)
);

SDFFR_X1 c4520(
.D(net4697),
.RN(net1887),
.SE(net4652),
.SI(net2851),
.CK(clk),
.Q(net4740),
.QN(net4739)
);

MUX2_X1 c4521(
.A(net1836),
.B(net4738),
.S(net3798),
.Z(net4741)
);

AOI221_X1 c4522(
.A(net3708),
.B1(net4668),
.B2(net4711),
.C1(net4739),
.C2(net2712),
.ZN(net4742)
);

OAI21_X4 c4523(
.A(net2844),
.B1(net2686),
.B2(net4726),
.ZN(net4743)
);

MUX2_X2 c4524(
.A(net3618),
.B(net2712),
.S(net10448),
.Z(net4744)
);

NAND3_X4 c4525(
.A1(net3782),
.A2(net3807),
.A3(net2814),
.ZN(net4745)
);

OR3_X4 c4526(
.A1(net4726),
.A2(net4741),
.A3(net3785),
.ZN(net4746)
);

DFFRS_X1 c4527(
.D(net3811),
.RN(net4462),
.SN(net867),
.CK(clk),
.Q(net4748),
.QN(net4747)
);

NOR2_X4 c4528(
.A1(net3788),
.A2(net4732),
.ZN(net4749)
);

INV_X1 c4529(
.A(net9601),
.ZN(net4750)
);

AND3_X2 c4530(
.A1(net4703),
.A2(net3759),
.A3(net4476),
.ZN(net4751)
);

OAI222_X1 c4531(
.A1(net3741),
.A2(net3762),
.B1(net4731),
.B2(net3782),
.C1(net3742),
.C2(net3797),
.ZN(net4752)
);

NOR2_X2 c4532(
.A1(net4723),
.A2(net1887),
.ZN(net4753)
);

XOR2_X2 c4533(
.A(net1827),
.B(net2737),
.Z(net4754)
);

XNOR2_X1 c4534(
.A(net10563),
.B(net11183),
.ZN(net4755)
);

OR2_X4 c4535(
.A1(net4032),
.A2(net4749),
.ZN(net4756)
);

DFFRS_X2 c4536(
.D(net3614),
.RN(net4729),
.SN(net2791),
.CK(clk),
.Q(net4758),
.QN(net4757)
);

OR2_X1 c4537(
.A1(net3618),
.A2(net4758),
.ZN(net4759)
);

NOR3_X1 c4538(
.A1(net3667),
.A2(net3818),
.A3(net708),
.ZN(net4760)
);

OR3_X2 c4539(
.A1(net3774),
.A2(net4705),
.A3(net4755),
.ZN(net4761)
);

OAI21_X2 c4540(
.A(net3736),
.B1(net4755),
.B2(net4717),
.ZN(net4762)
);

OAI21_X1 c4541(
.A(net4730),
.B1(net4707),
.B2(net11182),
.ZN(net4763)
);

AOI21_X2 c4542(
.A(net3810),
.B1(net4732),
.B2(net4740),
.ZN(net4764)
);

OAI222_X4 c4543(
.A1(net2791),
.A2(net4640),
.B1(net4754),
.B2(net4739),
.C1(net2789),
.C2(net4755),
.ZN(net4765)
);

SDFF_X1 c4544(
.D(net4749),
.SE(net2851),
.SI(net4731),
.CK(clk),
.Q(net4767),
.QN(net4766)
);

AOI21_X1 c4545(
.A(net4718),
.B1(net4760),
.B2(net4722),
.ZN(net4768)
);

AOI21_X4 c4546(
.A(net4726),
.B1(net10787),
.B2(net11183),
.ZN(net4769)
);

AND3_X1 c4547(
.A1(net3769),
.A2(net4719),
.A3(net807),
.ZN(net4770)
);

NAND3_X1 c4548(
.A1(net4756),
.A2(net4770),
.A3(net11184),
.ZN(net4771)
);

NOR3_X4 c4549(
.A1(net3369),
.A2(net4707),
.A3(net828),
.ZN(net4772)
);

NOR3_X2 c4550(
.A1(net4701),
.A2(net4767),
.A3(net10788),
.ZN(net4773)
);

AND3_X4 c4551(
.A1(net4704),
.A2(net4733),
.A3(net4757),
.ZN(net4774)
);

SDFF_X2 c4552(
.D(net3778),
.SE(net3742),
.SI(net3811),
.CK(clk),
.Q(net4776),
.QN(net4775)
);

DFFRS_X1 c4553(
.D(net1844),
.RN(net4758),
.SN(net4755),
.CK(clk),
.Q(net4778),
.QN(net4777)
);

DFFRS_X2 c4554(
.D(net4764),
.RN(net4773),
.SN(net10447),
.CK(clk),
.Q(net4780),
.QN(net4779)
);

SDFF_X1 c4555(
.D(net2838),
.SE(net2851),
.SI(net3825),
.CK(clk),
.Q(net4782),
.QN(net4781)
);

NAND3_X2 c4556(
.A1(net4711),
.A2(net4750),
.A3(net4747),
.ZN(net4783)
);

OR3_X1 c4557(
.A1(net4743),
.A2(net10538),
.A3(net10823),
.ZN(net4784)
);

OAI222_X2 c4558(
.A1(net1879),
.A2(net4778),
.B1(net4754),
.B2(net4755),
.C1(net3797),
.C2(net3766),
.ZN(net4785)
);

MUX2_X1 c4559(
.A(net807),
.B(net4749),
.S(net4781),
.Z(net4786)
);

SDFF_X2 c4560(
.D(net4742),
.SE(net4784),
.SI(net4757),
.CK(clk),
.Q(net4788),
.QN(net4787)
);

OAI21_X4 c4561(
.A(net4788),
.B1(net4771),
.B2(net4782),
.ZN(net4789)
);

MUX2_X2 c4562(
.A(net4725),
.B(net4777),
.S(net10720),
.Z(net4790)
);

NAND3_X4 c4563(
.A1(net4790),
.A2(net4787),
.A3(net3758),
.ZN(net4791)
);

OR3_X4 c4564(
.A1(net3699),
.A2(net4789),
.A3(net10619),
.ZN(net4792)
);

INV_X2 c4565(
.A(net3831),
.ZN(net4793)
);

INV_X8 c4566(
.A(net3904),
.ZN(net4794)
);

INV_X16 c4567(
.A(net3858),
.ZN(net4795)
);

INV_X32 c4568(
.A(net3851),
.ZN(net4796)
);

XNOR2_X2 c4569(
.A(net1960),
.B(net3908),
.ZN(net4797)
);

INV_X4 c4570(
.A(net3849),
.ZN(net4798)
);

INV_X1 c4571(
.A(net1004),
.ZN(net4799)
);

INV_X2 c4572(
.A(net1962),
.ZN(net4800)
);

AND2_X4 c4573(
.A1(net1891),
.A2(in24),
.ZN(net4801)
);

INV_X8 c4574(
.A(net1008),
.ZN(net4802)
);

INV_X16 c4575(
.A(net3868),
.ZN(net4803)
);

INV_X32 c4576(
.A(net3908),
.ZN(net4804)
);

INV_X4 c4577(
.A(net3898),
.ZN(net4805)
);

INV_X1 c4578(
.A(net1908),
.ZN(net4806)
);

INV_X2 c4579(
.A(in7),
.ZN(net4807)
);

INV_X8 c4580(
.A(net3848),
.ZN(net4808)
);

INV_X16 c4581(
.A(net4801),
.ZN(net4809)
);

INV_X32 c4582(
.A(net3878),
.ZN(net4810)
);

AND2_X1 c4583(
.A1(net3855),
.A2(net3898),
.ZN(net4811)
);

INV_X4 c4584(
.A(net3886),
.ZN(net4812)
);

INV_X1 c4585(
.A(net1936),
.ZN(net4813)
);

INV_X2 c4586(
.A(net2919),
.ZN(net4814)
);

INV_X8 c4587(
.A(net3855),
.ZN(net4815)
);

NAND2_X1 c4588(
.A1(net4803),
.A2(net4815),
.ZN(net4816)
);

INV_X16 c4589(
.A(net2898),
.ZN(net4817)
);

INV_X32 c4590(
.A(net4811),
.ZN(net4818)
);

INV_X4 c4591(
.A(net4809),
.ZN(net4819)
);

NAND2_X2 c4592(
.A1(in24),
.A2(net3855),
.ZN(net4820)
);

INV_X1 c4593(
.A(net4794),
.ZN(net4821)
);

NAND2_X4 c4594(
.A1(net4795),
.A2(net4819),
.ZN(net4822)
);

INV_X2 c4595(
.A(net3858),
.ZN(net4823)
);

AND2_X2 c4596(
.A1(net4816),
.A2(net2880),
.ZN(net4824)
);

INV_X8 c4597(
.A(net4821),
.ZN(net4825)
);

XOR2_X1 c4598(
.A(net4818),
.B(net3913),
.Z(net4826)
);

NOR2_X1 c4599(
.A1(net4812),
.A2(net4817),
.ZN(net4827)
);

AND3_X2 c4600(
.A1(net4819),
.A2(net4820),
.A3(net4817),
.ZN(net4828)
);

INV_X16 c4601(
.A(net9544),
.ZN(net4829)
);

INV_X32 c4602(
.A(net3864),
.ZN(net4830)
);

OR2_X2 c4603(
.A1(net4810),
.A2(net4822),
.ZN(net4831)
);

NOR2_X4 c4604(
.A1(net4817),
.A2(net4804),
.ZN(net4832)
);

INV_X4 c4605(
.A(net4820),
.ZN(net4833)
);

NOR3_X1 c4606(
.A1(net4806),
.A2(net4809),
.A3(net4828),
.ZN(net4834)
);

NOR2_X2 c4607(
.A1(net2898),
.A2(net4832),
.ZN(net4835)
);

OR3_X2 c4608(
.A1(net4823),
.A2(net3877),
.A3(net4800),
.ZN(net4836)
);

OAI21_X2 c4609(
.A(net4812),
.B1(net4815),
.B2(net4823),
.ZN(net4837)
);

XOR2_X2 c4610(
.A(net4828),
.B(net4801),
.Z(net4838)
);

INV_X1 c4611(
.A(net2936),
.ZN(net4839)
);

DFFS_X1 c4612(
.D(net4826),
.SN(net4836),
.CK(clk),
.Q(net4841),
.QN(net4840)
);

INV_X2 c4613(
.A(net4825),
.ZN(net4842)
);

XNOR2_X1 c4614(
.A(net4831),
.B(net4825),
.ZN(net4843)
);

OR2_X4 c4615(
.A1(net4821),
.A2(net4822),
.ZN(net4844)
);

OR2_X1 c4616(
.A1(net4836),
.A2(net4795),
.ZN(net4845)
);

XNOR2_X2 c4617(
.A(net4842),
.B(net4830),
.ZN(net4846)
);

INV_X8 c4618(
.A(net9545),
.ZN(net4847)
);

AND2_X4 c4619(
.A1(net4794),
.A2(net3908),
.ZN(net4848)
);

AND2_X1 c4620(
.A1(net4848),
.A2(net4833),
.ZN(net4849)
);

NAND2_X1 c4621(
.A1(net4796),
.A2(net3903),
.ZN(net4850)
);

NAND2_X2 c4622(
.A1(net4837),
.A2(net3904),
.ZN(net4851)
);

NAND2_X4 c4623(
.A1(net4828),
.A2(net4851),
.ZN(net4852)
);

AND2_X2 c4624(
.A1(net3877),
.A2(net4852),
.ZN(net4853)
);

XOR2_X1 c4625(
.A(net4811),
.B(net4814),
.Z(net4854)
);

OAI21_X1 c4626(
.A(net4833),
.B1(net4797),
.B2(net4812),
.ZN(net4855)
);

AOI21_X2 c4627(
.A(net4847),
.B1(net3886),
.B2(net4855),
.ZN(net4856)
);

NOR2_X1 c4628(
.A1(net4853),
.A2(net4854),
.ZN(net4857)
);

OR2_X2 c4629(
.A1(net3834),
.A2(net4823),
.ZN(net4858)
);

NOR2_X4 c4630(
.A1(net4850),
.A2(net4851),
.ZN(net4859)
);

AOI21_X1 c4631(
.A(net4803),
.B1(net4845),
.B2(net10503),
.ZN(net4860)
);

DFFS_X2 c4632(
.D(net3878),
.SN(net4858),
.CK(clk),
.Q(net4862),
.QN(net4861)
);

AOI222_X1 c4633(
.A1(net4848),
.A2(net4815),
.B1(net4853),
.B2(net4861),
.C1(net4838),
.C2(net3850),
.ZN(net4863)
);

SDFFR_X2 c4634(
.D(net4793),
.RN(net4829),
.SE(net4858),
.SI(net3899),
.CK(clk),
.Q(net4865),
.QN(net4864)
);

AOI21_X4 c4635(
.A(net4862),
.B1(net4835),
.B2(net4817),
.ZN(net4866)
);

AND3_X1 c4636(
.A1(net4851),
.A2(net4860),
.A3(net4827),
.ZN(net4867)
);

NOR2_X2 c4637(
.A1(net4829),
.A2(net4859),
.ZN(net4868)
);

XOR2_X2 c4638(
.A(net4861),
.B(net10503),
.Z(net4869)
);

AOI211_X4 c4639(
.A(net4804),
.B(net4842),
.C1(net4812),
.C2(net3848),
.ZN(net4870)
);

XNOR2_X1 c4640(
.A(net4870),
.B(net3854),
.ZN(net4871)
);

SDFFS_X1 c4641(
.D(net4858),
.SE(net4868),
.SI(net4831),
.SN(net4871),
.CK(clk),
.Q(net4873),
.QN(net4872)
);

AOI222_X4 c4642(
.A1(net4867),
.A2(net4852),
.B1(net4872),
.B2(net4810),
.C1(net4845),
.C2(net3850),
.ZN(net4874)
);

OR2_X4 c4643(
.A1(net4855),
.A2(net4851),
.ZN(net4875)
);

OR2_X1 c4644(
.A1(net4860),
.A2(net4859),
.ZN(net4876)
);

DFFRS_X1 c4645(
.D(net4870),
.RN(net4876),
.SN(net11187),
.CK(clk),
.Q(net4878),
.QN(net4877)
);

DFFRS_X2 c4646(
.D(net4876),
.RN(net4864),
.SN(net11186),
.CK(clk),
.Q(net4880),
.QN(net4879)
);

SDFFRS_X1 c4647(
.D(net4875),
.RN(net4843),
.SE(net4876),
.SI(net4871),
.SN(net4802),
.CK(clk),
.Q(net4882),
.QN(net4881)
);

XNOR2_X2 c4648(
.A(net3929),
.B(net2958),
.ZN(net4883)
);

NAND3_X1 c4649(
.A1(net3961),
.A2(net4834),
.A3(net4822),
.ZN(net4884)
);

INV_X16 c4650(
.A(net3964),
.ZN(net4885)
);

NOR3_X4 c4651(
.A1(net2029),
.A2(net2880),
.A3(net3929),
.ZN(net4886)
);

INV_X32 c4652(
.A(net4822),
.ZN(net4887)
);

AND2_X4 c4653(
.A1(net3917),
.A2(net3919),
.ZN(net4888)
);

INV_X4 c4654(
.A(net3942),
.ZN(net4889)
);

INV_X1 c4655(
.A(net2064),
.ZN(net4890)
);

INV_X2 c4656(
.A(net10340),
.ZN(net4891)
);

INV_X8 c4657(
.A(net4890),
.ZN(net4892)
);

INV_X16 c4658(
.A(net4887),
.ZN(net4893)
);

INV_X32 c4659(
.A(net9663),
.ZN(net4894)
);

AND2_X1 c4660(
.A1(net4816),
.A2(net3854),
.ZN(net4895)
);

INV_X4 c4661(
.A(net3829),
.ZN(net4896)
);

NAND2_X1 c4662(
.A1(net3001),
.A2(net4834),
.ZN(net4897)
);

INV_X1 c4663(
.A(net9699),
.ZN(net4898)
);

INV_X2 c4664(
.A(net3945),
.ZN(net4899)
);

INV_X8 c4665(
.A(net4891),
.ZN(net4900)
);

NAND2_X2 c4666(
.A1(net2958),
.A2(net3031),
.ZN(net4901)
);

INV_X16 c4667(
.A(net4892),
.ZN(net4902)
);

CLKGATETST_X1 c4668(
.E(net4826),
.SE(net4827),
.CK(clk),
.GCK(net4903)
);

INV_X32 c4669(
.A(net10784),
.ZN(net4904)
);

SDFF_X1 c4670(
.D(net4886),
.SE(net4902),
.SI(net4899),
.CK(clk),
.Q(net4906),
.QN(net4905)
);

INV_X4 c4671(
.A(net3962),
.ZN(net4907)
);

INV_X1 c4672(
.A(net4869),
.ZN(net4908)
);

INV_X2 c4673(
.A(net4895),
.ZN(net4909)
);

NAND2_X4 c4674(
.A1(net4835),
.A2(net4852),
.ZN(net4910)
);

SDFF_X2 c4675(
.D(net4852),
.SE(net2049),
.SI(net4884),
.CK(clk),
.Q(net4912),
.QN(net4911)
);

INV_X8 c4676(
.A(net2936),
.ZN(net4913)
);

AND2_X2 c4677(
.A1(net4907),
.A2(net4904),
.ZN(net4914)
);

XOR2_X1 c4678(
.A(net4880),
.B(net4852),
.Z(net4915)
);

INV_X16 c4679(
.A(net4896),
.ZN(net4916)
);

NOR2_X1 c4680(
.A1(net2880),
.A2(net3892),
.ZN(net4917)
);

INV_X32 c4681(
.A(net1908),
.ZN(net4918)
);

OR2_X2 c4682(
.A1(net4878),
.A2(net3935),
.ZN(net4919)
);

NOR2_X4 c4683(
.A1(net4906),
.A2(net4903),
.ZN(net4920)
);

NOR2_X2 c4684(
.A1(net4920),
.A2(net2064),
.ZN(net4921)
);

INV_X4 c4685(
.A(net4862),
.ZN(net4922)
);

INV_X1 c4686(
.A(net4916),
.ZN(net4923)
);

INV_X2 c4687(
.A(net4914),
.ZN(net4924)
);

INV_X8 c4688(
.A(net2036),
.ZN(net4925)
);

XOR2_X2 c4689(
.A(net4900),
.B(net4921),
.Z(net4926)
);

CLKGATETST_X2 c4690(
.E(net4897),
.SE(net4919),
.CK(clk),
.GCK(net4927)
);

XNOR2_X1 c4691(
.A(net4926),
.B(net4802),
.ZN(net4928)
);

OR2_X4 c4692(
.A1(net4883),
.A2(net4928),
.ZN(net4929)
);

INV_X16 c4693(
.A(net10136),
.ZN(net4930)
);

INV_X32 c4694(
.A(net4815),
.ZN(net4931)
);

NOR3_X2 c4695(
.A1(net4921),
.A2(net4899),
.A3(net4905),
.ZN(net4932)
);

DFFRS_X1 c4696(
.D(net4924),
.RN(net2993),
.SN(net4909),
.CK(clk),
.Q(net4934),
.QN(net4933)
);

AND3_X4 c4697(
.A1(net3031),
.A2(net4859),
.A3(net4919),
.ZN(net4935)
);

INV_X4 c4698(
.A(net9663),
.ZN(net4936)
);

OR2_X1 c4699(
.A1(net4817),
.A2(net10694),
.ZN(net4937)
);

CLKGATETST_X4 c4700(
.E(net4925),
.SE(net4879),
.CK(clk),
.GCK(net4938)
);

INV_X1 c4701(
.A(net10445),
.ZN(net4939)
);

XNOR2_X2 c4702(
.A(net4884),
.B(net4802),
.ZN(net4940)
);

INV_X2 c4703(
.A(net10112),
.ZN(net4941)
);

INV_X8 c4704(
.A(net4932),
.ZN(net4942)
);

AND2_X4 c4705(
.A1(net4928),
.A2(net4929),
.ZN(net4943)
);

NAND3_X2 c4706(
.A1(net4941),
.A2(net4895),
.A3(net4925),
.ZN(net4944)
);

AND2_X1 c4707(
.A1(net4922),
.A2(net3892),
.ZN(net4945)
);

NAND2_X1 c4708(
.A1(net4906),
.A2(net10610),
.ZN(net4946)
);

INV_X16 c4709(
.A(net4913),
.ZN(net4947)
);

INV_X32 c4710(
.A(net4947),
.ZN(net4948)
);

NAND2_X2 c4711(
.A1(net4802),
.A2(net4937),
.ZN(net4949)
);

OR3_X1 c4712(
.A1(net4946),
.A2(net4938),
.A3(net4904),
.ZN(net4950)
);

INV_X4 c4713(
.A(net9927),
.ZN(net4951)
);

NAND2_X4 c4714(
.A1(net4918),
.A2(net4908),
.ZN(net4952)
);

AND2_X2 c4715(
.A1(net4949),
.A2(net4928),
.ZN(net4953)
);

INV_X1 c4716(
.A(net10784),
.ZN(net4954)
);

XOR2_X1 c4717(
.A(net4937),
.B(net4833),
.Z(net4955)
);

MUX2_X1 c4718(
.A(net4951),
.B(net3943),
.S(net10847),
.Z(net4956)
);

NOR2_X1 c4719(
.A1(net4955),
.A2(net4948),
.ZN(net4957)
);

OR2_X2 c4720(
.A1(net4948),
.A2(net4934),
.ZN(net4958)
);

NOR2_X4 c4721(
.A1(net4952),
.A2(net4907),
.ZN(net4959)
);

NOR2_X2 c4722(
.A1(net4902),
.A2(net3965),
.ZN(net4960)
);

OAI21_X4 c4723(
.A(net3831),
.B1(net4928),
.B2(net4951),
.ZN(net4961)
);

OAI33_X1 c4724(
.A1(net4920),
.A2(net4961),
.A3(net4890),
.B1(net4933),
.B2(net2993),
.B3(net4928),
.ZN(net4962)
);

XOR2_X2 c4725(
.A(net4959),
.B(net4948),
.Z(net4963)
);

DFFRS_X2 c4726(
.D(net4953),
.RN(net4946),
.SN(net3848),
.CK(clk),
.Q(net4965),
.QN(net4964)
);

XNOR2_X1 c4727(
.A(net4963),
.B(net4938),
.ZN(net4966)
);

MUX2_X2 c4728(
.A(net4960),
.B(net4877),
.S(net10783),
.Z(net4967)
);

AOI222_X2 c4729(
.A1(net4960),
.A2(net4966),
.B1(net4933),
.B2(net3925),
.C1(net4900),
.C2(net10446),
.ZN(net4968)
);

SDFF_X1 c4730(
.D(net4827),
.SE(net4966),
.SI(net4963),
.CK(clk),
.Q(net4970),
.QN(net4969)
);

OR2_X4 c4731(
.A1(net3108),
.A2(net1927),
.ZN(net4971)
);

OR2_X1 c4732(
.A1(net2098),
.A2(net4930),
.ZN(net4972)
);

XNOR2_X2 c4733(
.A(net4083),
.B(net4972),
.ZN(net4973)
);

AND2_X4 c4734(
.A1(net3854),
.A2(net11152),
.ZN(net4974)
);

AND2_X1 c4735(
.A1(net4888),
.A2(net3956),
.ZN(net4975)
);

INV_X2 c4736(
.A(net2032),
.ZN(net4976)
);

INV_X8 c4737(
.A(net2884),
.ZN(net4977)
);

INV_X16 c4738(
.A(net4800),
.ZN(net4978)
);

INV_X32 c4739(
.A(net3974),
.ZN(net4979)
);

INV_X4 c4740(
.A(net10352),
.ZN(net4980)
);

INV_X1 c4741(
.A(net3052),
.ZN(net4981)
);

NAND2_X1 c4742(
.A1(net4974),
.A2(net4899),
.ZN(net4982)
);

INV_X2 c4743(
.A(net4972),
.ZN(net4983)
);

NAND2_X2 c4744(
.A1(net4978),
.A2(net4911),
.ZN(net4984)
);

NAND2_X4 c4745(
.A1(net3943),
.A2(net11049),
.ZN(net4985)
);

AND2_X2 c4746(
.A1(net4976),
.A2(net2098),
.ZN(net4986)
);

INV_X8 c4747(
.A(net9874),
.ZN(net4987)
);

INV_X16 c4748(
.A(net4057),
.ZN(net4988)
);

INV_X32 c4749(
.A(net4984),
.ZN(net4989)
);

INV_X4 c4750(
.A(net10635),
.ZN(net4990)
);

XOR2_X1 c4751(
.A(net2129),
.B(net4007),
.Z(net4991)
);

INV_X1 c4752(
.A(net3929),
.ZN(net4992)
);

INV_X2 c4753(
.A(net4991),
.ZN(net4993)
);

NAND3_X4 c4754(
.A1(net4797),
.A2(net4992),
.A3(net3965),
.ZN(net4994)
);

NOR2_X1 c4755(
.A1(net4982),
.A2(net4992),
.ZN(net4995)
);

INV_X8 c4756(
.A(net9656),
.ZN(net4996)
);

INV_X16 c4757(
.A(net4973),
.ZN(net4997)
);

INV_X32 c4758(
.A(net10830),
.ZN(net4998)
);

INV_X4 c4759(
.A(net4993),
.ZN(net4999)
);

OR2_X2 c4760(
.A1(net4026),
.A2(net4992),
.ZN(net5000)
);

INV_X1 c4761(
.A(net4973),
.ZN(net5001)
);

NOR2_X4 c4762(
.A1(net4834),
.A2(net4999),
.ZN(net5002)
);

INV_X2 c4763(
.A(net2919),
.ZN(net5003)
);

INV_X8 c4764(
.A(net9656),
.ZN(net5004)
);

INV_X16 c4765(
.A(net10013),
.ZN(net5005)
);

OR3_X4 c4766(
.A1(net4983),
.A2(net4942),
.A3(net5003),
.ZN(net5006)
);

INV_X32 c4767(
.A(net5003),
.ZN(net5007)
);

NOR2_X2 c4768(
.A1(net5007),
.A2(net4999),
.ZN(net5008)
);

AND3_X2 c4769(
.A1(net4992),
.A2(net4991),
.A3(net4838),
.ZN(net5009)
);

SDFF_X2 c4770(
.D(net3943),
.SE(net4994),
.SI(net4059),
.CK(clk),
.Q(net5011),
.QN(net5010)
);

XOR2_X2 c4771(
.A(net4067),
.B(net10904),
.Z(net5012)
);

OAI221_X1 c4772(
.A(net4912),
.B1(net4991),
.B2(net3913),
.C1(net4966),
.C2(net4993),
.ZN(net5013)
);

XNOR2_X1 c4773(
.A(net5005),
.B(net4905),
.ZN(net5014)
);

OR2_X4 c4774(
.A1(net4996),
.A2(net4969),
.ZN(net5015)
);

INV_X4 c4775(
.A(net10344),
.ZN(net5016)
);

OR2_X1 c4776(
.A1(net5000),
.A2(net5003),
.ZN(net5017)
);

NOR3_X1 c4777(
.A1(net4869),
.A2(net4047),
.A3(net4990),
.ZN(net5018)
);

INV_X1 c4778(
.A(net4084),
.ZN(net5019)
);

XNOR2_X2 c4779(
.A(net5001),
.B(net4993),
.ZN(net5020)
);

OR3_X2 c4780(
.A1(net5008),
.A2(net4062),
.A3(net4895),
.ZN(net5021)
);

AND2_X4 c4781(
.A1(net4059),
.A2(net4908),
.ZN(net5022)
);

AND2_X1 c4782(
.A1(net4998),
.A2(net4062),
.ZN(net5023)
);

INV_X2 c4783(
.A(net9751),
.ZN(net5024)
);

DFFRS_X1 c4784(
.D(net5008),
.RN(net3072),
.SN(net10419),
.CK(clk),
.Q(net5026),
.QN(net5025)
);

INV_X8 c4785(
.A(net5023),
.ZN(net5027)
);

INV_X16 c4786(
.A(net5017),
.ZN(net5028)
);

OAI221_X4 c4787(
.A(net5028),
.B1(net4993),
.B2(net5008),
.C1(net5003),
.C2(net4080),
.ZN(net5029)
);

INV_X32 c4788(
.A(net9750),
.ZN(net5030)
);

OAI21_X2 c4789(
.A(net5018),
.B1(net4888),
.B2(net5010),
.ZN(net5031)
);

OAI221_X2 c4790(
.A(net4993),
.B1(net3117),
.B2(net4986),
.C1(net3052),
.C2(net4990),
.ZN(net5032)
);

INV_X4 c4791(
.A(net3072),
.ZN(net5033)
);

DFFRS_X2 c4792(
.D(net4894),
.RN(net5025),
.SN(net5027),
.CK(clk),
.Q(net5035),
.QN(net5034)
);

INV_X1 c4793(
.A(net4987),
.ZN(net5036)
);

INV_X2 c4794(
.A(net5030),
.ZN(net5037)
);

INV_X8 c4795(
.A(net4976),
.ZN(net5038)
);

INV_X16 c4796(
.A(net9963),
.ZN(net5039)
);

INV_X32 c4797(
.A(net5039),
.ZN(net5040)
);

OAI21_X1 c4798(
.A(net3919),
.B1(net4973),
.B2(net5014),
.ZN(net5041)
);

NAND2_X1 c4799(
.A1(net5037),
.A2(net4990),
.ZN(net5042)
);

INV_X4 c4800(
.A(net9699),
.ZN(net5043)
);

INV_X1 c4801(
.A(net10939),
.ZN(net5044)
);

SDFF_X1 c4802(
.D(net5042),
.SE(net5027),
.SI(net5043),
.CK(clk),
.Q(net5046),
.QN(net5045)
);

NAND2_X2 c4803(
.A1(net5038),
.A2(net5043),
.ZN(net5047)
);

NAND2_X4 c4804(
.A1(net5041),
.A2(net4985),
.ZN(net5048)
);

AOI21_X2 c4805(
.A(net4979),
.B1(net4064),
.B2(net5040),
.ZN(net5049)
);

INV_X2 c4806(
.A(net10335),
.ZN(net5050)
);

AOI21_X1 c4807(
.A(net4988),
.B1(net5037),
.B2(net10660),
.ZN(net5051)
);

AOI21_X4 c4808(
.A(net5051),
.B1(net5003),
.B2(net4800),
.ZN(net5052)
);

AND2_X2 c4809(
.A1(net4084),
.A2(net10899),
.ZN(net5053)
);

INV_X8 c4810(
.A(net9873),
.ZN(net5054)
);

AND3_X1 c4811(
.A1(net4797),
.A2(net5053),
.A3(net10745),
.ZN(net5055)
);

INV_X16 c4812(
.A(net10938),
.ZN(net5056)
);

NAND3_X1 c4813(
.A1(net5056),
.A2(net5026),
.A3(net5042),
.ZN(net5057)
);

INV_X32 c4814(
.A(net10997),
.ZN(net5058)
);

XOR2_X1 c4815(
.A(net4133),
.B(net5016),
.Z(net5059)
);

NOR2_X1 c4816(
.A1(net4036),
.A2(net3153),
.ZN(net5060)
);

INV_X4 c4817(
.A(net4047),
.ZN(net5061)
);

OR2_X2 c4818(
.A1(net4938),
.A2(net1270),
.ZN(net5062)
);

NOR2_X4 c4819(
.A1(net4996),
.A2(net5058),
.ZN(net5063)
);

NOR2_X2 c4820(
.A1(net4148),
.A2(net4098),
.ZN(net5064)
);

XOR2_X2 c4821(
.A(net3935),
.B(net3101),
.Z(net5065)
);

INV_X1 c4822(
.A(net4131),
.ZN(net5066)
);

XNOR2_X1 c4823(
.A(net4895),
.B(net4934),
.ZN(net5067)
);

SDFF_X2 c4824(
.D(net4971),
.SE(net3211),
.SI(net3134),
.CK(clk),
.Q(net5069),
.QN(net5068)
);

INV_X2 c4825(
.A(net4062),
.ZN(net5070)
);

INV_X8 c4826(
.A(net10907),
.ZN(net5071)
);

OR2_X4 c4827(
.A1(net5066),
.A2(net10907),
.ZN(net5072)
);

OR2_X1 c4828(
.A1(net4001),
.A2(net4917),
.ZN(net5073)
);

INV_X16 c4829(
.A(net4058),
.ZN(net5074)
);

XNOR2_X2 c4830(
.A(net4087),
.B(net3857),
.ZN(net5075)
);

AND2_X4 c4831(
.A1(net5066),
.A2(net3100),
.ZN(net5076)
);

AND2_X1 c4832(
.A1(net3080),
.A2(net4939),
.ZN(net5077)
);

INV_X32 c4833(
.A(net4906),
.ZN(net5078)
);

NAND2_X1 c4834(
.A1(net251),
.A2(net5024),
.ZN(net5079)
);

NAND2_X2 c4835(
.A1(net4140),
.A2(net3060),
.ZN(net5080)
);

NAND2_X4 c4836(
.A1(net5058),
.A2(net4938),
.ZN(net5081)
);

AND2_X2 c4837(
.A1(net5080),
.A2(net4999),
.ZN(net5082)
);

XOR2_X1 c4838(
.A(net5024),
.B(net2959),
.Z(net5083)
);

NOR3_X4 c4839(
.A1(net5065),
.A2(net4080),
.A3(net5077),
.ZN(net5084)
);

INV_X4 c4840(
.A(net5044),
.ZN(net5085)
);

NOR2_X1 c4841(
.A1(net5081),
.A2(net5077),
.ZN(net5086)
);

OR2_X2 c4842(
.A1(net5067),
.A2(net3925),
.ZN(net5087)
);

NOR2_X4 c4843(
.A1(net5086),
.A2(net4031),
.ZN(net5088)
);

NOR2_X2 c4844(
.A1(net3100),
.A2(net3935),
.ZN(net5089)
);

XOR2_X2 c4845(
.A(net3913),
.B(net4986),
.Z(net5090)
);

XNOR2_X1 c4846(
.A(net5082),
.B(net2110),
.ZN(net5091)
);

NOR3_X2 c4847(
.A1(net5060),
.A2(net4134),
.A3(net5077),
.ZN(net5092)
);

INV_X1 c4848(
.A(net10359),
.ZN(net5093)
);

AND3_X4 c4849(
.A1(net3211),
.A2(net5082),
.A3(net3200),
.ZN(net5094)
);

NAND3_X2 c4850(
.A1(net5011),
.A2(net4153),
.A3(net5077),
.ZN(net5095)
);

OR2_X4 c4851(
.A1(net5071),
.A2(net5043),
.ZN(net5096)
);

OR3_X1 c4852(
.A1(net5083),
.A2(net4832),
.A3(net5059),
.ZN(net5097)
);

INV_X2 c4853(
.A(net10978),
.ZN(net5098)
);

OR2_X1 c4854(
.A1(net5060),
.A2(net10933),
.ZN(net5099)
);

INV_X8 c4855(
.A(net10916),
.ZN(net5100)
);

MUX2_X1 c4856(
.A(net5096),
.B(net5093),
.S(net4109),
.Z(net5101)
);

OAI21_X4 c4857(
.A(net4161),
.B1(net5097),
.B2(net4996),
.ZN(net5102)
);

XNOR2_X2 c4858(
.A(net4153),
.B(net5076),
.ZN(net5103)
);

AND2_X4 c4859(
.A1(net5093),
.A2(net10845),
.ZN(net5104)
);

AND2_X1 c4860(
.A1(net5103),
.A2(net5089),
.ZN(net5105)
);

NAND2_X1 c4861(
.A1(net4051),
.A2(net5040),
.ZN(net5106)
);

NAND2_X2 c4862(
.A1(net3860),
.A2(net5096),
.ZN(net5107)
);

NAND2_X4 c4863(
.A1(net5024),
.A2(net11153),
.ZN(net5108)
);

INV_X16 c4864(
.A(net11006),
.ZN(net5109)
);

INV_X32 c4865(
.A(net9651),
.ZN(net5110)
);

MUX2_X2 c4866(
.A(net5062),
.B(net5099),
.S(net5095),
.Z(net5111)
);

SDFFRS_X2 c4867(
.D(net5090),
.RN(net5011),
.SE(net4147),
.SI(net5077),
.SN(net5059),
.CK(clk),
.Q(net5113),
.QN(net5112)
);

INV_X4 c4868(
.A(net9852),
.ZN(net5114)
);

AND2_X2 c4869(
.A1(net4016),
.A2(net2121),
.ZN(net5115)
);

NAND3_X4 c4870(
.A1(net5109),
.A2(net5097),
.A3(net5044),
.ZN(net5116)
);

XOR2_X1 c4871(
.A(net4965),
.B(net5108),
.Z(net5117)
);

NOR2_X1 c4872(
.A1(net5078),
.A2(net5067),
.ZN(net5118)
);

OR2_X2 c4873(
.A1(net4939),
.A2(net5058),
.ZN(net5119)
);

NOR4_X1 c4874(
.A1(net5075),
.A2(net5108),
.A3(net5106),
.A4(net5107),
.ZN(net5120)
);

NOR2_X4 c4875(
.A1(net5096),
.A2(net5098),
.ZN(net5121)
);

OR3_X4 c4876(
.A1(net5119),
.A2(net5095),
.A3(net4148),
.ZN(net5122)
);

INV_X1 c4877(
.A(net10337),
.ZN(net5123)
);

NOR2_X2 c4878(
.A1(net5104),
.A2(net5076),
.ZN(net5124)
);

XOR2_X2 c4879(
.A(net5027),
.B(net5089),
.Z(net5125)
);

XNOR2_X1 c4880(
.A(net5067),
.B(net10951),
.ZN(net5126)
);

INV_X2 c4881(
.A(net9910),
.ZN(net5127)
);

AND3_X2 c4882(
.A1(net5098),
.A2(net4964),
.A3(net5126),
.ZN(net5128)
);

NOR3_X1 c4883(
.A1(net5085),
.A2(net5089),
.A3(net5118),
.ZN(net5129)
);

AOI211_X2 c4884(
.A(net5124),
.B(net3203),
.C1(net4095),
.C2(net5077),
.ZN(net5130)
);

OR2_X4 c4885(
.A1(net5106),
.A2(net5117),
.ZN(net5131)
);

OR3_X2 c4886(
.A1(net5073),
.A2(net5103),
.A3(net5070),
.ZN(net5132)
);

OR2_X1 c4887(
.A1(net5126),
.A2(net10700),
.ZN(net5133)
);

XNOR2_X2 c4888(
.A(net4988),
.B(net5096),
.ZN(net5134)
);

INV_X8 c4889(
.A(net9650),
.ZN(net5135)
);

OAI21_X2 c4890(
.A(net5100),
.B1(net5135),
.B2(net5128),
.ZN(net5136)
);

AOI22_X1 c4891(
.A1(net4127),
.A2(net5135),
.B1(net4134),
.B2(net11015),
.ZN(net5137)
);

AND4_X4 c4892(
.A1(net5134),
.A2(net5089),
.A3(net5066),
.A4(net4986),
.ZN(net5138)
);

NAND4_X1 c4893(
.A1(net5116),
.A2(net5070),
.A3(net4159),
.A4(net5024),
.ZN(net5139)
);

OAI21_X1 c4894(
.A(net5118),
.B1(net5123),
.B2(net11005),
.ZN(net5140)
);

AOI21_X2 c4895(
.A(net4986),
.B1(net4798),
.B2(net5128),
.ZN(net5141)
);

AOI21_X1 c4896(
.A(net5131),
.B1(net5134),
.B2(net5126),
.ZN(net5142)
);

INV_X16 c4897(
.A(net10569),
.ZN(net5143)
);

AND2_X4 c4898(
.A1(net4999),
.A2(net3278),
.ZN(net5144)
);

INV_X32 c4899(
.A(net9723),
.ZN(net5145)
);

INV_X4 c4900(
.A(net11189),
.ZN(net5146)
);

INV_X1 c4901(
.A(net9564),
.ZN(net5147)
);

AND2_X1 c4902(
.A1(net3299),
.A2(net4982),
.ZN(net5148)
);

INV_X2 c4903(
.A(net4172),
.ZN(net5149)
);

CLKGATETST_X8 c4904(
.E(net4220),
.SE(net5093),
.CK(clk),
.GCK(net5150)
);

DFFR_X1 c4905(
.D(net5129),
.RN(net4024),
.CK(clk),
.Q(net5152),
.QN(net5151)
);

INV_X8 c4906(
.A(net9791),
.ZN(net5153)
);

NAND2_X1 c4907(
.A1(net3857),
.A2(net11188),
.ZN(net5154)
);

INV_X16 c4908(
.A(net10907),
.ZN(net5155)
);

INV_X32 c4909(
.A(net4958),
.ZN(net5156)
);

NAND2_X2 c4910(
.A1(net3204),
.A2(net5115),
.ZN(net5157)
);

NAND2_X4 c4911(
.A1(net1297),
.A2(net4958),
.ZN(net5158)
);

INV_X4 c4912(
.A(net4982),
.ZN(net5159)
);

AND2_X2 c4913(
.A1(net5102),
.A2(net5097),
.ZN(net5160)
);

XOR2_X1 c4914(
.A(net5159),
.B(net2884),
.Z(net5161)
);

NOR2_X1 c4915(
.A1(net5121),
.A2(net4191),
.ZN(net5162)
);

DFFRS_X1 c4916(
.D(net5155),
.RN(net4220),
.SN(net4217),
.CK(clk),
.Q(net5164),
.QN(net5163)
);

OR2_X2 c4917(
.A1(net4095),
.A2(net5146),
.ZN(net5165)
);

NOR2_X4 c4918(
.A1(net4899),
.A2(net3228),
.ZN(net5166)
);

NOR2_X2 c4919(
.A1(net3228),
.A2(net5166),
.ZN(net5167)
);

XOR2_X2 c4920(
.A(net4191),
.B(net5155),
.Z(net5168)
);

XNOR2_X1 c4921(
.A(net3278),
.B(net251),
.ZN(net5169)
);

INV_X1 c4922(
.A(net10261),
.ZN(net5170)
);

OR2_X4 c4923(
.A1(net4217),
.A2(net5160),
.ZN(net5171)
);

OR2_X1 c4924(
.A1(net5087),
.A2(net5167),
.ZN(net5172)
);

XNOR2_X2 c4925(
.A(net5152),
.B(net5150),
.ZN(net5173)
);

INV_X2 c4926(
.A(net5173),
.ZN(net5174)
);

AND2_X4 c4927(
.A1(net5118),
.A2(net5155),
.ZN(net5175)
);

AND2_X1 c4928(
.A1(net3269),
.A2(net1927),
.ZN(net5176)
);

INV_X8 c4929(
.A(net3187),
.ZN(net5177)
);

NAND2_X1 c4930(
.A1(net4832),
.A2(net5064),
.ZN(net5178)
);

AOI21_X4 c4931(
.A(net4977),
.B1(net5153),
.B2(net5150),
.ZN(net5179)
);

INV_X16 c4932(
.A(net3060),
.ZN(net5180)
);

INV_X32 c4933(
.A(net10369),
.ZN(net5181)
);

INV_X4 c4934(
.A(net9934),
.ZN(net5182)
);

AND3_X1 c4935(
.A1(net5115),
.A2(net2261),
.A3(net5129),
.ZN(net5183)
);

NAND2_X2 c4936(
.A1(net2245),
.A2(net5151),
.ZN(net5184)
);

NAND2_X4 c4937(
.A1(net5150),
.A2(net5157),
.ZN(net5185)
);

INV_X1 c4938(
.A(net9564),
.ZN(net5186)
);

INV_X2 c4939(
.A(net10237),
.ZN(net5187)
);

DFFRS_X2 c4940(
.D(net5165),
.RN(net5186),
.SN(net5138),
.CK(clk),
.Q(net5189),
.QN(net5188)
);

NAND3_X1 c4941(
.A1(net5076),
.A2(net5168),
.A3(net5153),
.ZN(net5190)
);

INV_X8 c4942(
.A(net4175),
.ZN(net5191)
);

AND2_X2 c4943(
.A1(net5097),
.A2(net5174),
.ZN(net5192)
);

XOR2_X1 c4944(
.A(net5147),
.B(net5175),
.Z(net5193)
);

NOR2_X1 c4945(
.A1(net5186),
.A2(net5146),
.ZN(net5194)
);

OR2_X2 c4946(
.A1(net4209),
.A2(net5162),
.ZN(net5195)
);

INV_X16 c4947(
.A(net10979),
.ZN(net5196)
);

NOR2_X4 c4948(
.A1(net5193),
.A2(net1230),
.ZN(net5197)
);

NOR2_X2 c4949(
.A1(net5189),
.A2(net5167),
.ZN(net5198)
);

INV_X32 c4950(
.A(net10118),
.ZN(net5199)
);

AOI221_X4 c4951(
.A(net5180),
.B1(net5199),
.B2(net5187),
.C1(net5165),
.C2(net3209),
.ZN(net5200)
);

NOR3_X4 c4952(
.A1(net5170),
.A2(net5099),
.A3(net5182),
.ZN(net5201)
);

OAI222_X1 c4953(
.A1(net4196),
.A2(net3269),
.B1(net4134),
.B2(net4185),
.C1(net5160),
.C2(net5166),
.ZN(net5202)
);

NOR3_X2 c4954(
.A1(net5161),
.A2(net5168),
.A3(net2261),
.ZN(net5203)
);

XOR2_X2 c4955(
.A(net1230),
.B(net5198),
.Z(net5204)
);

XNOR2_X1 c4956(
.A(net5195),
.B(net5186),
.ZN(net5205)
);

OR2_X4 c4957(
.A1(net5198),
.A2(net10800),
.ZN(net5206)
);

OR2_X1 c4958(
.A1(net5184),
.A2(net5162),
.ZN(net5207)
);

AND3_X4 c4959(
.A1(net5187),
.A2(net4207),
.A3(net5199),
.ZN(net5208)
);

NAND3_X2 c4960(
.A1(net5192),
.A2(net3187),
.A3(net11190),
.ZN(net5209)
);

INV_X4 c4961(
.A(net10264),
.ZN(net5210)
);

XNOR2_X2 c4962(
.A(net5165),
.B(net10426),
.ZN(net5211)
);

OR4_X1 c4963(
.A1(net5200),
.A2(net3269),
.A3(net5210),
.A4(net4185),
.ZN(net5212)
);

OR3_X1 c4964(
.A1(net5204),
.A2(net5165),
.A3(net11132),
.ZN(net5213)
);

MUX2_X1 c4965(
.A(net5061),
.B(net5188),
.S(net11191),
.Z(net5214)
);

OAI21_X4 c4966(
.A(net5214),
.B1(net2261),
.B2(net10584),
.ZN(net5215)
);

AND2_X4 c4967(
.A1(net5196),
.A2(net5210),
.ZN(net5216)
);

MUX2_X2 c4968(
.A(net5191),
.B(net5189),
.S(net5165),
.Z(net5217)
);

AND2_X1 c4969(
.A1(net5153),
.A2(net11060),
.ZN(net5218)
);

INV_X1 c4970(
.A(net10291),
.ZN(net5219)
);

NAND2_X1 c4971(
.A1(net5198),
.A2(net5219),
.ZN(net5220)
);

SDFF_X1 c4972(
.D(net5138),
.SE(net5200),
.SI(net3248),
.CK(clk),
.Q(net5222),
.QN(net5221)
);

NAND3_X4 c4973(
.A1(net4205),
.A2(net5222),
.A3(net10426),
.ZN(net5223)
);

OAI222_X4 c4974(
.A1(net5199),
.A2(net2245),
.B1(net5221),
.B2(net5166),
.C1(net3925),
.C2(net11060),
.ZN(net5224)
);

OR3_X4 c4975(
.A1(net5222),
.A2(net5224),
.A3(net5220),
.ZN(net5225)
);

NAND2_X2 c4976(
.A1(net5169),
.A2(net3258),
.ZN(net5226)
);

AND3_X2 c4977(
.A1(net5218),
.A2(net5222),
.A3(net11132),
.ZN(net5227)
);

OAI222_X2 c4978(
.A1(net3258),
.A2(net5216),
.B1(net5221),
.B2(net5025),
.C1(net4217),
.C2(net11190),
.ZN(net5228)
);

NOR3_X1 c4979(
.A1(net5224),
.A2(net5223),
.A3(net4030),
.ZN(net5229)
);

INV_X2 c4980(
.A(net5226),
.ZN(net5230)
);

NAND2_X4 c4981(
.A1(net5194),
.A2(net5197),
.ZN(net5231)
);

INV_X8 c4982(
.A(net2295),
.ZN(net5232)
);

AND2_X2 c4983(
.A1(net5181),
.A2(net3376),
.ZN(net5233)
);

XOR2_X1 c4984(
.A(net4203),
.B(net4329),
.Z(net5234)
);

SDFF_X2 c4985(
.D(net4301),
.SE(net5233),
.SI(net5207),
.CK(clk),
.Q(net5236),
.QN(net5235)
);

NOR2_X1 c4986(
.A1(net5223),
.A2(net4279),
.ZN(net5237)
);

INV_X16 c4987(
.A(net5197),
.ZN(net5238)
);

INV_X32 c4988(
.A(net9630),
.ZN(net5239)
);

OR2_X2 c4989(
.A1(net4198),
.A2(net4272),
.ZN(net5240)
);

INV_X4 c4990(
.A(net9630),
.ZN(net5241)
);

OR3_X2 c4991(
.A1(net5232),
.A2(net4207),
.A3(net4185),
.ZN(net5242)
);

OAI21_X2 c4992(
.A(net5237),
.B1(net5216),
.B2(net4312),
.ZN(net5243)
);

INV_X1 c4993(
.A(net11045),
.ZN(net5244)
);

INV_X2 c4994(
.A(net9707),
.ZN(net5245)
);

NOR2_X4 c4995(
.A1(net5243),
.A2(net5128),
.ZN(net5246)
);

INV_X8 c4996(
.A(net1279),
.ZN(net5247)
);

OAI21_X1 c4997(
.A(net3376),
.B1(net5230),
.B2(net5228),
.ZN(net5248)
);

NOR2_X2 c4998(
.A1(net4214),
.A2(net1392),
.ZN(net5249)
);

XOR2_X2 c4999(
.A(net5234),
.B(net4336),
.Z(net5250)
);

XNOR2_X1 c5000(
.A(net5145),
.B(net5239),
.ZN(net5251)
);

INV_X16 c5001(
.A(net5247),
.ZN(net5252)
);

OR2_X4 c5002(
.A1(net4317),
.A2(net4279),
.ZN(net5253)
);

INV_X32 c5003(
.A(net9723),
.ZN(net5254)
);

INV_X4 c5004(
.A(net5252),
.ZN(net5255)
);

OR2_X1 c5005(
.A1(net4240),
.A2(net5220),
.ZN(net5256)
);

INV_X1 c5006(
.A(net10153),
.ZN(net5257)
);

INV_X2 c5007(
.A(net5254),
.ZN(net5258)
);

AOI21_X2 c5008(
.A(net4291),
.B1(net5252),
.B2(net11086),
.ZN(net5259)
);

XNOR2_X2 c5009(
.A(net5197),
.B(net11086),
.ZN(net5260)
);

AOI21_X1 c5010(
.A(net5230),
.B1(net5241),
.B2(net3376),
.ZN(net5261)
);

AOI21_X4 c5011(
.A(net5246),
.B1(net5245),
.B2(net4312),
.ZN(net5262)
);

AND2_X4 c5012(
.A1(net5016),
.A2(net4177),
.ZN(net5263)
);

DFFRS_X1 c5013(
.D(net4177),
.RN(net5223),
.SN(net5262),
.CK(clk),
.Q(net5265),
.QN(net5264)
);

INV_X8 c5014(
.A(net5093),
.ZN(net5266)
);

INV_X16 c5015(
.A(net4318),
.ZN(net5267)
);

AND2_X1 c5016(
.A1(net5092),
.A2(net5263),
.ZN(net5268)
);

NAND2_X1 c5017(
.A1(net3362),
.A2(net5182),
.ZN(net5269)
);

INV_X32 c5018(
.A(net9733),
.ZN(net5270)
);

NAND2_X2 c5019(
.A1(net5258),
.A2(net4203),
.ZN(net5271)
);

NAND2_X4 c5020(
.A1(net5255),
.A2(net5266),
.ZN(net5272)
);

INV_X4 c5021(
.A(net10231),
.ZN(net5273)
);

AND2_X2 c5022(
.A1(net5260),
.A2(net11066),
.ZN(net5274)
);

INV_X1 c5023(
.A(net10293),
.ZN(net5275)
);

AND3_X1 c5024(
.A1(net5267),
.A2(net5263),
.A3(net5272),
.ZN(net5276)
);

NAND3_X1 c5025(
.A1(net5257),
.A2(net4279),
.A3(net4205),
.ZN(net5277)
);

INV_X2 c5026(
.A(net10080),
.ZN(net5278)
);

INV_X8 c5027(
.A(net10258),
.ZN(net5279)
);

NOR3_X4 c5028(
.A1(net5272),
.A2(net5260),
.A3(net5223),
.ZN(net5280)
);

AOI221_X2 c5029(
.A(net5262),
.B1(net4284),
.B2(net5206),
.C1(net5241),
.C2(net5239),
.ZN(net5281)
);

NOR3_X2 c5030(
.A1(net5259),
.A2(net5263),
.A3(net4284),
.ZN(net5282)
);

XOR2_X1 c5031(
.A(net3357),
.B(net4312),
.Z(net5283)
);

DFFR_X2 c5032(
.D(net2376),
.RN(net3169),
.CK(clk),
.Q(net5285),
.QN(net5284)
);

INV_X16 c5033(
.A(net11045),
.ZN(net5286)
);

NOR2_X1 c5034(
.A1(net5286),
.A2(net5133),
.ZN(net5287)
);

AND3_X4 c5035(
.A1(net4280),
.A2(net5287),
.A3(net5093),
.ZN(net5288)
);

OR2_X2 c5036(
.A1(net5270),
.A2(net3357),
.ZN(net5289)
);

NOR2_X4 c5037(
.A1(net4340),
.A2(net5272),
.ZN(net5290)
);

NOR2_X2 c5038(
.A1(net5248),
.A2(net5185),
.ZN(net5291)
);

DFFS_X1 c5039(
.D(net5233),
.SN(net5243),
.CK(clk),
.Q(net5293),
.QN(net5292)
);

NAND3_X2 c5040(
.A1(net4205),
.A2(net4336),
.A3(net11004),
.ZN(net5294)
);

XOR2_X2 c5041(
.A(net4311),
.B(net5219),
.Z(net5295)
);

OR3_X1 c5042(
.A1(net5293),
.A2(net5242),
.A3(net10746),
.ZN(net5296)
);

XNOR2_X1 c5043(
.A(net5293),
.B(net4945),
.ZN(net5297)
);

OR2_X4 c5044(
.A1(net5287),
.A2(net465),
.ZN(net5298)
);

MUX2_X1 c5045(
.A(net5295),
.B(net5294),
.S(net5016),
.Z(net5299)
);

OR2_X1 c5046(
.A1(net5297),
.A2(net5285),
.ZN(net5300)
);

XNOR2_X2 c5047(
.A(net4345),
.B(net5285),
.ZN(net5301)
);

AND2_X4 c5048(
.A1(net5251),
.A2(net5297),
.ZN(net5302)
);

INV_X32 c5049(
.A(net10152),
.ZN(net5303)
);

INV_X4 c5050(
.A(net11130),
.ZN(net5304)
);

DFFRS_X2 c5051(
.D(net5298),
.RN(net5297),
.SN(net5269),
.CK(clk),
.Q(net5306),
.QN(net5305)
);

AOI221_X1 c5052(
.A(net5136),
.B1(net5305),
.B2(net2376),
.C1(net5279),
.C2(net5253),
.ZN(net5307)
);

OAI221_X1 c5053(
.A(net4184),
.B1(net5099),
.B2(net4303),
.C1(net5279),
.C2(net3209),
.ZN(net5308)
);

OAI21_X4 c5054(
.A(net5240),
.B1(net5272),
.B2(net5297),
.ZN(net5309)
);

AND2_X1 c5055(
.A1(net5275),
.A2(net5302),
.ZN(net5310)
);

OAI221_X4 c5056(
.A(net5299),
.B1(net5310),
.B2(net5307),
.C1(net5266),
.C2(net5279),
.ZN(net5311)
);

NAND2_X1 c5057(
.A1(net5244),
.A2(net10567),
.ZN(net5312)
);

MUX2_X2 c5058(
.A(net5312),
.B(net5310),
.S(net5279),
.Z(net5313)
);

NAND3_X4 c5059(
.A1(net5273),
.A2(net5313),
.A3(net5286),
.ZN(net5314)
);

AOI222_X1 c5060(
.A1(net5278),
.A2(net5314),
.B1(net5271),
.B2(net5292),
.C1(net5264),
.C2(net5284),
.ZN(net5315)
);

NAND2_X2 c5061(
.A1(net5313),
.A2(net5314),
.ZN(net5316)
);

AOI222_X4 c5062(
.A1(net5316),
.A2(net5313),
.B1(net5314),
.B2(net4273),
.C1(net5284),
.C2(net10679),
.ZN(net5317)
);

NAND2_X4 c5063(
.A1(net4272),
.A2(net4363),
.ZN(net5318)
);

AND2_X2 c5064(
.A1(net5265),
.A2(net11032),
.ZN(net5319)
);

INV_X1 c5065(
.A(net937),
.ZN(net5320)
);

INV_X2 c5066(
.A(net4841),
.ZN(net5321)
);

INV_X8 c5067(
.A(net2454),
.ZN(net5322)
);

XOR2_X1 c5068(
.A(net4419),
.B(net5300),
.Z(net5323)
);

INV_X16 c5069(
.A(net5063),
.ZN(net5324)
);

NOR2_X1 c5070(
.A1(net4185),
.A2(net4414),
.ZN(net5325)
);

INV_X32 c5071(
.A(net4207),
.ZN(net5326)
);

INV_X4 c5072(
.A(net4917),
.ZN(net5327)
);

INV_X1 c5073(
.A(net9684),
.ZN(net5328)
);

OR2_X2 c5074(
.A1(net5263),
.A2(net4414),
.ZN(net5329)
);

NOR2_X4 c5075(
.A1(net4382),
.A2(net4207),
.ZN(net5330)
);

INV_X2 c5076(
.A(net9684),
.ZN(net5331)
);

INV_X8 c5077(
.A(net4414),
.ZN(net5332)
);

INV_X16 c5078(
.A(net5146),
.ZN(net5333)
);

INV_X32 c5079(
.A(net11116),
.ZN(net5334)
);

INV_X4 c5080(
.A(net4347),
.ZN(net5335)
);

INV_X1 c5081(
.A(net5271),
.ZN(net5336)
);

INV_X2 c5082(
.A(net5306),
.ZN(net5337)
);

INV_X8 c5083(
.A(net3387),
.ZN(net5338)
);

OR3_X4 c5084(
.A1(net5332),
.A2(net548),
.A3(net5338),
.ZN(net5339)
);

INV_X16 c5085(
.A(net5318),
.ZN(net5340)
);

NOR2_X2 c5086(
.A1(net5300),
.A2(net4409),
.ZN(net5341)
);

INV_X32 c5087(
.A(net9702),
.ZN(net5342)
);

INV_X4 c5088(
.A(net4363),
.ZN(net5343)
);

INV_X1 c5089(
.A(net5178),
.ZN(net5344)
);

SDFF_X1 c5090(
.D(net5327),
.SE(net5277),
.SI(net5207),
.CK(clk),
.Q(net5346),
.QN(net5345)
);

INV_X2 c5091(
.A(net10814),
.ZN(net5347)
);

INV_X8 c5092(
.A(net5329),
.ZN(net5348)
);

INV_X16 c5093(
.A(net10056),
.ZN(net5349)
);

OAI221_X2 c5094(
.A(net5128),
.B1(net3397),
.B2(net5346),
.C1(net5099),
.C2(net5321),
.ZN(net5350)
);

INV_X32 c5095(
.A(net4384),
.ZN(net5351)
);

XOR2_X2 c5096(
.A(net4344),
.B(net5349),
.Z(net5352)
);

OAI22_X1 c5097(
.A1(net5348),
.A2(net5338),
.B1(net5263),
.B2(net2491),
.ZN(net5353)
);

XNOR2_X1 c5098(
.A(net4276),
.B(net4382),
.ZN(net5354)
);

SDFFS_X2 c5099(
.D(net3429),
.SE(net5306),
.SI(net4413),
.SN(net5321),
.CK(clk),
.Q(net5356),
.QN(net5355)
);

OR2_X4 c5100(
.A1(net5347),
.A2(net4384),
.ZN(net5357)
);

OR2_X1 c5101(
.A1(net5277),
.A2(net4360),
.ZN(net5358)
);

INV_X4 c5102(
.A(net9735),
.ZN(net5359)
);

AND3_X2 c5103(
.A1(net5342),
.A2(net4276),
.A3(net4207),
.ZN(net5360)
);

XNOR2_X2 c5104(
.A(net1471),
.B(net5334),
.ZN(net5361)
);

INV_X1 c5105(
.A(net5304),
.ZN(net5362)
);

DFFS_X2 c5106(
.D(net5362),
.SN(net2473),
.CK(clk),
.Q(net5364),
.QN(net5363)
);

AND2_X4 c5107(
.A1(net5341),
.A2(net5360),
.ZN(net5365)
);

AND2_X1 c5108(
.A1(net5330),
.A2(net4432),
.ZN(net5366)
);

NAND2_X1 c5109(
.A1(net4383),
.A2(net5366),
.ZN(net5367)
);

INV_X2 c5110(
.A(net10141),
.ZN(net5368)
);

NAND2_X2 c5111(
.A1(net5319),
.A2(net5279),
.ZN(net5369)
);

NOR3_X1 c5112(
.A1(net5350),
.A2(net5368),
.A3(net5264),
.ZN(net5370)
);

NAND2_X4 c5113(
.A1(net5301),
.A2(net4384),
.ZN(net5371)
);

INV_X8 c5114(
.A(net10303),
.ZN(net5372)
);

SDFFR_X1 c5115(
.D(net5360),
.RN(net5265),
.SE(net5366),
.SI(net5321),
.CK(clk),
.Q(net5374),
.QN(net5373)
);

AND2_X2 c5116(
.A1(net5370),
.A2(net5236),
.ZN(net5375)
);

XOR2_X1 c5117(
.A(net5343),
.B(net5354),
.Z(net5376)
);

NOR2_X1 c5118(
.A1(net5336),
.A2(net4298),
.ZN(net5377)
);

INV_X16 c5119(
.A(net10029),
.ZN(net5378)
);

OR2_X2 c5120(
.A1(net5372),
.A2(net5377),
.ZN(net5379)
);

INV_X32 c5121(
.A(net10430),
.ZN(net5380)
);

OR3_X2 c5122(
.A1(net3348),
.A2(net5368),
.A3(net5373),
.ZN(net5381)
);

CLKGATETST_X1 c5123(
.E(net5379),
.SE(net5366),
.CK(clk),
.GCK(net5382)
);

INV_X4 c5124(
.A(net5382),
.ZN(net5383)
);

INV_X1 c5125(
.A(net5374),
.ZN(net5384)
);

NOR2_X4 c5126(
.A1(net5368),
.A2(net4185),
.ZN(net5385)
);

NOR2_X2 c5127(
.A1(net5324),
.A2(net5235),
.ZN(net5386)
);

AND4_X2 c5128(
.A1(net5220),
.A2(net4276),
.A3(net5368),
.A4(net5305),
.ZN(net5387)
);

OAI21_X2 c5129(
.A(net5358),
.B1(net4203),
.B2(net5382),
.ZN(net5388)
);

XOR2_X2 c5130(
.A(net5388),
.B(net5380),
.Z(net5389)
);

AND4_X1 c5131(
.A1(net5108),
.A2(net2481),
.A3(net5378),
.A4(net5166),
.ZN(net5390)
);

XNOR2_X1 c5132(
.A(net5326),
.B(net5385),
.ZN(net5391)
);

INV_X2 c5133(
.A(net10273),
.ZN(net5392)
);

OAI21_X1 c5134(
.A(net4298),
.B1(net5388),
.B2(net5385),
.ZN(net5393)
);

OR2_X4 c5135(
.A1(net5392),
.A2(net5383),
.ZN(net5394)
);

SDFF_X2 c5136(
.D(net5391),
.SE(net5241),
.SI(net10429),
.CK(clk),
.Q(net5396),
.QN(net5395)
);

OR2_X1 c5137(
.A1(net5382),
.A2(net10757),
.ZN(net5397)
);

CLKGATETST_X2 c5138(
.E(net5393),
.SE(net5356),
.CK(clk),
.GCK(net5398)
);

CLKGATETST_X4 c5139(
.E(net5353),
.SE(net4430),
.CK(clk),
.GCK(net5399)
);

AOI21_X2 c5140(
.A(net5390),
.B1(net5398),
.B2(net4418),
.ZN(net5400)
);

INV_X8 c5141(
.A(net10300),
.ZN(net5401)
);

AOI21_X1 c5142(
.A(net5400),
.B1(net5396),
.B2(net4344),
.ZN(net5402)
);

XNOR2_X2 c5143(
.A(net5397),
.B(net5396),
.ZN(net5403)
);

INV_X16 c5144(
.A(net10942),
.ZN(net5404)
);

AND2_X4 c5145(
.A1(net5403),
.A2(net5404),
.ZN(net5405)
);

INV_X32 c5146(
.A(net5383),
.ZN(net5406)
);

INV_X4 c5147(
.A(net9622),
.ZN(net5407)
);

INV_X1 c5148(
.A(net5371),
.ZN(net5408)
);

INV_X2 c5149(
.A(net5338),
.ZN(net5409)
);

INV_X8 c5150(
.A(net10227),
.ZN(net5410)
);

AND2_X1 c5151(
.A1(net5369),
.A2(net5381),
.ZN(net5411)
);

NAND2_X1 c5152(
.A1(net4515),
.A2(net5339),
.ZN(net5412)
);

AOI21_X4 c5153(
.A(net2594),
.B1(net4420),
.B2(net4461),
.ZN(net5413)
);

INV_X16 c5154(
.A(net9622),
.ZN(net5414)
);

INV_X32 c5155(
.A(net4456),
.ZN(net5415)
);

NAND2_X2 c5156(
.A1(net4333),
.A2(net5333),
.ZN(net5416)
);

AND3_X1 c5157(
.A1(net5410),
.A2(net5241),
.A3(net5401),
.ZN(net5417)
);

INV_X4 c5158(
.A(net10970),
.ZN(net5418)
);

NAND2_X4 c5159(
.A1(net5415),
.A2(net5279),
.ZN(net5419)
);

INV_X1 c5160(
.A(net5207),
.ZN(net5420)
);

INV_X2 c5161(
.A(net9735),
.ZN(net5421)
);

AND2_X2 c5162(
.A1(net4518),
.A2(net5285),
.ZN(net5422)
);

INV_X8 c5163(
.A(net5416),
.ZN(net5423)
);

XOR2_X1 c5164(
.A(net5361),
.B(net4477),
.Z(net5424)
);

INV_X16 c5165(
.A(net10186),
.ZN(net5425)
);

INV_X32 c5166(
.A(net4409),
.ZN(net5426)
);

INV_X4 c5167(
.A(net5422),
.ZN(net5427)
);

INV_X1 c5168(
.A(net5418),
.ZN(net5428)
);

INV_X2 c5169(
.A(net3538),
.ZN(net5429)
);

INV_X8 c5170(
.A(net11004),
.ZN(net5430)
);

NOR2_X1 c5171(
.A1(net5409),
.A2(net4371),
.ZN(net5431)
);

OR2_X2 c5172(
.A1(net5430),
.A2(net10513),
.ZN(net5432)
);

INV_X16 c5173(
.A(net10025),
.ZN(net5433)
);

NAND3_X1 c5174(
.A1(net5352),
.A2(net5253),
.A3(net5431),
.ZN(net5434)
);

NOR2_X4 c5175(
.A1(net5426),
.A2(net3544),
.ZN(net5435)
);

NOR2_X2 c5176(
.A1(net5430),
.A2(net5241),
.ZN(net5436)
);

INV_X32 c5177(
.A(net3521),
.ZN(net5437)
);

XOR2_X2 c5178(
.A(net5421),
.B(net4395),
.Z(net5438)
);

DFFRS_X1 c5179(
.D(net5408),
.RN(net4471),
.SN(net5414),
.CK(clk),
.Q(net5440),
.QN(net5439)
);

XNOR2_X1 c5180(
.A(net5423),
.B(net5438),
.ZN(net5441)
);

OR2_X4 c5181(
.A1(net5424),
.A2(net5253),
.ZN(net5442)
);

OR2_X1 c5182(
.A1(net5441),
.A2(net5422),
.ZN(net5443)
);

XNOR2_X2 c5183(
.A(net4371),
.B(net5422),
.ZN(net5444)
);

AND2_X4 c5184(
.A1(net2592),
.A2(net5431),
.ZN(net5445)
);

AND2_X1 c5185(
.A1(net4160),
.A2(net5424),
.ZN(net5446)
);

NAND2_X1 c5186(
.A1(net5428),
.A2(net2546),
.ZN(net5447)
);

NAND2_X2 c5187(
.A1(net5417),
.A2(net5380),
.ZN(net5448)
);

NAND2_X4 c5188(
.A1(net5446),
.A2(net5439),
.ZN(net5449)
);

AND2_X2 c5189(
.A1(net5419),
.A2(net4441),
.ZN(net5450)
);

XOR2_X1 c5190(
.A(net5413),
.B(net5279),
.Z(net5451)
);

INV_X4 c5191(
.A(net9780),
.ZN(net5452)
);

INV_X1 c5192(
.A(net5279),
.ZN(net5453)
);

NOR2_X1 c5193(
.A1(net5404),
.A2(net5438),
.ZN(net5454)
);

NOR3_X4 c5194(
.A1(net5429),
.A2(net3548),
.A3(net3544),
.ZN(net5455)
);

INV_X2 c5195(
.A(net10278),
.ZN(net5456)
);

INV_X8 c5196(
.A(net11085),
.ZN(net5457)
);

INV_X16 c5197(
.A(net11102),
.ZN(net5458)
);

OR2_X2 c5198(
.A1(net5339),
.A2(net5444),
.ZN(net5459)
);

INV_X32 c5199(
.A(net4441),
.ZN(net5460)
);

NOR2_X4 c5200(
.A1(net5450),
.A2(net10408),
.ZN(net5461)
);

NOR2_X2 c5201(
.A1(net5458),
.A2(net5406),
.ZN(net5462)
);

XOR2_X2 c5202(
.A(net5462),
.B(net2593),
.Z(net5463)
);

NOR3_X2 c5203(
.A1(net5448),
.A2(net5381),
.A3(net5359),
.ZN(net5464)
);

XNOR2_X1 c5204(
.A(net1392),
.B(net5458),
.ZN(net5465)
);

INV_X4 c5205(
.A(net5241),
.ZN(net5466)
);

OR2_X4 c5206(
.A1(net4491),
.A2(net1542),
.ZN(net5467)
);

OR2_X1 c5207(
.A1(net5420),
.A2(net5430),
.ZN(net5468)
);

AOI22_X4 c5208(
.A1(net5199),
.A2(net5452),
.B1(net5112),
.B2(net5284),
.ZN(net5469)
);

XNOR2_X2 c5209(
.A(net5450),
.B(net5468),
.ZN(net5470)
);

INV_X1 c5210(
.A(net11083),
.ZN(net5471)
);

AND3_X4 c5211(
.A1(net5468),
.A2(net4425),
.A3(net4395),
.ZN(net5472)
);

NAND3_X2 c5212(
.A1(net5470),
.A2(net5456),
.A3(net5471),
.ZN(net5473)
);

AND2_X4 c5213(
.A1(net5472),
.A2(net5460),
.ZN(net5474)
);

AND2_X1 c5214(
.A1(net5457),
.A2(net5474),
.ZN(net5475)
);

NAND2_X1 c5215(
.A1(net5333),
.A2(net5468),
.ZN(net5476)
);

OR3_X1 c5216(
.A1(net4474),
.A2(net5437),
.A3(net3538),
.ZN(net5477)
);

NAND2_X2 c5217(
.A1(net5438),
.A2(net5415),
.ZN(net5478)
);

MUX2_X1 c5218(
.A(net5432),
.B(net5424),
.S(net10647),
.Z(net5479)
);

DFFRS_X2 c5219(
.D(net5479),
.RN(net5477),
.SN(net5476),
.CK(clk),
.Q(net5481),
.QN(net5480)
);

NAND2_X4 c5220(
.A1(net4098),
.A2(net5446),
.ZN(net5482)
);

OAI33_X1 c5221(
.A1(net5478),
.A2(net5456),
.A3(net5469),
.B1(net5438),
.B2(net4460),
.B3(net5471),
.ZN(net5483)
);

AND2_X2 c5222(
.A1(net5433),
.A2(net5471),
.ZN(net5484)
);

SDFFRS_X1 c5223(
.D(net5414),
.RN(net5435),
.SE(net5477),
.SI(net5474),
.SN(net5417),
.CK(clk),
.Q(net5486),
.QN(net5485)
);

XOR2_X1 c5224(
.A(net4420),
.B(net5479),
.Z(net5487)
);

SDFFRS_X2 c5225(
.D(net5452),
.RN(net5380),
.SE(net5479),
.SI(net5439),
.SN(net5474),
.CK(clk),
.Q(net5489),
.QN(net5488)
);

AOI221_X4 c5226(
.A(net5473),
.B1(net4441),
.B2(net5440),
.C1(net5471),
.C2(net5284),
.ZN(net5490)
);

SDFF_X1 c5227(
.D(net5487),
.SE(net5476),
.SI(net5486),
.CK(clk),
.Q(net5492),
.QN(net5491)
);

SDFF_X2 c5228(
.D(net5490),
.SE(net5454),
.SI(net5164),
.CK(clk),
.Q(net5494),
.QN(net5493)
);

NOR2_X1 c5229(
.A1(net4596),
.A2(net5435),
.ZN(net5495)
);

OR2_X2 c5230(
.A1(net4569),
.A2(net1114),
.ZN(net5496)
);

INV_X2 c5231(
.A(net10104),
.ZN(out25)
);

NOR2_X4 c5232(
.A1(net5434),
.A2(net2490),
.ZN(net5497)
);

INV_X8 c5233(
.A(net11073),
.ZN(net5498)
);

OAI21_X4 c5234(
.A(net3557),
.B1(net5442),
.B2(net5495),
.ZN(net5499)
);

INV_X16 c5235(
.A(net10903),
.ZN(net5500)
);

NOR2_X2 c5236(
.A1(net5484),
.A2(net5476),
.ZN(net5501)
);

XOR2_X2 c5237(
.A(net5498),
.B(net4544),
.Z(net5502)
);

XNOR2_X1 c5238(
.A(net3594),
.B(net11100),
.ZN(net5503)
);

OR2_X4 c5239(
.A1(net2492),
.A2(net5493),
.ZN(net5504)
);

OR2_X1 c5240(
.A1(net5500),
.A2(net5285),
.ZN(net5505)
);

XNOR2_X2 c5241(
.A(net4598),
.B(net5503),
.ZN(net5506)
);

INV_X32 c5242(
.A(net5445),
.ZN(net5507)
);

AND2_X4 c5243(
.A1(net4595),
.A2(net4569),
.ZN(net5508)
);

AND2_X1 c5244(
.A1(net4527),
.A2(net4551),
.ZN(net5509)
);

NAND2_X1 c5245(
.A1(net4461),
.A2(net10482),
.ZN(net5510)
);

NAND2_X2 c5246(
.A1(net4402),
.A2(net2492),
.ZN(net5511)
);

INV_X4 c5247(
.A(net4573),
.ZN(net5512)
);

NAND2_X4 c5248(
.A1(net5401),
.A2(net5512),
.ZN(net5513)
);

AND2_X2 c5249(
.A1(net4533),
.A2(net4499),
.ZN(net5514)
);

XOR2_X1 c5250(
.A(net708),
.B(net10748),
.Z(net5515)
);

NOR2_X1 c5251(
.A1(net5497),
.A2(net5471),
.ZN(net5516)
);

INV_X1 c5252(
.A(net5506),
.ZN(net5517)
);

OR2_X2 c5253(
.A1(net5435),
.A2(net3625),
.ZN(net5518)
);

NOR2_X4 c5254(
.A1(net5517),
.A2(net4499),
.ZN(net5519)
);

NOR2_X2 c5255(
.A1(net4577),
.A2(net3571),
.ZN(net5520)
);

INV_X2 c5256(
.A(net4205),
.ZN(net5521)
);

XOR2_X2 c5257(
.A(net4551),
.B(net10461),
.Z(net5522)
);

XNOR2_X1 c5258(
.A(net5436),
.B(net3617),
.ZN(net5523)
);

INV_X8 c5259(
.A(net4467),
.ZN(net5524)
);

OR2_X4 c5260(
.A1(net4603),
.A2(net5160),
.ZN(net5525)
);

INV_X16 c5261(
.A(net9870),
.ZN(net5526)
);

INV_X32 c5262(
.A(net11062),
.ZN(net5527)
);

OR2_X1 c5263(
.A1(net5467),
.A2(net3576),
.ZN(net5528)
);

INV_X4 c5264(
.A(net11133),
.ZN(net5529)
);

XNOR2_X2 c5265(
.A(net5501),
.B(net4273),
.ZN(net5530)
);

AND2_X4 c5266(
.A1(net4539),
.A2(net10481),
.ZN(net5531)
);

AND2_X1 c5267(
.A1(net5453),
.A2(net4577),
.ZN(net5532)
);

NAND2_X1 c5268(
.A1(net5521),
.A2(net4329),
.ZN(net5533)
);

NAND2_X2 c5269(
.A1(net5514),
.A2(net5531),
.ZN(net5534)
);

INV_X1 c5270(
.A(net11079),
.ZN(net5535)
);

NAND2_X4 c5271(
.A1(net5502),
.A2(net5496),
.ZN(net5536)
);

INV_X2 c5272(
.A(net10105),
.ZN(net5537)
);

INV_X8 c5273(
.A(net10266),
.ZN(net5538)
);

AND2_X2 c5274(
.A1(net4559),
.A2(net4479),
.ZN(net5539)
);

XOR2_X1 c5275(
.A(net5523),
.B(net5512),
.Z(net5540)
);

INV_X16 c5276(
.A(net9966),
.ZN(net5541)
);

MUX2_X2 c5277(
.A(net4506),
.B(net699),
.S(net4594),
.Z(net5542)
);

NOR2_X1 c5278(
.A1(net5540),
.A2(net5026),
.ZN(net5543)
);

CLKGATETST_X8 c5279(
.E(net4597),
.SE(net5525),
.CK(clk),
.GCK(net5544)
);

INV_X32 c5280(
.A(net5529),
.ZN(net5545)
);

INV_X4 c5281(
.A(net5536),
.ZN(net5546)
);

OR2_X2 c5282(
.A1(net5542),
.A2(net5544),
.ZN(net5547)
);

NOR2_X4 c5283(
.A1(net5522),
.A2(net4551),
.ZN(net5548)
);

NOR2_X2 c5284(
.A1(net5548),
.A2(net5492),
.ZN(net5549)
);

XOR2_X2 c5285(
.A(net5511),
.B(net5547),
.Z(net5550)
);

XNOR2_X1 c5286(
.A(net4539),
.B(net5538),
.ZN(net5551)
);

OR2_X4 c5287(
.A1(net2490),
.A2(net5351),
.ZN(net5552)
);

OR2_X1 c5288(
.A1(net4582),
.A2(net5544),
.ZN(net5553)
);

XNOR2_X2 c5289(
.A(net5546),
.B(net5492),
.ZN(net5554)
);

NAND3_X4 c5290(
.A1(net5532),
.A2(net5549),
.A3(net5544),
.ZN(net5555)
);

AND2_X4 c5291(
.A1(net5547),
.A2(net5555),
.ZN(net5556)
);

AND2_X1 c5292(
.A1(net4432),
.A2(net5435),
.ZN(net5557)
);

INV_X1 c5293(
.A(net11058),
.ZN(net5558)
);

NAND2_X1 c5294(
.A1(net5545),
.A2(net5386),
.ZN(net5559)
);

AOI222_X2 c5295(
.A1(net5496),
.A2(net5559),
.B1(net4550),
.B2(net5509),
.C1(net5488),
.C2(net10944),
.ZN(net5560)
);

NAND2_X2 c5296(
.A1(net5552),
.A2(net5551),
.ZN(net5561)
);

INV_X2 c5297(
.A(net10043),
.ZN(net5562)
);

OR3_X4 c5298(
.A1(net5560),
.A2(net5524),
.A3(net4031),
.ZN(net5563)
);

OAI222_X1 c5299(
.A1(net3561),
.A2(net5559),
.B1(net5560),
.B2(out25),
.C1(net5544),
.C2(net4544),
.ZN(net5564)
);

AND3_X2 c5300(
.A1(net5558),
.A2(net5172),
.A3(net5553),
.ZN(net5565)
);

INV_X8 c5301(
.A(net11073),
.ZN(net5566)
);

NOR3_X1 c5302(
.A1(net5508),
.A2(net5563),
.A3(net5566),
.ZN(net5567)
);

DFFRS_X1 c5303(
.D(net5550),
.RN(net5547),
.SN(net5566),
.CK(clk),
.Q(net5569),
.QN(net5568)
);

AOI221_X2 c5304(
.A(net5026),
.B1(net5559),
.B2(net5562),
.C1(net5544),
.C2(out25),
.ZN(net5570)
);

OAI222_X4 c5305(
.A1(net5526),
.A2(net5565),
.B1(net5566),
.B2(net4432),
.C1(net5345),
.C2(net10944),
.ZN(net5571)
);

NAND2_X4 c5306(
.A1(net5527),
.A2(net5566),
.ZN(net5572)
);

OAI222_X2 c5307(
.A1(net5572),
.A2(net4471),
.B1(net5509),
.B2(net4460),
.C1(net5544),
.C2(net10587),
.ZN(net5573)
);

OR3_X2 c5308(
.A1(net5359),
.A2(net5567),
.A3(net11029),
.ZN(net5574)
);

AOI221_X1 c5309(
.A(net5570),
.B1(net5560),
.B2(net4569),
.C1(net5566),
.C2(net4528),
.ZN(net5575)
);

OAI21_X2 c5310(
.A(net5573),
.B1(net5574),
.B2(net5541),
.ZN(net5576)
);

DFFRS_X2 c5311(
.D(net5576),
.RN(net5566),
.SN(net5445),
.CK(clk),
.Q(net5578),
.QN(net5577)
);

AND2_X2 c5312(
.A1(net4550),
.A2(net3672),
.ZN(net5579)
);

OAI221_X1 c5313(
.A(net4615),
.B1(net4550),
.B2(net4616),
.C1(net5395),
.C2(net3691),
.ZN(net5580)
);

INV_X16 c5314(
.A(net10363),
.ZN(net5581)
);

XOR2_X1 c5315(
.A(net4675),
.B(net3690),
.Z(net5582)
);

INV_X32 c5316(
.A(net11043),
.ZN(net5583)
);

OAI21_X1 c5317(
.A(net5583),
.B1(net4600),
.B2(net5265),
.ZN(net5584)
);

NOR2_X1 c5318(
.A1(net5504),
.A2(net3698),
.ZN(net5585)
);

OR2_X2 c5319(
.A1(net4499),
.A2(net5582),
.ZN(net5586)
);

INV_X4 c5320(
.A(net9919),
.ZN(net5587)
);

INV_X1 c5321(
.A(net10942),
.ZN(net5588)
);

NOR2_X4 c5322(
.A1(net3727),
.A2(net3713),
.ZN(net5589)
);

NOR2_X2 c5323(
.A1(net4635),
.A2(net5512),
.ZN(net5590)
);

INV_X2 c5324(
.A(net10994),
.ZN(net5591)
);

XOR2_X2 c5325(
.A(net5365),
.B(net5582),
.Z(net5592)
);

XNOR2_X1 c5326(
.A(net3713),
.B(net5533),
.ZN(net5593)
);

OR2_X4 c5327(
.A1(net5535),
.A2(net5553),
.ZN(net5594)
);

OR2_X1 c5328(
.A1(net3447),
.A2(net5567),
.ZN(net5595)
);

XNOR2_X2 c5329(
.A(net3678),
.B(net828),
.ZN(net5596)
);

AND2_X4 c5330(
.A1(net5442),
.A2(net5594),
.ZN(net5597)
);

AND2_X1 c5331(
.A1(net5471),
.A2(net5588),
.ZN(net5598)
);

NAND2_X1 c5332(
.A1(net5567),
.A2(net4600),
.ZN(net5599)
);

NAND2_X2 c5333(
.A1(net5598),
.A2(net5583),
.ZN(net5600)
);

NAND2_X4 c5334(
.A1(net5496),
.A2(net5567),
.ZN(net5601)
);

INV_X8 c5335(
.A(net10960),
.ZN(net5602)
);

INV_X16 c5336(
.A(net9714),
.ZN(net5603)
);

AOI21_X2 c5337(
.A(net5351),
.B1(net2481),
.B2(net5489),
.ZN(net5604)
);

AND2_X2 c5338(
.A1(net465),
.A2(net5595),
.ZN(net5605)
);

AOI21_X1 c5339(
.A(net3690),
.B1(net5578),
.B2(net4650),
.ZN(net5606)
);

XOR2_X1 c5340(
.A(net3696),
.B(net3107),
.Z(net5607)
);

NOR2_X1 c5341(
.A1(net4612),
.A2(net5537),
.ZN(net5608)
);

INV_X32 c5342(
.A(net11119),
.ZN(net5609)
);

OR2_X2 c5343(
.A1(net3706),
.A2(net4273),
.ZN(net5610)
);

NOR2_X4 c5344(
.A1(net5554),
.A2(net4676),
.ZN(net5611)
);

AOI21_X4 c5345(
.A(net3718),
.B1(net3447),
.B2(net10388),
.ZN(net5612)
);

NOR2_X2 c5346(
.A1(net4681),
.A2(net4651),
.ZN(net5613)
);

XOR2_X2 c5347(
.A(net5595),
.B(net5613),
.Z(net5614)
);

AND3_X1 c5348(
.A1(net4551),
.A2(net5509),
.A3(net5533),
.ZN(net5615)
);

XNOR2_X1 c5349(
.A(net4594),
.B(net5590),
.ZN(net5616)
);

OR2_X4 c5350(
.A1(net5608),
.A2(net4612),
.ZN(net5617)
);

NAND3_X1 c5351(
.A1(net5582),
.A2(net5609),
.A3(net5172),
.ZN(net5618)
);

SDFF_X1 c5352(
.D(net1720),
.SE(net5597),
.SI(net3641),
.CK(clk),
.Q(net5620),
.QN(net5619)
);

OR2_X1 c5353(
.A1(net4623),
.A2(net5519),
.ZN(net5621)
);

XNOR2_X2 c5354(
.A(net5581),
.B(net5595),
.ZN(net5622)
);

AND2_X4 c5355(
.A1(net5603),
.A2(net5620),
.ZN(net5623)
);

INV_X4 c5356(
.A(net9689),
.ZN(net5624)
);

AND2_X1 c5357(
.A1(net5601),
.A2(net5609),
.ZN(net5625)
);

NAND2_X1 c5358(
.A1(net5617),
.A2(net10463),
.ZN(net5626)
);

NAND2_X2 c5359(
.A1(net5587),
.A2(net10538),
.ZN(net5627)
);

NAND2_X4 c5360(
.A1(net5610),
.A2(net5596),
.ZN(net5628)
);

SDFF_X2 c5361(
.D(net5346),
.SE(net5619),
.SI(net3696),
.CK(clk),
.Q(net5630),
.QN(net5629)
);

AND2_X2 c5362(
.A1(net5600),
.A2(net5628),
.ZN(net5631)
);

NOR3_X4 c5363(
.A1(net771),
.A2(net5596),
.A3(net5471),
.ZN(net5632)
);

XOR2_X1 c5364(
.A(net4273),
.B(net5629),
.Z(net5633)
);

DFFR_X1 c5365(
.D(net5495),
.RN(net5626),
.CK(clk),
.Q(net5635),
.QN(net5634)
);

INV_X1 c5366(
.A(net10055),
.ZN(net5636)
);

NOR2_X1 c5367(
.A1(net5585),
.A2(net5583),
.ZN(net5637)
);

OR2_X2 c5368(
.A1(net5625),
.A2(net5637),
.ZN(net5638)
);

NOR2_X4 c5369(
.A1(net5489),
.A2(net5637),
.ZN(net5639)
);

NOR3_X2 c5370(
.A1(net4604),
.A2(net5637),
.A3(net5635),
.ZN(net5640)
);

NOR2_X2 c5371(
.A1(net3448),
.A2(net5583),
.ZN(net5641)
);

DFFR_X2 c5372(
.D(net2481),
.RN(net5611),
.CK(clk),
.Q(net5643),
.QN(net5642)
);

INV_X2 c5373(
.A(net10142),
.ZN(net5644)
);

AND3_X4 c5374(
.A1(net4585),
.A2(net5614),
.A3(net5582),
.ZN(net5645)
);

DFFRS_X1 c5375(
.D(net5602),
.RN(net5644),
.SN(net5638),
.CK(clk),
.Q(net5647),
.QN(net5646)
);

INV_X8 c5376(
.A(net10180),
.ZN(net5648)
);

XOR2_X2 c5377(
.A(net5579),
.B(net5589),
.Z(net5649)
);

XNOR2_X1 c5378(
.A(net5406),
.B(net5639),
.ZN(net5650)
);

OR2_X4 c5379(
.A1(net5639),
.A2(net5628),
.ZN(net5651)
);

NAND3_X2 c5380(
.A1(net5537),
.A2(net5624),
.A3(net5650),
.ZN(net5652)
);

OR2_X1 c5381(
.A1(net5652),
.A2(net5412),
.ZN(net5653)
);

XNOR2_X2 c5382(
.A(net5386),
.B(net5631),
.ZN(net5654)
);

AND2_X4 c5383(
.A1(net5646),
.A2(net10387),
.ZN(net5655)
);

OAI221_X4 c5384(
.A(net5614),
.B1(net5655),
.B2(net4615),
.C1(net5582),
.C2(net5640),
.ZN(net5656)
);

SDFFRS_X1 c5385(
.D(net5640),
.RN(net5591),
.SE(net5655),
.SI(net5639),
.SN(net5632),
.CK(clk),
.Q(net5658),
.QN(net5657)
);

AND2_X1 c5386(
.A1(net5593),
.A2(net5599),
.ZN(net5659)
);

NAND2_X1 c5387(
.A1(net5648),
.A2(net10572),
.ZN(net5660)
);

NAND2_X2 c5388(
.A1(net5641),
.A2(net5615),
.ZN(net5661)
);

NAND2_X4 c5389(
.A1(net2696),
.A2(net5650),
.ZN(net5662)
);

OR3_X1 c5390(
.A1(net5609),
.A2(net5638),
.A3(net5657),
.ZN(net5663)
);

MUX2_X1 c5391(
.A(net5659),
.B(net5595),
.S(net10805),
.Z(net5664)
);

OAI221_X2 c5392(
.A(net4687),
.B1(net5651),
.B2(net4640),
.C1(net5657),
.C2(net5634),
.ZN(net5665)
);

AND2_X2 c5393(
.A1(net5553),
.A2(net5660),
.ZN(net5666)
);

INV_X16 c5394(
.A(net11043),
.ZN(net5667)
);

OAI21_X4 c5395(
.A(net1857),
.B1(net3768),
.B2(net5642),
.ZN(net5668)
);

XOR2_X1 c5396(
.A(net3651),
.B(net5395),
.Z(net5669)
);

NOR2_X1 c5397(
.A1(net4476),
.A2(net11169),
.ZN(net5670)
);

OR2_X2 c5398(
.A1(net5665),
.A2(net3737),
.ZN(net5671)
);

NOR2_X4 c5399(
.A1(net5643),
.A2(net4601),
.ZN(net5672)
);

INV_X32 c5400(
.A(net9648),
.ZN(net5673)
);

OAI22_X4 c5401(
.A1(net4753),
.A2(net4715),
.B1(net2808),
.B2(net4700),
.ZN(net5674)
);

AOI222_X1 c5402(
.A1(net3766),
.A2(net4693),
.B1(net4683),
.B2(net5577),
.C1(net4755),
.C2(net11182),
.ZN(net5675)
);

DFFS_X1 c5403(
.D(net5507),
.SN(net4702),
.CK(clk),
.Q(net5677),
.QN(net5676)
);

MUX2_X2 c5404(
.A(net5396),
.B(net4786),
.S(net4773),
.Z(net5678)
);

NAND3_X4 c5405(
.A1(net1816),
.A2(net3820),
.A3(net3672),
.ZN(net5679)
);

OR3_X4 c5406(
.A1(net4724),
.A2(net4786),
.A3(net11184),
.ZN(net5680)
);

DFFRS_X2 c5407(
.D(net4769),
.RN(net4712),
.SN(net5662),
.CK(clk),
.Q(net5682),
.QN(net5681)
);

INV_X4 c5408(
.A(net10166),
.ZN(net5683)
);

NOR2_X2 c5409(
.A1(net4699),
.A2(net3822),
.ZN(net5684)
);

XOR2_X2 c5410(
.A(net4786),
.B(net4724),
.Z(net5685)
);

XNOR2_X1 c5411(
.A(net2686),
.B(net4528),
.ZN(net5686)
);

OR2_X4 c5412(
.A1(net4601),
.A2(net10562),
.ZN(net5687)
);

OR2_X1 c5413(
.A1(net5684),
.A2(net5507),
.ZN(out16)
);

AND3_X2 c5414(
.A1(net5662),
.A2(net3812),
.A3(net10677),
.ZN(net5688)
);

NOR3_X1 c5415(
.A1(net2782),
.A2(net5662),
.A3(net5682),
.ZN(net5689)
);

OR3_X2 c5416(
.A1(net4683),
.A2(net5680),
.A3(net2674),
.ZN(net5690)
);

XNOR2_X2 c5417(
.A(net5669),
.B(net2814),
.ZN(net5691)
);

AND2_X4 c5418(
.A1(net4776),
.A2(net5647),
.ZN(net5692)
);

AND2_X1 c5419(
.A1(net4736),
.A2(net4748),
.ZN(net5693)
);

NAND2_X1 c5420(
.A1(net3786),
.A2(net11185),
.ZN(net5694)
);

OAI21_X2 c5421(
.A(net3812),
.B1(net3766),
.B2(net4754),
.ZN(net5695)
);

SDFF_X1 c5422(
.D(net3792),
.SE(net5665),
.SI(net3825),
.CK(clk),
.Q(net5697),
.QN(net5696)
);

NAND2_X2 c5423(
.A1(net4616),
.A2(net699),
.ZN(net5698)
);

NAND2_X4 c5424(
.A1(net5685),
.A2(net5679),
.ZN(net5699)
);

AND2_X2 c5425(
.A1(net5680),
.A2(net5509),
.ZN(net5700)
);

OAI21_X1 c5426(
.A(net5596),
.B1(net4649),
.B2(net4692),
.ZN(net5701)
);

AOI21_X2 c5427(
.A(net3785),
.B1(net5681),
.B2(net10648),
.ZN(net5702)
);

AOI21_X1 c5428(
.A(net5623),
.B1(net2712),
.B2(net4260),
.ZN(net5703)
);

XOR2_X1 c5429(
.A(net5679),
.B(net11185),
.Z(net5704)
);

NOR2_X1 c5430(
.A1(net5701),
.A2(net3794),
.ZN(net5705)
);

AOI21_X4 c5431(
.A(net5693),
.B1(net2781),
.B2(net3781),
.ZN(net5706)
);

DFFS_X2 c5432(
.D(net3746),
.SN(net5596),
.CK(clk),
.Q(net5708),
.QN(net5707)
);

AND3_X1 c5433(
.A1(net4762),
.A2(net2809),
.A3(net3781),
.ZN(net5709)
);

INV_X1 c5434(
.A(net9987),
.ZN(net5710)
);

OR2_X2 c5435(
.A1(net3821),
.A2(net11157),
.ZN(net5711)
);

NAND3_X1 c5436(
.A1(net1779),
.A2(net5704),
.A3(net10476),
.ZN(net5712)
);

SDFF_X2 c5437(
.D(net4754),
.SE(net5701),
.SI(net3797),
.CK(clk),
.Q(net5714),
.QN(net5713)
);

NOR3_X4 c5438(
.A1(net4649),
.A2(net2674),
.A3(net4601),
.ZN(net5715)
);

NOR2_X4 c5439(
.A1(net2558),
.A2(net5712),
.ZN(net5716)
);

NOR3_X2 c5440(
.A1(net5683),
.A2(net4717),
.A3(net11183),
.ZN(net5717)
);

AND3_X4 c5441(
.A1(net4716),
.A2(net4754),
.A3(net4712),
.ZN(net5718)
);

DFFRS_X1 c5442(
.D(net5618),
.RN(net5708),
.SN(net5701),
.CK(clk),
.Q(net5720),
.QN(net5719)
);

NOR2_X2 c5443(
.A1(net5706),
.A2(net5707),
.ZN(net5721)
);

NAND3_X2 c5444(
.A1(net5697),
.A2(net4699),
.A3(net5701),
.ZN(net5722)
);

XOR2_X2 c5445(
.A(net5716),
.B(net5643),
.Z(net5723)
);

DFFRS_X2 c5446(
.D(net5674),
.RN(net5715),
.SN(net3791),
.CK(clk),
.Q(net5725),
.QN(net5724)
);

INV_X2 c5447(
.A(net9647),
.ZN(net5726)
);

OR3_X1 c5448(
.A1(net5726),
.A2(net2781),
.A3(net10726),
.ZN(net5727)
);

XNOR2_X1 c5449(
.A(net3737),
.B(net4717),
.ZN(net5728)
);

OR2_X4 c5450(
.A1(net5702),
.A2(net2814),
.ZN(net5729)
);

MUX2_X1 c5451(
.A(net5700),
.B(net5701),
.S(net5696),
.Z(net5730)
);

INV_X8 c5452(
.A(net10089),
.ZN(net5731)
);

OR2_X1 c5453(
.A1(net5727),
.A2(net5700),
.ZN(net5732)
);

SDFF_X1 c5454(
.D(net5694),
.SE(net5732),
.SI(net4775),
.CK(clk),
.Q(net5734),
.QN(net5733)
);

OAI21_X4 c5455(
.A(net5729),
.B1(net5692),
.B2(net11169),
.ZN(net5735)
);

SDFF_X2 c5456(
.D(net5703),
.SE(net5715),
.SI(net5723),
.CK(clk),
.Q(net5737),
.QN(net5736)
);

DFFRS_X1 c5457(
.D(net5715),
.RN(net3758),
.SN(net5623),
.CK(clk),
.Q(net5739),
.QN(net5738)
);

MUX2_X2 c5458(
.A(net5734),
.B(net5713),
.S(net5692),
.Z(net5740)
);

NAND3_X4 c5459(
.A1(net3672),
.A2(net4755),
.A3(net5733),
.ZN(net5741)
);

OR3_X4 c5460(
.A1(net4702),
.A2(net5699),
.A3(net5679),
.ZN(net5742)
);

XNOR2_X2 c5461(
.A(net5737),
.B(net5733),
.ZN(net5743)
);

AND3_X2 c5462(
.A1(net5741),
.A2(net5647),
.A3(net5723),
.ZN(net5744)
);

DFFRS_X2 c5463(
.D(net4743),
.RN(net5735),
.SN(net5712),
.CK(clk),
.Q(net5746),
.QN(net5745)
);

INV_X16 c5464(
.A(net9965),
.ZN(net5747)
);

AND2_X4 c5465(
.A1(net4744),
.A2(net5730),
.ZN(net5748)
);

SDFF_X1 c5466(
.D(net5728),
.SE(net5736),
.SI(net5716),
.CK(clk),
.Q(net5750),
.QN(net5749)
);

NOR3_X1 c5467(
.A1(net4783),
.A2(net5644),
.A3(net5744),
.ZN(net5751)
);

OR3_X2 c5468(
.A1(net5721),
.A2(net5741),
.A3(net5723),
.ZN(net5752)
);

OAI21_X2 c5469(
.A(net5679),
.B1(net5734),
.B2(net5685),
.ZN(net5753)
);

SDFF_X2 c5470(
.D(net5740),
.SE(net4702),
.SI(net10695),
.CK(clk),
.Q(net5755),
.QN(net5754)
);

AOI22_X2 c5471(
.A1(net5711),
.A2(net5714),
.B1(net5754),
.B2(net11168),
.ZN(net5756)
);

AND2_X1 c5472(
.A1(net4746),
.A2(net5727),
.ZN(net5757)
);

OAI21_X1 c5473(
.A(net5691),
.B1(net5719),
.B2(net10795),
.ZN(net5758)
);

AOI222_X4 c5474(
.A1(net5665),
.A2(net5719),
.B1(out25),
.B2(net5681),
.C1(net10749),
.C2(net11157),
.ZN(net5759)
);

OAI33_X1 c5475(
.A1(net5757),
.A2(net5758),
.A3(net5755),
.B1(net5596),
.B2(net3640),
.B3(out25),
.ZN(net5760)
);

AOI21_X2 c5476(
.A(net5753),
.B1(net5756),
.B2(net11194),
.ZN(net5761)
);

AOI21_X1 c5477(
.A(net5726),
.B1(net5761),
.B2(net11195),
.ZN(net5762)
);

NAND2_X1 c5478(
.A1(net4854),
.A2(net2901),
.ZN(net5763)
);

INV_X32 c5479(
.A(net4824),
.ZN(net5764)
);

INV_X4 c5480(
.A(net4846),
.ZN(net5765)
);

INV_X1 c5481(
.A(net4824),
.ZN(net5766)
);

INV_X2 c5482(
.A(net4839),
.ZN(net5767)
);

INV_X8 c5483(
.A(net2901),
.ZN(net5768)
);

INV_X16 c5484(
.A(net4808),
.ZN(net5769)
);

INV_X32 c5485(
.A(net5765),
.ZN(net5770)
);

INV_X4 c5486(
.A(net3843),
.ZN(net5771)
);

CLKGATETST_X1 c5487(
.E(net4813),
.SE(net4871),
.CK(clk),
.GCK(net5772)
);

INV_X1 c5488(
.A(net4856),
.ZN(net5773)
);

INV_X2 c5489(
.A(net5770),
.ZN(net5774)
);

INV_X8 c5490(
.A(net4875),
.ZN(net5775)
);

INV_X16 c5491(
.A(net3874),
.ZN(net5776)
);

NAND2_X2 c5492(
.A1(net4807),
.A2(net5776),
.ZN(net5777)
);

NAND2_X4 c5493(
.A1(net4806),
.A2(net5776),
.ZN(net5778)
);

INV_X32 c5494(
.A(net4866),
.ZN(net5779)
);

AND2_X2 c5495(
.A1(net4845),
.A2(net2859),
.ZN(net5780)
);

INV_X4 c5496(
.A(net3913),
.ZN(net5781)
);

INV_X1 c5497(
.A(net976),
.ZN(net5782)
);

INV_X2 c5498(
.A(net9673),
.ZN(net5783)
);

INV_X8 c5499(
.A(net4866),
.ZN(net5784)
);

INV_X16 c5500(
.A(net9673),
.ZN(net5785)
);

INV_X32 c5501(
.A(net5773),
.ZN(net5786)
);

INV_X4 c5502(
.A(net9701),
.ZN(net5787)
);

XOR2_X1 c5503(
.A(net1004),
.B(net4808),
.Z(net5788)
);

CLKGATETST_X2 c5504(
.E(net5766),
.SE(net4864),
.CK(clk),
.GCK(net5789)
);

INV_X1 c5505(
.A(net5779),
.ZN(net5790)
);

INV_X2 c5506(
.A(net4849),
.ZN(net5791)
);

CLKGATETST_X4 c5507(
.E(net5770),
.SE(net3850),
.CK(clk),
.GCK(net5792)
);

AOI21_X4 c5508(
.A(net5773),
.B1(net4856),
.B2(net4805),
.ZN(net5793)
);

NOR2_X1 c5509(
.A1(net5785),
.A2(net5770),
.ZN(net5794)
);

INV_X8 c5510(
.A(net4882),
.ZN(net5795)
);

OR2_X2 c5511(
.A1(net5791),
.A2(net4865),
.ZN(net5796)
);

INV_X16 c5512(
.A(net10412),
.ZN(net5797)
);

INV_X32 c5513(
.A(net3898),
.ZN(net5798)
);

INV_X4 c5514(
.A(net5792),
.ZN(net5799)
);

AND3_X1 c5515(
.A1(net5798),
.A2(net5770),
.A3(net5786),
.ZN(net5800)
);

NOR2_X4 c5516(
.A1(net3843),
.A2(net4845),
.ZN(net5801)
);

INV_X1 c5517(
.A(net5796),
.ZN(net5802)
);

INV_X2 c5518(
.A(net5772),
.ZN(net5803)
);

INV_X8 c5519(
.A(net9857),
.ZN(net5804)
);

INV_X16 c5520(
.A(net5798),
.ZN(net5805)
);

INV_X32 c5521(
.A(net5777),
.ZN(net5806)
);

NOR2_X2 c5522(
.A1(net5802),
.A2(net5784),
.ZN(net5807)
);

INV_X4 c5523(
.A(net4818),
.ZN(net5808)
);

INV_X1 c5524(
.A(net5804),
.ZN(net5809)
);

INV_X2 c5525(
.A(net9739),
.ZN(net5810)
);

XOR2_X2 c5526(
.A(net5785),
.B(net5786),
.Z(net5811)
);

XNOR2_X1 c5527(
.A(net1978),
.B(net5793),
.ZN(net5812)
);

NAND3_X1 c5528(
.A1(net5799),
.A2(net5809),
.A3(net4798),
.ZN(net5813)
);

CLKGATETST_X8 c5529(
.E(net4813),
.SE(net5764),
.CK(clk),
.GCK(net5814)
);

INV_X8 c5530(
.A(net9760),
.ZN(net5815)
);

INV_X16 c5531(
.A(net5793),
.ZN(net5816)
);

INV_X32 c5532(
.A(net4839),
.ZN(net5817)
);

INV_X4 c5533(
.A(net5789),
.ZN(net5818)
);

INV_X1 c5534(
.A(net5787),
.ZN(net5819)
);

INV_X2 c5535(
.A(net5814),
.ZN(net5820)
);

OR2_X4 c5536(
.A1(net5811),
.A2(net5820),
.ZN(net5821)
);

DFFR_X1 c5537(
.D(net5816),
.RN(net2901),
.CK(clk),
.Q(net5823),
.QN(net5822)
);

INV_X8 c5538(
.A(net5782),
.ZN(net5824)
);

INV_X16 c5539(
.A(net5813),
.ZN(net5825)
);

INV_X32 c5540(
.A(net9808),
.ZN(net5826)
);

DFFRS_X1 c5541(
.D(net5812),
.RN(net5826),
.SN(net5795),
.CK(clk),
.Q(net5828),
.QN(net5827)
);

NOR3_X4 c5542(
.A1(net5809),
.A2(net5798),
.A3(net5826),
.ZN(net5829)
);

NOR3_X2 c5543(
.A1(net5800),
.A2(net5792),
.A3(net5799),
.ZN(net5830)
);

AND3_X4 c5544(
.A1(net5817),
.A2(net5829),
.A3(net5818),
.ZN(net5831)
);

DFFRS_X2 c5545(
.D(net5826),
.RN(net5789),
.SN(net5771),
.CK(clk),
.Q(net5833),
.QN(net5832)
);

DFFR_X2 c5546(
.D(net5768),
.RN(net5831),
.CK(clk),
.Q(net5835),
.QN(net5834)
);

OR2_X1 c5547(
.A1(net5828),
.A2(net5834),
.ZN(net5836)
);

NAND3_X2 c5548(
.A1(net5789),
.A2(net5818),
.A3(net5826),
.ZN(net5837)
);

OR3_X1 c5549(
.A1(net5829),
.A2(net5797),
.A3(net10421),
.ZN(net5838)
);

SDFFR_X2 c5550(
.D(net5831),
.RN(net5814),
.SE(net5763),
.SI(net5818),
.CK(clk),
.Q(net5840),
.QN(net5839)
);

MUX2_X1 c5551(
.A(net4814),
.B(net4881),
.S(net5834),
.Z(net5841)
);

XNOR2_X2 c5552(
.A(net5817),
.B(net10421),
.ZN(net5842)
);

OAI21_X4 c5553(
.A(net5819),
.B1(net5841),
.B2(net3912),
.ZN(net5843)
);

AOI222_X2 c5554(
.A1(net5803),
.A2(net5832),
.B1(net5814),
.B2(net5786),
.C1(net5808),
.C2(net4871),
.ZN(net5844)
);

MUX2_X2 c5555(
.A(net5810),
.B(net5839),
.S(net5837),
.Z(net5845)
);

SDFF_X1 c5556(
.D(net5841),
.SE(net3874),
.SI(net5808),
.CK(clk),
.Q(net5847),
.QN(net5846)
);

AND2_X4 c5557(
.A1(net5845),
.A2(net5796),
.ZN(net5848)
);

NAND3_X4 c5558(
.A1(net5825),
.A2(net5848),
.A3(net1004),
.ZN(net5849)
);

SDFFS_X1 c5559(
.D(net5847),
.SE(net5842),
.SI(net5845),
.SN(net5849),
.CK(clk),
.Q(net5851),
.QN(net5850)
);

NAND4_X4 c5560(
.A1(net5820),
.A2(net5846),
.A3(net5777),
.A4(net5848),
.ZN(net5852)
);

INV_X4 c5561(
.A(net4898),
.ZN(net5853)
);

INV_X1 c5562(
.A(net10807),
.ZN(net5854)
);

AND2_X1 c5563(
.A1(net5778),
.A2(net4890),
.ZN(net5855)
);

NAND2_X1 c5564(
.A1(net2049),
.A2(net4957),
.ZN(net5856)
);

INV_X2 c5565(
.A(net4859),
.ZN(net5857)
);

DFFS_X1 c5566(
.D(net4948),
.SN(net5764),
.CK(clk),
.Q(net5859),
.QN(net5858)
);

NAND2_X2 c5567(
.A1(net5764),
.A2(net10847),
.ZN(net5860)
);

OR3_X4 c5568(
.A1(net4951),
.A2(net5788),
.A3(net4904),
.ZN(net5861)
);

NAND2_X4 c5569(
.A1(net5780),
.A2(net4909),
.ZN(net5862)
);

AND2_X2 c5570(
.A1(net4833),
.A2(net5858),
.ZN(net5863)
);

XOR2_X1 c5571(
.A(net3925),
.B(net4838),
.Z(net5864)
);

NOR2_X1 c5572(
.A1(net5851),
.A2(net2049),
.ZN(net5865)
);

INV_X8 c5573(
.A(net9582),
.ZN(net5866)
);

OR2_X2 c5574(
.A1(net4929),
.A2(net5797),
.ZN(net5867)
);

NOR2_X4 c5575(
.A1(net3899),
.A2(net4872),
.ZN(net5868)
);

INV_X16 c5576(
.A(net4955),
.ZN(net5869)
);

NOR2_X2 c5577(
.A1(net3933),
.A2(net4951),
.ZN(net5870)
);

XOR2_X2 c5578(
.A(net4844),
.B(net5827),
.Z(net5871)
);

INV_X32 c5579(
.A(net10778),
.ZN(net5872)
);

INV_X4 c5580(
.A(net9582),
.ZN(net5873)
);

XNOR2_X1 c5581(
.A(net4844),
.B(net10437),
.ZN(net5874)
);

OR2_X4 c5582(
.A1(net5842),
.A2(net5778),
.ZN(net5875)
);

INV_X1 c5583(
.A(net5806),
.ZN(net5876)
);

AND3_X2 c5584(
.A1(net5875),
.A2(net3933),
.A3(net4885),
.ZN(net5877)
);

INV_X2 c5585(
.A(net10255),
.ZN(net5878)
);

INV_X8 c5586(
.A(net4904),
.ZN(net5879)
);

INV_X16 c5587(
.A(net10374),
.ZN(net5880)
);

NOR3_X1 c5588(
.A1(net5769),
.A2(net5764),
.A3(net1898),
.ZN(net5881)
);

INV_X32 c5589(
.A(net5833),
.ZN(net5882)
);

INV_X4 c5590(
.A(net930),
.ZN(net5883)
);

INV_X1 c5591(
.A(net9759),
.ZN(net5884)
);

INV_X2 c5592(
.A(net3007),
.ZN(net5885)
);

INV_X8 c5593(
.A(net10030),
.ZN(net5886)
);

DFFS_X2 c5594(
.D(net5878),
.SN(net2993),
.CK(clk),
.Q(net5888),
.QN(net5887)
);

OR2_X1 c5595(
.A1(net4844),
.A2(net2859),
.ZN(net5889)
);

XNOR2_X2 c5596(
.A(net4918),
.B(net4898),
.ZN(net5890)
);

AND2_X4 c5597(
.A1(net5863),
.A2(net5886),
.ZN(net5891)
);

AND2_X1 c5598(
.A1(net5888),
.A2(net5863),
.ZN(net5892)
);

INV_X16 c5599(
.A(net5854),
.ZN(net5893)
);

INV_X32 c5600(
.A(net9739),
.ZN(net5894)
);

INV_X4 c5601(
.A(net10376),
.ZN(net5895)
);

NAND2_X1 c5602(
.A1(net5883),
.A2(net10682),
.ZN(net5896)
);

NAND2_X2 c5603(
.A1(net5884),
.A2(net4930),
.ZN(net5897)
);

NAND2_X4 c5604(
.A1(net5883),
.A2(net5869),
.ZN(net5898)
);

AND2_X2 c5605(
.A1(net5885),
.A2(net3007),
.ZN(net5899)
);

INV_X1 c5606(
.A(net5882),
.ZN(net5900)
);

INV_X2 c5607(
.A(net9928),
.ZN(net5901)
);

XOR2_X1 c5608(
.A(net4873),
.B(net5879),
.Z(net5902)
);

SDFF_X2 c5609(
.D(net5887),
.SE(net5899),
.SI(net4936),
.CK(clk),
.Q(net5904),
.QN(net5903)
);

NOR2_X1 c5610(
.A1(net5797),
.A2(net4954),
.ZN(net5905)
);

INV_X8 c5611(
.A(net5805),
.ZN(net5906)
);

INV_X16 c5612(
.A(net5892),
.ZN(net5907)
);

OR3_X2 c5613(
.A1(net5876),
.A2(net5891),
.A3(net5864),
.ZN(net5908)
);

CLKGATETST_X1 c5614(
.E(net5868),
.SE(net5906),
.CK(clk),
.GCK(net5909)
);

OR2_X2 c5615(
.A1(net5905),
.A2(net4969),
.ZN(net5910)
);

INV_X32 c5616(
.A(net10807),
.ZN(net5911)
);

NOR2_X4 c5617(
.A1(net5910),
.A2(net5855),
.ZN(net5912)
);

OAI21_X2 c5618(
.A(net3981),
.B1(net5905),
.B2(net5904),
.ZN(net5913)
);

NOR2_X2 c5619(
.A1(net5912),
.A2(net5910),
.ZN(net5914)
);

OAI211_X2 c5620(
.A(net4909),
.B(net5876),
.C1(net5850),
.C2(net147),
.ZN(net5915)
);

OAI21_X1 c5621(
.A(net5893),
.B1(net5898),
.B2(net4889),
.ZN(net5916)
);

INV_X4 c5622(
.A(net9945),
.ZN(net5917)
);

XOR2_X2 c5623(
.A(net5895),
.B(net5886),
.Z(net5918)
);

XNOR2_X1 c5624(
.A(net5894),
.B(net5876),
.ZN(net5919)
);

AOI21_X2 c5625(
.A(net5855),
.B1(net5898),
.B2(net10555),
.ZN(net5920)
);

OR2_X4 c5626(
.A1(net5896),
.A2(net5898),
.ZN(net5921)
);

SDFFS_X2 c5627(
.D(net5914),
.SE(net5870),
.SI(net5904),
.SN(net5849),
.CK(clk),
.Q(net5923),
.QN(net5922)
);

OR2_X1 c5628(
.A1(net5916),
.A2(net4927),
.ZN(net5924)
);

INV_X1 c5629(
.A(net10778),
.ZN(net5925)
);

AOI21_X1 c5630(
.A(net5852),
.B1(net5910),
.B2(net10776),
.ZN(net5926)
);

XNOR2_X2 c5631(
.A(net5900),
.B(net3965),
.ZN(net5927)
);

AND2_X4 c5632(
.A1(net5906),
.A2(net4871),
.ZN(net5928)
);

OR4_X2 c5633(
.A1(net5920),
.A2(net5884),
.A3(net3007),
.A4(net5899),
.ZN(net5929)
);

AOI21_X4 c5634(
.A(net5925),
.B1(net5923),
.B2(net10712),
.ZN(net5930)
);

DFFRS_X1 c5635(
.D(net5764),
.RN(net5882),
.SN(net10682),
.CK(clk),
.Q(net5932),
.QN(net5931)
);

INV_X2 c5636(
.A(net10260),
.ZN(net5933)
);

DFFRS_X2 c5637(
.D(net5931),
.RN(net5862),
.SN(net10778),
.CK(clk),
.Q(net5935),
.QN(net5934)
);

AND3_X1 c5638(
.A1(net5927),
.A2(net5907),
.A3(net4910),
.ZN(net5936)
);

NAND3_X1 c5639(
.A1(net5932),
.A2(net4873),
.A3(net5806),
.ZN(net5937)
);

AND2_X1 c5640(
.A1(net5937),
.A2(net5925),
.ZN(net5938)
);

NOR3_X4 c5641(
.A1(net5918),
.A2(net5923),
.A3(net5937),
.ZN(net5939)
);

SDFFR_X1 c5642(
.D(net5930),
.RN(net5920),
.SE(net3850),
.SI(net5937),
.CK(clk),
.Q(net5941),
.QN(net5940)
);

OAI222_X1 c5643(
.A1(net5939),
.A2(net2993),
.B1(net5862),
.B2(net5899),
.C1(net5937),
.C2(net5783),
.ZN(net5942)
);

INV_X8 c5644(
.A(net4930),
.ZN(net5943)
);

INV_X16 c5645(
.A(net3990),
.ZN(net5944)
);

NAND2_X1 c5646(
.A1(net3848),
.A2(net3007),
.ZN(net5945)
);

NAND2_X2 c5647(
.A1(net4931),
.A2(net5865),
.ZN(net5946)
);

INV_X32 c5648(
.A(net9741),
.ZN(net5947)
);

INV_X4 c5649(
.A(net9646),
.ZN(net5948)
);

INV_X1 c5650(
.A(net11199),
.ZN(net5949)
);

INV_X2 c5651(
.A(net4817),
.ZN(net5950)
);

INV_X8 c5652(
.A(net3965),
.ZN(net5951)
);

NOR3_X2 c5653(
.A1(net4954),
.A2(net5949),
.A3(net5052),
.ZN(net5952)
);

AOI211_X1 c5654(
.A(net5052),
.B(net4930),
.C1(net5946),
.C2(net4080),
.ZN(net5953)
);

NAND2_X4 c5655(
.A1(net5901),
.A2(net5952),
.ZN(net5954)
);

AND2_X2 c5656(
.A1(net5909),
.A2(net4871),
.ZN(net5955)
);

INV_X16 c5657(
.A(net9645),
.ZN(net5956)
);

INV_X32 c5658(
.A(net5946),
.ZN(net5957)
);

XOR2_X1 c5659(
.A(net4082),
.B(net11199),
.Z(net5958)
);

INV_X4 c5660(
.A(net9717),
.ZN(net5959)
);

INV_X1 c5661(
.A(net4956),
.ZN(net5960)
);

NOR2_X1 c5662(
.A1(net5952),
.A2(net5956),
.ZN(net5961)
);

OR2_X2 c5663(
.A1(net5897),
.A2(net5827),
.ZN(net5962)
);

INV_X2 c5664(
.A(net5956),
.ZN(net5963)
);

INV_X8 c5665(
.A(net5865),
.ZN(net5964)
);

INV_X16 c5666(
.A(net9913),
.ZN(net5965)
);

NOR2_X4 c5667(
.A1(net3113),
.A2(net5040),
.ZN(net5966)
);

NAND4_X2 c5668(
.A1(net5964),
.A2(net5946),
.A3(net5952),
.A4(net5949),
.ZN(net5967)
);

OR4_X4 c5669(
.A1(net5946),
.A2(net5909),
.A3(net5866),
.A4(net5956),
.ZN(net5968)
);

NOR2_X2 c5670(
.A1(net5957),
.A2(net4923),
.ZN(net5969)
);

INV_X32 c5671(
.A(net10012),
.ZN(net5970)
);

XOR2_X2 c5672(
.A(net5960),
.B(net5949),
.Z(net5971)
);

XNOR2_X1 c5673(
.A(net4871),
.B(net3007),
.ZN(net5972)
);

INV_X4 c5674(
.A(net4892),
.ZN(net5973)
);

INV_X1 c5675(
.A(net10770),
.ZN(net5974)
);

OR2_X4 c5676(
.A1(net5954),
.A2(net5945),
.ZN(net5975)
);

OR2_X1 c5677(
.A1(net5971),
.A2(net3007),
.ZN(net5976)
);

AND3_X4 c5678(
.A1(net5004),
.A2(net4025),
.A3(net5886),
.ZN(net5977)
);

INV_X2 c5679(
.A(net5966),
.ZN(net5978)
);

INV_X8 c5680(
.A(net10694),
.ZN(net5979)
);

INV_X16 c5681(
.A(net10904),
.ZN(net5980)
);

INV_X32 c5682(
.A(net9917),
.ZN(net5981)
);

INV_X4 c5683(
.A(net5969),
.ZN(net5982)
);

XNOR2_X2 c5684(
.A(net5945),
.B(net5960),
.ZN(net5983)
);

INV_X1 c5685(
.A(net5772),
.ZN(net5984)
);

NAND3_X2 c5686(
.A1(net5052),
.A2(net5040),
.A3(net10568),
.ZN(net5985)
);

INV_X2 c5687(
.A(net9796),
.ZN(net5986)
);

INV_X8 c5688(
.A(net10076),
.ZN(net5987)
);

OR3_X1 c5689(
.A1(net5947),
.A2(net5986),
.A3(net4933),
.ZN(net5988)
);

INV_X16 c5690(
.A(net5890),
.ZN(net5989)
);

AND2_X4 c5691(
.A1(net5961),
.A2(net5870),
.ZN(net5990)
);

INV_X32 c5692(
.A(net10436),
.ZN(net5991)
);

AND2_X1 c5693(
.A1(net5978),
.A2(net5949),
.ZN(net5992)
);

INV_X4 c5694(
.A(net5984),
.ZN(net5993)
);

NAND2_X1 c5695(
.A1(net5907),
.A2(net5956),
.ZN(net5994)
);

MUX2_X1 c5696(
.A(net5980),
.B(net4990),
.S(net11198),
.Z(net5995)
);

OAI21_X4 c5697(
.A(net5986),
.B1(net5993),
.B2(net4985),
.ZN(net5996)
);

NAND2_X2 c5698(
.A1(net5974),
.A2(net4985),
.ZN(net5997)
);

NAND2_X4 c5699(
.A1(net5962),
.A2(net5943),
.ZN(net5998)
);

INV_X1 c5700(
.A(net5979),
.ZN(net5999)
);

AND2_X2 c5701(
.A1(net5987),
.A2(net5938),
.ZN(net6000)
);

INV_X2 c5702(
.A(net5054),
.ZN(net6001)
);

XOR2_X1 c5703(
.A(net5967),
.B(net6000),
.Z(net6002)
);

NOR2_X1 c5704(
.A1(net5997),
.A2(net5945),
.ZN(net6003)
);

OR2_X2 c5705(
.A1(net4923),
.A2(net6000),
.ZN(net6004)
);

MUX2_X2 c5706(
.A(net5993),
.B(net4080),
.S(net6000),
.Z(net6005)
);

INV_X8 c5707(
.A(net10869),
.ZN(net6006)
);

OAI22_X2 c5708(
.A1(net5022),
.A2(net5801),
.B1(net5865),
.B2(net5052),
.ZN(net6007)
);

NOR2_X4 c5709(
.A1(net5996),
.A2(net4908),
.ZN(net6008)
);

INV_X16 c5710(
.A(net9962),
.ZN(net6009)
);

INV_X32 c5711(
.A(net6009),
.ZN(net6010)
);

INV_X4 c5712(
.A(net9922),
.ZN(net6011)
);

NOR2_X2 c5713(
.A1(net6005),
.A2(net5033),
.ZN(net6012)
);

XOR2_X2 c5714(
.A(net5880),
.B(net5954),
.Z(net6013)
);

INV_X1 c5715(
.A(net11054),
.ZN(net6014)
);

NAND3_X4 c5716(
.A1(net5015),
.A2(net6013),
.A3(net6005),
.ZN(net6015)
);

XNOR2_X1 c5717(
.A(net6011),
.B(net6013),
.ZN(net6016)
);

SDFF_X1 c5718(
.D(net6002),
.SE(net5983),
.SI(net6014),
.CK(clk),
.Q(net6018),
.QN(net6017)
);

OR3_X4 c5719(
.A1(net5963),
.A2(net5965),
.A3(net5952),
.ZN(net6019)
);

SDFF_X2 c5720(
.D(net6008),
.SE(net5983),
.SI(net5944),
.CK(clk),
.Q(net6021),
.QN(net6020)
);

AND3_X2 c5721(
.A1(net6006),
.A2(net5952),
.A3(net5052),
.ZN(net6022)
);

OR2_X4 c5722(
.A1(net6014),
.A2(net11137),
.ZN(net6023)
);

OR2_X1 c5723(
.A1(net6022),
.A2(net10457),
.ZN(net6024)
);

XNOR2_X2 c5724(
.A(net5986),
.B(net10745),
.ZN(net6025)
);

NOR3_X1 c5725(
.A1(net6001),
.A2(net6002),
.A3(net6025),
.ZN(net6026)
);

DFFRS_X1 c5726(
.D(net6025),
.RN(net6026),
.SN(net6016),
.CK(clk),
.Q(net6028),
.QN(net6027)
);

OR3_X2 c5727(
.A1(net5819),
.A2(net4931),
.A3(net5995),
.ZN(net6029)
);

SDFFR_X2 c5728(
.D(net5060),
.RN(net5837),
.SE(net4147),
.SI(net3007),
.CK(clk),
.Q(net6031),
.QN(net6030)
);

INV_X2 c5729(
.A(net5970),
.ZN(net6032)
);

INV_X8 c5730(
.A(net10984),
.ZN(net6033)
);

INV_X16 c5731(
.A(net6000),
.ZN(net6034)
);

AND2_X4 c5732(
.A1(net5938),
.A2(net5110),
.ZN(net6035)
);

INV_X32 c5733(
.A(net5873),
.ZN(net6036)
);

INV_X4 c5734(
.A(net3210),
.ZN(net6037)
);

AND2_X1 c5735(
.A1(net1236),
.A2(net5107),
.ZN(net6038)
);

INV_X1 c5736(
.A(net2171),
.ZN(net6039)
);

INV_X2 c5737(
.A(net9642),
.ZN(net6040)
);

INV_X8 c5738(
.A(net9642),
.ZN(net6041)
);

NAND2_X1 c5739(
.A1(net5081),
.A2(net6023),
.ZN(net6042)
);

CLKGATETST_X2 c5740(
.E(net2229),
.SE(net278),
.CK(clk),
.GCK(net6043)
);

INV_X16 c5741(
.A(net9797),
.ZN(net6044)
);

INV_X32 c5742(
.A(net5117),
.ZN(net6045)
);

NAND2_X2 c5743(
.A1(net5828),
.A2(net5995),
.ZN(net6046)
);

INV_X4 c5744(
.A(net6032),
.ZN(net6047)
);

NAND2_X4 c5745(
.A1(net6039),
.A2(net5043),
.ZN(net6048)
);

AND2_X2 c5746(
.A1(net5140),
.A2(net3200),
.ZN(net6049)
);

INV_X1 c5747(
.A(net5126),
.ZN(net6050)
);

AOI221_X4 c5748(
.A(net6049),
.B1(net5123),
.B2(net2110),
.C1(net4099),
.C2(net6047),
.ZN(net6051)
);

INV_X2 c5749(
.A(net5043),
.ZN(net6052)
);

INV_X8 c5750(
.A(net10066),
.ZN(net6053)
);

XOR2_X1 c5751(
.A(net4109),
.B(net6031),
.Z(net6054)
);

INV_X16 c5752(
.A(net6053),
.ZN(net6055)
);

INV_X32 c5753(
.A(net6035),
.ZN(net6056)
);

INV_X4 c5754(
.A(net2195),
.ZN(net6057)
);

NOR2_X1 c5755(
.A1(net5991),
.A2(net3175),
.ZN(net6058)
);

OR2_X2 c5756(
.A1(net6033),
.A2(net4970),
.ZN(net6059)
);

NOR2_X4 c5757(
.A1(net6048),
.A2(net5060),
.ZN(net6060)
);

NOR2_X2 c5758(
.A1(net4908),
.A2(net6048),
.ZN(net6061)
);

XOR2_X2 c5759(
.A(net6044),
.B(net5135),
.Z(net6062)
);

XNOR2_X1 c5760(
.A(net6047),
.B(net5081),
.ZN(net6063)
);

INV_X1 c5761(
.A(net10324),
.ZN(net6064)
);

OR2_X4 c5762(
.A1(net1203),
.A2(net6064),
.ZN(net6065)
);

INV_X2 c5763(
.A(net4970),
.ZN(net6066)
);

INV_X8 c5764(
.A(net9721),
.ZN(net6067)
);

CLKGATETST_X4 c5765(
.E(net5095),
.SE(net4099),
.CK(clk),
.GCK(net6068)
);

OR2_X1 c5766(
.A1(net6055),
.A2(net6048),
.ZN(net6069)
);

INV_X16 c5767(
.A(net6067),
.ZN(net6070)
);

XNOR2_X2 c5768(
.A(net6042),
.B(net6069),
.ZN(net6071)
);

INV_X32 c5769(
.A(net6062),
.ZN(net6072)
);

INV_X4 c5770(
.A(net5077),
.ZN(net6073)
);

AND2_X4 c5771(
.A1(net6037),
.A2(net6068),
.ZN(net6074)
);

OAI21_X2 c5772(
.A(net6032),
.B1(net5992),
.B2(net6052),
.ZN(net6075)
);

OAI211_X4 c5773(
.A(net5137),
.B(net5869),
.C1(net6052),
.C2(net5922),
.ZN(net6076)
);

AND2_X1 c5774(
.A1(net5921),
.A2(net5994),
.ZN(net6077)
);

NAND2_X1 c5775(
.A1(net5788),
.A2(net6010),
.ZN(net6078)
);

INV_X1 c5776(
.A(net6078),
.ZN(net6079)
);

NAND2_X2 c5777(
.A1(net4168),
.A2(net5072),
.ZN(net6080)
);

INV_X2 c5778(
.A(net5059),
.ZN(net6081)
);

INV_X8 c5779(
.A(net6064),
.ZN(net6082)
);

NAND2_X4 c5780(
.A1(net4121),
.A2(net6045),
.ZN(net6083)
);

INV_X16 c5781(
.A(net6061),
.ZN(net6084)
);

AND2_X2 c5782(
.A1(net6045),
.A2(net6047),
.ZN(net6085)
);

INV_X32 c5783(
.A(net5120),
.ZN(net6086)
);

XOR2_X1 c5784(
.A(net6039),
.B(net5123),
.Z(net6087)
);

NOR2_X1 c5785(
.A1(net6075),
.A2(net3925),
.ZN(net6088)
);

INV_X4 c5786(
.A(net11072),
.ZN(net6089)
);

OAI211_X1 c5787(
.A(net6082),
.B(net6060),
.C1(net6030),
.C2(net6074),
.ZN(net6090)
);

OR2_X2 c5788(
.A1(net6066),
.A2(net3134),
.ZN(net6091)
);

INV_X1 c5789(
.A(net6072),
.ZN(net6092)
);

OAI21_X1 c5790(
.A(net6056),
.B1(net6087),
.B2(net6069),
.ZN(net6093)
);

NOR2_X4 c5791(
.A1(net6050),
.A2(net6060),
.ZN(net6094)
);

NOR2_X2 c5792(
.A1(net2166),
.A2(net6094),
.ZN(net6095)
);

XOR2_X2 c5793(
.A(net6083),
.B(net11126),
.Z(net6096)
);

XNOR2_X1 c5794(
.A(net6088),
.B(net6085),
.ZN(net6097)
);

INV_X2 c5795(
.A(net10149),
.ZN(net6098)
);

AOI21_X2 c5796(
.A(net5990),
.B1(net6068),
.B2(net6085),
.ZN(net6099)
);

AOI21_X1 c5797(
.A(net6094),
.B1(net6099),
.B2(net5140),
.ZN(net6100)
);

AOI21_X4 c5798(
.A(net4011),
.B1(net6084),
.B2(net6098),
.ZN(net6101)
);

OR2_X4 c5799(
.A1(net6090),
.A2(net6088),
.ZN(net6102)
);

OR2_X1 c5800(
.A1(net6034),
.A2(net5950),
.ZN(net6103)
);

NOR4_X4 c5801(
.A1(net6058),
.A2(net6093),
.A3(net6103),
.A4(net6096),
.ZN(net6104)
);

AOI221_X2 c5802(
.A(net5981),
.B1(net3134),
.B2(net5114),
.C1(net6028),
.C2(net6103),
.ZN(net6105)
);

AND3_X1 c5803(
.A1(net6059),
.A2(net6047),
.A3(net10909),
.ZN(net6106)
);

INV_X8 c5804(
.A(net10327),
.ZN(net6107)
);

NAND3_X1 c5805(
.A1(net5992),
.A2(net6107),
.A3(net11097),
.ZN(net6108)
);

XNOR2_X2 c5806(
.A(net6106),
.B(net6096),
.ZN(net6109)
);

AND2_X4 c5807(
.A1(net5034),
.A2(net11097),
.ZN(net6110)
);

AOI221_X1 c5808(
.A(net6080),
.B1(net6054),
.B2(net6103),
.C1(net3200),
.C2(net3134),
.ZN(net6111)
);

OAI221_X1 c5809(
.A(net6092),
.B1(net5043),
.B2(net6103),
.C1(net4134),
.C2(net10634),
.ZN(net6112)
);

AND2_X1 c5810(
.A1(net4216),
.A2(net5069),
.ZN(net6113)
);

NAND2_X1 c5811(
.A1(net5944),
.A2(net11121),
.ZN(net6114)
);

INV_X16 c5812(
.A(net4927),
.ZN(net6115)
);

NOR3_X4 c5813(
.A1(net5123),
.A2(net5211),
.A3(net6096),
.ZN(net6116)
);

NAND2_X2 c5814(
.A1(net5848),
.A2(net5205),
.ZN(net6117)
);

NAND2_X4 c5815(
.A1(net5853),
.A2(net5157),
.ZN(net6118)
);

INV_X32 c5816(
.A(net5968),
.ZN(net6119)
);

NOR3_X2 c5817(
.A1(net4942),
.A2(net6081),
.A3(net5994),
.ZN(net6120)
);

AND2_X2 c5818(
.A1(net6115),
.A2(net5175),
.ZN(net6121)
);

INV_X4 c5819(
.A(net11060),
.ZN(net6122)
);

INV_X1 c5820(
.A(net9540),
.ZN(net6123)
);

AND3_X4 c5821(
.A1(net5069),
.A2(net5072),
.A3(net5167),
.ZN(net6124)
);

INV_X2 c5822(
.A(net9539),
.ZN(net6125)
);

INV_X8 c5823(
.A(net11132),
.ZN(net6126)
);

XOR2_X1 c5824(
.A(net3200),
.B(net5886),
.Z(net6127)
);

INV_X16 c5825(
.A(net5205),
.ZN(net6128)
);

INV_X32 c5826(
.A(net6063),
.ZN(net6129)
);

NOR2_X1 c5827(
.A1(net6123),
.A2(net5160),
.ZN(net6130)
);

INV_X4 c5828(
.A(net6113),
.ZN(net6131)
);

INV_X1 c5829(
.A(net10102),
.ZN(net6132)
);

OR2_X2 c5830(
.A1(net5157),
.A2(net5968),
.ZN(net6133)
);

CLKGATETST_X8 c5831(
.E(net6065),
.SE(net5209),
.CK(clk),
.GCK(net6134)
);

INV_X2 c5832(
.A(net6040),
.ZN(net6135)
);

INV_X8 c5833(
.A(net10263),
.ZN(net6136)
);

INV_X16 c5834(
.A(net10845),
.ZN(net6137)
);

INV_X32 c5835(
.A(net6068),
.ZN(net6138)
);

INV_X4 c5836(
.A(net5064),
.ZN(net6139)
);

INV_X1 c5837(
.A(net10803),
.ZN(net6140)
);

NOR2_X4 c5838(
.A1(net5948),
.A2(net6134),
.ZN(net6141)
);

NOR2_X2 c5839(
.A1(net6114),
.A2(net6135),
.ZN(net6142)
);

XOR2_X2 c5840(
.A(net5870),
.B(net6129),
.Z(net6143)
);

INV_X2 c5841(
.A(net10320),
.ZN(net6144)
);

XNOR2_X1 c5842(
.A(net5168),
.B(net2110),
.ZN(net6145)
);

OR2_X4 c5843(
.A1(net6110),
.A2(net6142),
.ZN(net6146)
);

OR2_X1 c5844(
.A1(net6121),
.A2(net6146),
.ZN(net6147)
);

XNOR2_X2 c5845(
.A(net4093),
.B(net6036),
.ZN(net6148)
);

AND2_X4 c5846(
.A1(net5149),
.A2(net5848),
.ZN(net6149)
);

AND2_X1 c5847(
.A1(net5201),
.A2(net6074),
.ZN(net6150)
);

NAND2_X1 c5848(
.A1(net4251),
.A2(net3200),
.ZN(net6151)
);

NAND2_X2 c5849(
.A1(net3248),
.A2(net6113),
.ZN(net6152)
);

NAND2_X4 c5850(
.A1(net6077),
.A2(net5114),
.ZN(net6153)
);

AND2_X2 c5851(
.A1(net4134),
.A2(net5064),
.ZN(net6154)
);

DFFRS_X2 c5852(
.D(net6120),
.RN(net6137),
.SN(net6151),
.CK(clk),
.Q(net6156),
.QN(net6155)
);

XOR2_X1 c5853(
.A(net6148),
.B(net6063),
.Z(net6157)
);

NAND3_X2 c5854(
.A1(net6124),
.A2(net6119),
.A3(net6148),
.ZN(net6158)
);

NOR2_X1 c5855(
.A1(net6128),
.A2(net6148),
.ZN(net6159)
);

OR3_X1 c5856(
.A1(net6125),
.A2(net6152),
.A3(net6154),
.ZN(net6160)
);

OR2_X2 c5857(
.A1(net6127),
.A2(net6154),
.ZN(net6161)
);

INV_X8 c5858(
.A(net10179),
.ZN(net6162)
);

NOR2_X4 c5859(
.A1(net6126),
.A2(net6155),
.ZN(net6163)
);

INV_X16 c5860(
.A(net5950),
.ZN(net6164)
);

INV_X32 c5861(
.A(net6135),
.ZN(net6165)
);

NOR2_X2 c5862(
.A1(net6145),
.A2(net6144),
.ZN(net6166)
);

XOR2_X2 c5863(
.A(net4146),
.B(net6096),
.Z(net6167)
);

MUX2_X1 c5864(
.A(net6167),
.B(net5228),
.S(net6143),
.Z(net6168)
);

XNOR2_X1 c5865(
.A(net6140),
.B(net6115),
.ZN(net6169)
);

SDFF_X1 c5866(
.D(net6166),
.SE(net6133),
.SI(net6160),
.CK(clk),
.Q(net6171),
.QN(net6170)
);

OR2_X4 c5867(
.A1(net6165),
.A2(net6159),
.ZN(net6172)
);

OR2_X1 c5868(
.A1(net6142),
.A2(net4134),
.ZN(net6173)
);

XNOR2_X2 c5869(
.A(net6146),
.B(net6134),
.ZN(net6174)
);

OAI21_X4 c5870(
.A(net6109),
.B1(net6172),
.B2(net6140),
.ZN(net6175)
);

MUX2_X2 c5871(
.A(net6119),
.B(net6156),
.S(net5219),
.Z(net6176)
);

NAND3_X4 c5872(
.A1(net6151),
.A2(net6170),
.A3(net6161),
.ZN(net6177)
);

AND2_X4 c5873(
.A1(net6131),
.A2(net6169),
.ZN(net6178)
);

OR3_X4 c5874(
.A1(net6162),
.A2(net6147),
.A3(net6136),
.ZN(net6179)
);

AND3_X2 c5875(
.A1(net6161),
.A2(net6165),
.A3(net4222),
.ZN(net6180)
);

NOR3_X1 c5876(
.A1(net6169),
.A2(net6139),
.A3(net6179),
.ZN(net6181)
);

OR3_X2 c5877(
.A1(net6164),
.A2(net6156),
.A3(net6126),
.ZN(net6182)
);

OAI21_X2 c5878(
.A(net6041),
.B1(net6182),
.B2(net6165),
.ZN(net6183)
);

INV_X4 c5879(
.A(net11134),
.ZN(net6184)
);

OAI21_X1 c5880(
.A(net4096),
.B1(net6155),
.B2(net5219),
.ZN(net6185)
);

AOI21_X2 c5881(
.A(net6178),
.B1(net6079),
.B2(net10928),
.ZN(net6186)
);

AOI21_X1 c5882(
.A(net6154),
.B1(net6186),
.B2(net10845),
.ZN(net6187)
);

AND2_X1 c5883(
.A1(net6174),
.A2(net6152),
.ZN(net6188)
);

OAI221_X4 c5884(
.A(net6079),
.B1(net6180),
.B2(net6185),
.C1(net6188),
.C2(net6016),
.ZN(net6189)
);

SDFF_X2 c5885(
.D(net3999),
.SE(net6172),
.SI(net6183),
.CK(clk),
.Q(net6191),
.QN(net6190)
);

AOI21_X4 c5886(
.A(net6163),
.B1(net6174),
.B2(net10983),
.ZN(net6192)
);

AND3_X1 c5887(
.A1(net5040),
.A2(net6186),
.A3(net6188),
.ZN(net6193)
);

NAND3_X1 c5888(
.A1(net6187),
.A2(net6160),
.A3(net6184),
.ZN(net6194)
);

NOR3_X4 c5889(
.A1(net4113),
.A2(net6194),
.A3(net6185),
.ZN(net6195)
);

NOR3_X2 c5890(
.A1(net6192),
.A2(net6193),
.A3(net6185),
.ZN(net6196)
);

SDFFRS_X2 c5891(
.D(net5141),
.RN(net6184),
.SE(net5157),
.SI(net6196),
.SN(net6179),
.CK(clk),
.Q(net6198),
.QN(net6197)
);

AND3_X4 c5892(
.A1(net6198),
.A2(net6196),
.A3(net10899),
.ZN(net6199)
);

INV_X1 c5893(
.A(net10983),
.ZN(net6200)
);

NAND2_X1 c5894(
.A1(net6081),
.A2(net1392),
.ZN(net6201)
);

INV_X2 c5895(
.A(net1381),
.ZN(net6202)
);

INV_X8 c5896(
.A(net9733),
.ZN(net6203)
);

INV_X16 c5897(
.A(net9680),
.ZN(net6204)
);

INV_X32 c5898(
.A(net5219),
.ZN(net6205)
);

INV_X4 c5899(
.A(net6139),
.ZN(net6206)
);

NAND2_X2 c5900(
.A1(net5244),
.A2(net6180),
.ZN(net6207)
);

NAND3_X2 c5901(
.A1(net6203),
.A2(net6144),
.A3(net6149),
.ZN(net6208)
);

DFFRS_X1 c5902(
.D(net6205),
.RN(net6093),
.SN(net6201),
.CK(clk),
.Q(net6210),
.QN(net6209)
);

INV_X1 c5903(
.A(net6188),
.ZN(net6211)
);

NAND2_X4 c5904(
.A1(net5303),
.A2(net6016),
.ZN(net6212)
);

AND2_X2 c5905(
.A1(net6188),
.A2(net10614),
.ZN(net6213)
);

INV_X2 c5906(
.A(net5228),
.ZN(net6214)
);

OR3_X1 c5907(
.A1(net5294),
.A2(net4261),
.A3(net4312),
.ZN(net6215)
);

INV_X8 c5908(
.A(net9679),
.ZN(net6216)
);

DFFR_X1 c5909(
.D(net6130),
.RN(net6216),
.CK(clk),
.Q(net6218),
.QN(net6217)
);

INV_X16 c5910(
.A(net11071),
.ZN(net6219)
);

INV_X32 c5911(
.A(net9707),
.ZN(net6220)
);

XOR2_X1 c5912(
.A(net6216),
.B(net1236),
.Z(net6221)
);

INV_X4 c5913(
.A(net10081),
.ZN(net6222)
);

INV_X1 c5914(
.A(net5239),
.ZN(net6223)
);

INV_X2 c5915(
.A(net5818),
.ZN(net6224)
);

DFFR_X2 c5916(
.D(net5311),
.RN(net6212),
.CK(clk),
.Q(net6226),
.QN(net6225)
);

INV_X8 c5917(
.A(net6150),
.ZN(net6227)
);

NOR2_X1 c5918(
.A1(net5242),
.A2(net11071),
.ZN(net6228)
);

OR2_X2 c5919(
.A1(net5127),
.A2(net6200),
.ZN(net6229)
);

NOR2_X4 c5920(
.A1(net6219),
.A2(net6139),
.ZN(net6230)
);

INV_X16 c5921(
.A(net9749),
.ZN(net6231)
);

NOR2_X2 c5922(
.A1(net6204),
.A2(net5236),
.ZN(net6232)
);

MUX2_X1 c5923(
.A(net6220),
.B(net5239),
.S(net6016),
.Z(net6233)
);

OAI21_X4 c5924(
.A(net6230),
.B1(net6203),
.B2(net6225),
.ZN(net6234)
);

DFFS_X1 c5925(
.D(net5209),
.SN(net6218),
.CK(clk),
.Q(net6236),
.QN(net6235)
);

XOR2_X2 c5926(
.A(net5216),
.B(net6083),
.Z(net6237)
);

XNOR2_X1 c5927(
.A(net6217),
.B(net10454),
.ZN(net6238)
);

OR2_X4 c5928(
.A1(net6206),
.A2(net6215),
.ZN(net6239)
);

INV_X32 c5929(
.A(net4284),
.ZN(net6240)
);

OR2_X1 c5930(
.A1(net4312),
.A2(net6238),
.ZN(net6241)
);

DFFS_X2 c5931(
.D(net6207),
.SN(net6200),
.CK(clk),
.Q(net6243),
.QN(net6242)
);

XNOR2_X2 c5932(
.A(net5302),
.B(net4145),
.ZN(net6244)
);

AND2_X4 c5933(
.A1(net6215),
.A2(net4338),
.ZN(net6245)
);

NOR4_X2 c5934(
.A1(net6224),
.A2(net6226),
.A3(net5296),
.A4(net6180),
.ZN(net6246)
);

AOI211_X4 c5935(
.A(net6223),
.B(net6230),
.C1(net6188),
.C2(net6213),
.ZN(net6247)
);

AND2_X1 c5936(
.A1(net3210),
.A2(net6204),
.ZN(net6248)
);

INV_X4 c5937(
.A(net10020),
.ZN(net6249)
);

NAND2_X1 c5938(
.A1(net6209),
.A2(net10454),
.ZN(net6250)
);

NAND2_X2 c5939(
.A1(net4291),
.A2(net6200),
.ZN(net6251)
);

INV_X1 c5940(
.A(net6250),
.ZN(net6252)
);

MUX2_X2 c5941(
.A(net6203),
.B(net5242),
.S(net10933),
.Z(net6253)
);

NAND2_X4 c5942(
.A1(net6229),
.A2(net5190),
.ZN(net6254)
);

INV_X2 c5943(
.A(net11130),
.ZN(net6255)
);

AND2_X2 c5944(
.A1(net6237),
.A2(net5166),
.ZN(net6256)
);

XOR2_X1 c5945(
.A(net6227),
.B(net6238),
.Z(net6257)
);

INV_X8 c5946(
.A(net10294),
.ZN(net6258)
);

NOR2_X1 c5947(
.A1(net6231),
.A2(net6257),
.ZN(net6259)
);

OR2_X2 c5948(
.A1(net6241),
.A2(net6223),
.ZN(net6260)
);

NOR2_X4 c5949(
.A1(net6214),
.A2(net6260),
.ZN(net6261)
);

NOR2_X2 c5950(
.A1(net5250),
.A2(net6083),
.ZN(net6262)
);

CLKGATETST_X1 c5951(
.E(net4304),
.SE(net6196),
.CK(clk),
.GCK(net6263)
);

XOR2_X2 c5952(
.A(net6262),
.B(net6230),
.Z(net6264)
);

XNOR2_X1 c5953(
.A(net5310),
.B(net6243),
.ZN(net6265)
);

OR2_X4 c5954(
.A1(net6252),
.A2(net6263),
.ZN(net6266)
);

OAI221_X2 c5955(
.A(net6257),
.B1(net6036),
.B2(net5303),
.C1(net6264),
.C2(net5284),
.ZN(net6267)
);

NOR4_X1 c5956(
.A1(net6144),
.A2(net6263),
.A3(net6264),
.A4(net6267),
.ZN(net6268)
);

INV_X16 c5957(
.A(net6264),
.ZN(net6269)
);

NAND3_X4 c5958(
.A1(net6211),
.A2(net6263),
.A3(net6222),
.ZN(net6270)
);

OR2_X1 c5959(
.A1(net6263),
.A2(net6206),
.ZN(net6271)
);

XNOR2_X2 c5960(
.A(net4279),
.B(net6259),
.ZN(net6272)
);

AND2_X4 c5961(
.A1(net6271),
.A2(net6240),
.ZN(net6273)
);

OAI222_X4 c5962(
.A1(net4288),
.A2(net6236),
.B1(net6267),
.B2(net5239),
.C1(net5315),
.C2(net6253),
.ZN(net6274)
);

AOI211_X2 c5963(
.A(net5872),
.B(net4342),
.C1(net6229),
.C2(net6083),
.ZN(net6275)
);

AND2_X1 c5964(
.A1(net5162),
.A2(net6225),
.ZN(net6276)
);

OR3_X4 c5965(
.A1(net6247),
.A2(net6229),
.A3(net6264),
.ZN(net6277)
);

AND3_X2 c5966(
.A1(net6258),
.A2(net6275),
.A3(net6273),
.ZN(net6278)
);

AOI22_X1 c5967(
.A1(net6269),
.A2(net6223),
.B1(net6267),
.B2(net5283),
.ZN(net6279)
);

NOR3_X1 c5968(
.A1(net6268),
.A2(net6277),
.A3(net5294),
.ZN(net6280)
);

NAND2_X1 c5969(
.A1(net6245),
.A2(net11100),
.ZN(net6281)
);

NAND2_X2 c5970(
.A1(net6272),
.A2(net6259),
.ZN(net6282)
);

OR3_X2 c5971(
.A1(net6270),
.A2(net6281),
.A3(net10756),
.ZN(net6283)
);

NAND2_X4 c5972(
.A1(net6200),
.A2(net6282),
.ZN(net6284)
);

OAI21_X2 c5973(
.A(net6278),
.B1(net6260),
.B2(net6277),
.ZN(net6285)
);

OAI21_X1 c5974(
.A(net6281),
.B1(net6266),
.B2(net6275),
.ZN(net6286)
);

AOI221_X4 c5975(
.A(net6267),
.B1(net3383),
.B2(net6286),
.C1(net6183),
.C2(net11032),
.ZN(net6287)
);

AND2_X2 c5976(
.A1(net5099),
.A2(net6270),
.ZN(net6288)
);

INV_X32 c5977(
.A(net9846),
.ZN(net6289)
);

INV_X4 c5978(
.A(net6234),
.ZN(net6290)
);

INV_X1 c5979(
.A(net9588),
.ZN(net6291)
);

XOR2_X1 c5980(
.A(net5334),
.B(net6218),
.Z(net6292)
);

NOR2_X1 c5981(
.A1(net6255),
.A2(net6242),
.ZN(net6293)
);

OR2_X2 c5982(
.A1(net6259),
.A2(net6201),
.ZN(net6294)
);

INV_X2 c5983(
.A(net6201),
.ZN(net6295)
);

NOR2_X4 c5984(
.A1(net5283),
.A2(net10711),
.ZN(net6296)
);

INV_X8 c5985(
.A(net10041),
.ZN(net6297)
);

INV_X16 c5986(
.A(net6294),
.ZN(net6298)
);

INV_X32 c5987(
.A(net5344),
.ZN(net6299)
);

NOR2_X2 c5988(
.A1(net6202),
.A2(net5321),
.ZN(net6300)
);

INV_X4 c5989(
.A(net5399),
.ZN(net6301)
);

INV_X1 c5990(
.A(net6292),
.ZN(net6302)
);

XOR2_X2 c5991(
.A(net6236),
.B(net6270),
.Z(net6303)
);

AOI21_X2 c5992(
.A(net6267),
.B1(net6301),
.B2(net5355),
.ZN(net6304)
);

XNOR2_X1 c5993(
.A(net5378),
.B(net6293),
.ZN(net6305)
);

INV_X2 c5994(
.A(net6291),
.ZN(net6306)
);

OR2_X4 c5995(
.A1(net5886),
.A2(net5266),
.ZN(net6307)
);

OR2_X1 c5996(
.A1(net5323),
.A2(net6074),
.ZN(net6308)
);

XNOR2_X2 c5997(
.A(net5337),
.B(net6180),
.ZN(net6309)
);

INV_X8 c5998(
.A(net6180),
.ZN(net6310)
);

AOI21_X1 c5999(
.A(net6270),
.B1(net6253),
.B2(net5166),
.ZN(net6311)
);

INV_X16 c6000(
.A(net5405),
.ZN(net6312)
);

DFFRS_X2 c6001(
.D(net5889),
.RN(net6312),
.SN(net5340),
.CK(clk),
.Q(net6314),
.QN(net6313)
);

AND2_X4 c6002(
.A1(net6300),
.A2(net5253),
.ZN(net6315)
);

INV_X32 c6003(
.A(net10197),
.ZN(net6316)
);

AND2_X1 c6004(
.A1(net4360),
.A2(net6302),
.ZN(net6317)
);

NAND2_X1 c6005(
.A1(net2473),
.A2(net4388),
.ZN(net6318)
);

INV_X4 c6006(
.A(net9588),
.ZN(net6319)
);

NAND2_X2 c6007(
.A1(net6243),
.A2(net5346),
.ZN(net6320)
);

NAND2_X4 c6008(
.A1(net6293),
.A2(net6302),
.ZN(net6321)
);

AND2_X2 c6009(
.A1(net6286),
.A2(net4350),
.ZN(net6322)
);

INV_X1 c6010(
.A(net10602),
.ZN(net6323)
);

INV_X2 c6011(
.A(net10276),
.ZN(net6324)
);

XOR2_X1 c6012(
.A(net6074),
.B(net6322),
.Z(net6325)
);

INV_X8 c6013(
.A(net6320),
.ZN(net6326)
);

NOR2_X1 c6014(
.A1(net6319),
.A2(net4360),
.ZN(net6327)
);

OR2_X2 c6015(
.A1(net6289),
.A2(net5886),
.ZN(net6328)
);

NOR2_X4 c6016(
.A1(net6321),
.A2(net6198),
.ZN(net6329)
);

AND4_X4 c6017(
.A1(net6295),
.A2(net5156),
.A3(net5163),
.A4(net6222),
.ZN(net6330)
);

NOR2_X2 c6018(
.A1(net4416),
.A2(net6286),
.ZN(net6331)
);

XOR2_X2 c6019(
.A(net6261),
.B(net6267),
.Z(net6332)
);

XNOR2_X1 c6020(
.A(net6327),
.B(net5253),
.ZN(net6333)
);

OR2_X4 c6021(
.A1(net5953),
.A2(net6329),
.ZN(net6334)
);

AOI21_X4 c6022(
.A(net5266),
.B1(net5331),
.B2(net5405),
.ZN(net6335)
);

INV_X16 c6023(
.A(net9948),
.ZN(net6336)
);

AND3_X1 c6024(
.A1(net5377),
.A2(net6325),
.A3(net6138),
.ZN(net6337)
);

OR2_X1 c6025(
.A1(net6319),
.A2(net10786),
.ZN(net6338)
);

XNOR2_X2 c6026(
.A(net5266),
.B(net10602),
.ZN(net6339)
);

AND2_X4 c6027(
.A1(net6326),
.A2(net10438),
.ZN(net6340)
);

AND2_X1 c6028(
.A1(net5357),
.A2(net6286),
.ZN(net6341)
);

NAND2_X1 c6029(
.A1(net5384),
.A2(net6316),
.ZN(net6342)
);

NAND3_X1 c6030(
.A1(net6325),
.A2(net6336),
.A3(net6313),
.ZN(net6343)
);

INV_X32 c6031(
.A(net11114),
.ZN(net6344)
);

NAND2_X2 c6032(
.A1(net6341),
.A2(net6158),
.ZN(net6345)
);

INV_X4 c6033(
.A(net10123),
.ZN(net6346)
);

NAND2_X4 c6034(
.A1(net6340),
.A2(net4425),
.ZN(net6347)
);

AND2_X2 c6035(
.A1(net5823),
.A2(net5321),
.ZN(net6348)
);

SDFFS_X1 c6036(
.D(net6138),
.SE(net6344),
.SI(net5953),
.SN(net5166),
.CK(clk),
.Q(net6350),
.QN(net6349)
);

NOR3_X4 c6037(
.A1(net4388),
.A2(net6339),
.A3(net6344),
.ZN(net6351)
);

XOR2_X1 c6038(
.A(net6287),
.B(net5399),
.Z(net6352)
);

NOR2_X1 c6039(
.A1(net6317),
.A2(net6344),
.ZN(net6353)
);

OR2_X2 c6040(
.A1(net6304),
.A2(net6295),
.ZN(net6354)
);

NOR2_X4 c6041(
.A1(net6346),
.A2(net6351),
.ZN(net6355)
);

NOR2_X2 c6042(
.A1(net5354),
.A2(net6233),
.ZN(net6356)
);

INV_X1 c6043(
.A(net10908),
.ZN(net6357)
);

NOR3_X2 c6044(
.A1(net6336),
.A2(net6351),
.A3(net6342),
.ZN(net6358)
);

XOR2_X2 c6045(
.A(net6338),
.B(net6355),
.Z(net6359)
);

AND3_X4 c6046(
.A1(net6314),
.A2(net5344),
.A3(net6356),
.ZN(net6360)
);

INV_X2 c6047(
.A(net10246),
.ZN(net6361)
);

AOI221_X2 c6048(
.A(net6348),
.B1(net6355),
.B2(net6359),
.C1(net6316),
.C2(net6356),
.ZN(net6362)
);

XNOR2_X1 c6049(
.A(net6347),
.B(net6349),
.ZN(net6363)
);

OR2_X4 c6050(
.A1(net6335),
.A2(net6351),
.ZN(net6364)
);

AOI221_X1 c6051(
.A(net6331),
.B1(net5378),
.B2(net6348),
.C1(net6344),
.C2(net6359),
.ZN(net6365)
);

SDFF_X1 c6052(
.D(net6365),
.SE(net6331),
.SI(net6359),
.CK(clk),
.Q(net6367),
.QN(net6366)
);

OR2_X1 c6053(
.A1(net6355),
.A2(net6335),
.ZN(net6368)
);

SDFFRS_X1 c6054(
.D(net6322),
.RN(net6357),
.SE(net6353),
.SI(net6366),
.SN(net6253),
.CK(clk),
.Q(net6370),
.QN(net6369)
);

XNOR2_X2 c6055(
.A(net6352),
.B(net6366),
.ZN(net6371)
);

AND2_X4 c6056(
.A1(net6363),
.A2(net6317),
.ZN(net6372)
);

INV_X8 c6057(
.A(net9800),
.ZN(net6373)
);

OAI221_X1 c6058(
.A(net6343),
.B1(net6373),
.B2(net6297),
.C1(net6361),
.C2(net5345),
.ZN(net6374)
);

INV_X16 c6059(
.A(net10036),
.ZN(net6375)
);

INV_X32 c6060(
.A(net6364),
.ZN(net6376)
);

INV_X4 c6061(
.A(net6299),
.ZN(net6377)
);

AND2_X1 c6062(
.A1(net5385),
.A2(net5307),
.ZN(net6378)
);

NAND3_X2 c6063(
.A1(net4395),
.A2(net5474),
.A3(net10408),
.ZN(net6379)
);

INV_X1 c6064(
.A(net9638),
.ZN(net6380)
);

NAND2_X1 c6065(
.A1(net5253),
.A2(net5466),
.ZN(net6381)
);

INV_X2 c6066(
.A(net3399),
.ZN(net6382)
);

INV_X8 c6067(
.A(net10185),
.ZN(net6383)
);

NAND2_X2 c6068(
.A1(net6185),
.A2(net6357),
.ZN(net6384)
);

OR3_X1 c6069(
.A1(net6376),
.A2(net6384),
.A3(net6383),
.ZN(net6385)
);

NAND2_X4 c6070(
.A1(net4477),
.A2(net5160),
.ZN(net6386)
);

INV_X16 c6071(
.A(net3548),
.ZN(net6387)
);

AND2_X2 c6072(
.A1(net5437),
.A2(net5425),
.ZN(net6388)
);

INV_X32 c6073(
.A(net6375),
.ZN(net6389)
);

MUX2_X1 c6074(
.A(net5456),
.B(net4499),
.S(net6382),
.Z(net6390)
);

INV_X4 c6075(
.A(net5164),
.ZN(net6391)
);

INV_X1 c6076(
.A(net10218),
.ZN(net6392)
);

INV_X2 c6077(
.A(net10024),
.ZN(net6393)
);

XOR2_X1 c6078(
.A(net6357),
.B(net6381),
.Z(net6394)
);

INV_X8 c6079(
.A(net6298),
.ZN(net6395)
);

NOR2_X1 c6080(
.A1(net6308),
.A2(net6316),
.ZN(net6396)
);

OR2_X2 c6081(
.A1(net6396),
.A2(net5381),
.ZN(net6397)
);

NOR2_X4 c6082(
.A1(net6368),
.A2(net6337),
.ZN(net6398)
);

INV_X16 c6083(
.A(net10088),
.ZN(net6399)
);

INV_X32 c6084(
.A(net6392),
.ZN(net6400)
);

INV_X4 c6085(
.A(net10284),
.ZN(net6401)
);

INV_X1 c6086(
.A(net9637),
.ZN(net6402)
);

OAI21_X4 c6087(
.A(net4395),
.B1(net6390),
.B2(net4329),
.ZN(net6403)
);

NOR2_X2 c6088(
.A1(net5466),
.A2(net4379),
.ZN(net6404)
);

XOR2_X2 c6089(
.A(net6393),
.B(net6388),
.Z(net6405)
);

XNOR2_X1 c6090(
.A(net5356),
.B(net6404),
.ZN(net6406)
);

OR2_X4 c6091(
.A1(net5427),
.A2(net6404),
.ZN(net6407)
);

MUX2_X2 c6092(
.A(net5465),
.B(net6378),
.S(net5432),
.Z(net6408)
);

INV_X2 c6093(
.A(net10250),
.ZN(net6409)
);

OR2_X1 c6094(
.A1(net6394),
.A2(net6405),
.ZN(net6410)
);

XNOR2_X2 c6095(
.A(net6377),
.B(net6147),
.ZN(net6411)
);

AND2_X4 c6096(
.A1(net6404),
.A2(net6342),
.ZN(net6412)
);

SDFF_X2 c6097(
.D(net6339),
.SE(net6409),
.SI(net6403),
.CK(clk),
.Q(net6414),
.QN(net6413)
);

AND2_X1 c6098(
.A1(net1579),
.A2(net11036),
.ZN(net6415)
);

INV_X8 c6099(
.A(net11036),
.ZN(net6416)
);

NAND2_X1 c6100(
.A1(net6402),
.A2(net5307),
.ZN(net6417)
);

INV_X16 c6101(
.A(net10022),
.ZN(net6418)
);

NAND2_X2 c6102(
.A1(net6415),
.A2(net5160),
.ZN(net6419)
);

NAND2_X4 c6103(
.A1(net5432),
.A2(net6415),
.ZN(net6420)
);

AND2_X2 c6104(
.A1(net6323),
.A2(net5359),
.ZN(net6421)
);

NAND3_X4 c6105(
.A1(net6256),
.A2(net6404),
.A3(net10758),
.ZN(net6422)
);

DFFRS_X1 c6106(
.D(net5431),
.RN(net6402),
.SN(net6419),
.CK(clk),
.Q(net6424),
.QN(net6423)
);

XOR2_X1 c6107(
.A(net6406),
.B(net10497),
.Z(net6425)
);

NOR2_X1 c6108(
.A1(net6389),
.A2(net11036),
.ZN(net6426)
);

OR2_X2 c6109(
.A1(net2593),
.A2(net6426),
.ZN(net6427)
);

NOR2_X4 c6110(
.A1(net4510),
.A2(net6412),
.ZN(net6428)
);

NOR2_X2 c6111(
.A1(net6426),
.A2(net10615),
.ZN(net6429)
);

XOR2_X2 c6112(
.A(net6389),
.B(net5385),
.Z(net6430)
);

XNOR2_X1 c6113(
.A(net6420),
.B(net6401),
.ZN(net6431)
);

INV_X32 c6114(
.A(net10046),
.ZN(net6432)
);

OR2_X4 c6115(
.A1(net6421),
.A2(net6429),
.ZN(net6433)
);

OR2_X1 c6116(
.A1(net2546),
.A2(net6364),
.ZN(net6434)
);

OR3_X4 c6117(
.A1(net6430),
.A2(net5437),
.A3(net6083),
.ZN(net6435)
);

OAI222_X2 c6118(
.A1(net6422),
.A2(net6083),
.B1(net6394),
.B2(net5355),
.C1(net5345),
.C2(net6405),
.ZN(net6436)
);

XNOR2_X2 c6119(
.A(net6409),
.B(net6393),
.ZN(net6437)
);

DFFRS_X2 c6120(
.D(net6431),
.RN(net6378),
.SN(net5440),
.CK(clk),
.Q(net6439),
.QN(net6438)
);

NAND4_X1 c6121(
.A1(net6384),
.A2(net6437),
.A3(net6436),
.A4(net6438),
.ZN(net6440)
);

AOI222_X1 c6122(
.A1(net6437),
.A2(net6404),
.B1(net6423),
.B2(net6412),
.C1(net5485),
.C2(net6342),
.ZN(net6441)
);

AND3_X2 c6123(
.A1(net5356),
.A2(net6426),
.A3(net10631),
.ZN(net6442)
);

NOR3_X1 c6124(
.A1(net6312),
.A2(net6403),
.A3(net6429),
.ZN(net6443)
);

INV_X4 c6125(
.A(net10969),
.ZN(net6444)
);

AND2_X4 c6126(
.A1(net6429),
.A2(net6420),
.ZN(net6445)
);

OR4_X1 c6127(
.A1(net5321),
.A2(net3532),
.A3(net5486),
.A4(net11109),
.ZN(net6446)
);

OR3_X2 c6128(
.A1(net6445),
.A2(net6429),
.A3(net10496),
.ZN(net6447)
);

OAI21_X2 c6129(
.A(net6436),
.B1(net6439),
.B2(net6426),
.ZN(net6448)
);

OAI21_X1 c6130(
.A(net6445),
.B1(net4329),
.B2(net10759),
.ZN(net6449)
);

AND2_X1 c6131(
.A1(net6424),
.A2(net10831),
.ZN(net6450)
);

AOI21_X2 c6132(
.A(net6324),
.B1(net6426),
.B2(net6450),
.ZN(net6451)
);

OAI221_X4 c6133(
.A(net6016),
.B1(net6406),
.B2(net6429),
.C1(net6450),
.C2(net6381),
.ZN(net6452)
);

NAND2_X1 c6134(
.A1(net6424),
.A2(net6376),
.ZN(net6453)
);

INV_X1 c6135(
.A(net10348),
.ZN(net6454)
);

INV_X2 c6136(
.A(net9974),
.ZN(net6455)
);

AOI21_X1 c6137(
.A(net6406),
.B1(net6450),
.B2(net6429),
.ZN(net6456)
);

SDFF_X1 c6138(
.D(net6455),
.SE(net6456),
.SI(net4479),
.CK(clk),
.Q(net6458),
.QN(net6457)
);

AOI21_X4 c6139(
.A(net6306),
.B1(net6432),
.B2(net6413),
.ZN(net6459)
);

AND3_X1 c6140(
.A1(net6407),
.A2(net6458),
.A3(net6450),
.ZN(net6460)
);

SDFF_X2 c6141(
.D(net6459),
.SE(net6453),
.SI(net6450),
.CK(clk),
.Q(net6462),
.QN(net6461)
);

INV_X8 c6142(
.A(net11071),
.ZN(net6463)
);

INV_X16 c6143(
.A(net5494),
.ZN(net6464)
);

INV_X32 c6144(
.A(net10298),
.ZN(net6465)
);

INV_X4 c6145(
.A(net11133),
.ZN(net6466)
);

INV_X1 c6146(
.A(net9757),
.ZN(net6467)
);

NAND2_X2 c6147(
.A1(net5285),
.A2(net6466),
.ZN(net6468)
);

INV_X2 c6148(
.A(net5575),
.ZN(net6469)
);

NAND2_X4 c6149(
.A1(net4544),
.A2(net5503),
.ZN(net6470)
);

INV_X8 c6150(
.A(net10754),
.ZN(net6471)
);

AND2_X2 c6151(
.A1(net5359),
.A2(net10708),
.ZN(net6472)
);

INV_X16 c6152(
.A(net5440),
.ZN(net6473)
);

XOR2_X1 c6153(
.A(net5160),
.B(net6466),
.Z(net6474)
);

CLKGATETST_X2 c6154(
.E(net5565),
.SE(net5515),
.CK(clk),
.GCK(net6475)
);

INV_X32 c6155(
.A(net9635),
.ZN(net6476)
);

NOR2_X1 c6156(
.A1(net6390),
.A2(net5486),
.ZN(net6477)
);

OR2_X2 c6157(
.A1(net6475),
.A2(net10733),
.ZN(net6478)
);

NOR2_X4 c6158(
.A1(net5505),
.A2(net4544),
.ZN(net6479)
);

NOR2_X2 c6159(
.A1(net6462),
.A2(net4425),
.ZN(net6480)
);

INV_X4 c6160(
.A(net9871),
.ZN(net6481)
);

XOR2_X2 c6161(
.A(net5941),
.B(net5491),
.Z(net6482)
);

XNOR2_X1 c6162(
.A(net5524),
.B(net4379),
.ZN(net6483)
);

OR2_X4 c6163(
.A1(net6449),
.A2(net5380),
.ZN(net6484)
);

INV_X1 c6164(
.A(net9967),
.ZN(net6485)
);

INV_X2 c6165(
.A(net9635),
.ZN(net6486)
);

OR2_X1 c6166(
.A1(net5359),
.A2(net6467),
.ZN(net6487)
);

XNOR2_X2 c6167(
.A(net6468),
.B(net5562),
.ZN(net6488)
);

AND2_X4 c6168(
.A1(net5510),
.A2(net6475),
.ZN(net6489)
);

AND2_X1 c6169(
.A1(net6480),
.A2(net6472),
.ZN(net6490)
);

NAND2_X1 c6170(
.A1(net6083),
.A2(net5530),
.ZN(net6491)
);

INV_X8 c6171(
.A(net5380),
.ZN(net6492)
);

NAND2_X2 c6172(
.A1(net4572),
.A2(net6470),
.ZN(net6493)
);

INV_X16 c6173(
.A(net11058),
.ZN(net6494)
);

INV_X32 c6174(
.A(net4379),
.ZN(net6495)
);

NAND2_X4 c6175(
.A1(net6382),
.A2(net5531),
.ZN(net6496)
);

OAI221_X2 c6176(
.A(net6465),
.B1(net6466),
.B2(net6467),
.C1(net6337),
.C2(net11071),
.ZN(net6497)
);

AND2_X2 c6177(
.A1(net3617),
.A2(net6495),
.ZN(net6498)
);

XOR2_X1 c6178(
.A(net6494),
.B(net5494),
.Z(net6499)
);

NOR2_X1 c6179(
.A1(net5541),
.A2(net4031),
.ZN(net6500)
);

OR2_X2 c6180(
.A1(net6500),
.A2(net5439),
.ZN(net6501)
);

NAND3_X1 c6181(
.A1(net6493),
.A2(net6483),
.A3(net5544),
.ZN(net6502)
);

INV_X4 c6182(
.A(net6470),
.ZN(net6503)
);

NOR2_X4 c6183(
.A1(net6498),
.A2(net4540),
.ZN(net6504)
);

NOR2_X2 c6184(
.A1(net4591),
.A2(net6502),
.ZN(net6505)
);

INV_X1 c6185(
.A(net6383),
.ZN(net6506)
);

XOR2_X2 c6186(
.A(net6486),
.B(net5285),
.Z(net6507)
);

XNOR2_X1 c6187(
.A(net3624),
.B(net6494),
.ZN(net6508)
);

NOR3_X4 c6188(
.A1(net6496),
.A2(net6462),
.A3(net6475),
.ZN(net6509)
);

NOR3_X2 c6189(
.A1(net6463),
.A2(net6485),
.A3(net11080),
.ZN(net6510)
);

OR2_X4 c6190(
.A1(net6482),
.A2(net6500),
.ZN(net6511)
);

OR2_X1 c6191(
.A1(net6495),
.A2(net6510),
.ZN(net6512)
);

XNOR2_X2 c6192(
.A(net6503),
.B(net6510),
.ZN(net6513)
);

AND2_X4 c6193(
.A1(net6380),
.A2(net5493),
.ZN(net6514)
);

AND2_X1 c6194(
.A1(net6427),
.A2(net6487),
.ZN(net6515)
);

INV_X2 c6195(
.A(net6481),
.ZN(net6516)
);

INV_X8 c6196(
.A(net9997),
.ZN(net6517)
);

NAND2_X1 c6197(
.A1(net6507),
.A2(net6489),
.ZN(net6518)
);

NAND2_X2 c6198(
.A1(net6490),
.A2(net6457),
.ZN(net6519)
);

INV_X16 c6199(
.A(net11073),
.ZN(net6520)
);

AND3_X4 c6200(
.A1(net6519),
.A2(net6520),
.A3(net6405),
.ZN(net6521)
);

NAND2_X4 c6201(
.A1(net6499),
.A2(net6520),
.ZN(net6522)
);

NAND3_X2 c6202(
.A1(net6471),
.A2(net6507),
.A3(net5565),
.ZN(net6523)
);

INV_X32 c6203(
.A(net11062),
.ZN(net6524)
);

AND2_X2 c6204(
.A1(net6506),
.A2(net6463),
.ZN(net6525)
);

XOR2_X1 c6205(
.A(net6512),
.B(net6316),
.Z(net6526)
);

OR3_X1 c6206(
.A1(net6478),
.A2(net6518),
.A3(net6496),
.ZN(net6527)
);

NOR2_X1 c6207(
.A1(net6475),
.A2(net6427),
.ZN(net6528)
);

OR2_X2 c6208(
.A1(net6515),
.A2(net6470),
.ZN(net6529)
);

NOR2_X4 c6209(
.A1(net6522),
.A2(net6503),
.ZN(net6530)
);

MUX2_X1 c6210(
.A(net6516),
.B(net6518),
.S(net6520),
.Z(net6531)
);

NOR2_X2 c6211(
.A1(net6524),
.A2(net6515),
.ZN(net6532)
);

OAI21_X4 c6212(
.A(net6531),
.B1(net6520),
.B2(net10619),
.ZN(net6533)
);

MUX2_X2 c6213(
.A(net6458),
.B(net6525),
.S(net5973),
.Z(net6534)
);

AOI222_X4 c6214(
.A1(net6502),
.A2(net6531),
.B1(net6487),
.B2(net6083),
.C1(net2569),
.C2(net5544),
.ZN(net6535)
);

NAND3_X4 c6215(
.A1(net6531),
.A2(net6533),
.A3(net6518),
.ZN(net6536)
);

OR3_X4 c6216(
.A1(net6419),
.A2(net6380),
.A3(net6510),
.ZN(net6537)
);

AND3_X2 c6217(
.A1(net6290),
.A2(net6507),
.A3(net6484),
.ZN(net6538)
);

NOR3_X1 c6218(
.A1(net6528),
.A2(net1708),
.A3(net11139),
.ZN(net6539)
);

OR3_X2 c6219(
.A1(net6513),
.A2(net6530),
.A3(net6534),
.ZN(net6540)
);

OAI33_X1 c6220(
.A1(net6536),
.A2(net6515),
.A3(net6533),
.B1(net6452),
.B2(net6525),
.B3(net6467),
.ZN(net6541)
);

AOI222_X2 c6221(
.A1(net6538),
.A2(net6483),
.B1(net6405),
.B2(net6464),
.C1(net11139),
.C2(net11200),
.ZN(net6542)
);

OAI21_X2 c6222(
.A(net6532),
.B1(net6495),
.B2(net11200),
.ZN(net6543)
);

OAI21_X1 c6223(
.A(net6539),
.B1(net6542),
.B2(net11201),
.ZN(net6544)
);

AOI21_X2 c6224(
.A(net6520),
.B1(net6543),
.B2(net11201),
.ZN(net6545)
);

AOI21_X1 c6225(
.A(net5649),
.B1(net3698),
.B2(net5633),
.ZN(net6546)
);

XOR2_X2 c6226(
.A(net2674),
.B(net6546),
.Z(net6547)
);

XNOR2_X1 c6227(
.A(net5572),
.B(net5346),
.ZN(net6548)
);

INV_X4 c6228(
.A(net10370),
.ZN(net6549)
);

INV_X1 c6229(
.A(net5627),
.ZN(net6550)
);

OR2_X4 c6230(
.A1(net4600),
.A2(net5491),
.ZN(net6551)
);

INV_X2 c6231(
.A(net9653),
.ZN(net6552)
);

OR2_X1 c6232(
.A1(net5492),
.A2(out1),
.ZN(net6553)
);

INV_X8 c6233(
.A(net10942),
.ZN(net6554)
);

INV_X16 c6234(
.A(net9713),
.ZN(net6555)
);

INV_X32 c6235(
.A(net5973),
.ZN(net6556)
);

XNOR2_X2 c6236(
.A(net6551),
.B(net6467),
.ZN(net6557)
);

AND2_X4 c6237(
.A1(net5307),
.A2(net6464),
.ZN(net6558)
);

AND2_X1 c6238(
.A1(net6483),
.A2(net5590),
.ZN(net6559)
);

NAND2_X1 c6239(
.A1(net6552),
.A2(net6550),
.ZN(net6560)
);

NAND2_X2 c6240(
.A1(net4528),
.A2(net11080),
.ZN(net6561)
);

INV_X4 c6241(
.A(net9824),
.ZN(net6562)
);

INV_X1 c6242(
.A(net3656),
.ZN(net6563)
);

NAND2_X4 c6243(
.A1(net3723),
.A2(net4678),
.ZN(net6564)
);

DFFRS_X1 c6244(
.D(net5534),
.RN(net5627),
.SN(net6381),
.CK(clk),
.Q(net6566),
.QN(net6565)
);

INV_X2 c6245(
.A(net9654),
.ZN(net6567)
);

INV_X8 c6246(
.A(net6492),
.ZN(net6568)
);

AND2_X2 c6247(
.A1(net6473),
.A2(net6550),
.ZN(net6569)
);

XOR2_X1 c6248(
.A(net6562),
.B(net4655),
.Z(net6570)
);

INV_X16 c6249(
.A(net10051),
.ZN(net6571)
);

NOR2_X1 c6250(
.A1(net5661),
.A2(net6561),
.ZN(net6572)
);

OR2_X2 c6251(
.A1(net6552),
.A2(out0),
.ZN(net6573)
);

NOR2_X4 c6252(
.A1(net6539),
.A2(net6464),
.ZN(net6574)
);

INV_X32 c6253(
.A(net9905),
.ZN(net6575)
);

NOR2_X2 c6254(
.A1(net5584),
.A2(net6562),
.ZN(net6576)
);

AOI21_X4 c6255(
.A(net6574),
.B1(net6576),
.B2(net6565),
.ZN(net6577)
);

XOR2_X2 c6256(
.A(net6565),
.B(net11109),
.Z(net6578)
);

AND3_X1 c6257(
.A1(net6577),
.A2(net6569),
.A3(net5534),
.ZN(net6579)
);

INV_X4 c6258(
.A(net6510),
.ZN(net6580)
);

XNOR2_X1 c6259(
.A(net6570),
.B(net6476),
.ZN(net6581)
);

SDFFRS_X2 c6260(
.D(net6276),
.RN(net5597),
.SE(net6557),
.SI(net6562),
.SN(net5632),
.CK(clk),
.Q(net6583),
.QN(net6582)
);

OR2_X4 c6261(
.A1(net5606),
.A2(net4638),
.ZN(net6584)
);

OR2_X1 c6262(
.A1(net5531),
.A2(net5627),
.ZN(net6585)
);

INV_X1 c6263(
.A(net6416),
.ZN(net6586)
);

XNOR2_X2 c6264(
.A(net6568),
.B(net5635),
.ZN(net6587)
);

INV_X2 c6265(
.A(net6557),
.ZN(net6588)
);

DFFRS_X2 c6266(
.D(net6581),
.RN(net6557),
.SN(net6464),
.CK(clk),
.Q(net6590),
.QN(net6589)
);

NAND3_X1 c6267(
.A1(net5611),
.A2(net3723),
.A3(net5634),
.ZN(net6591)
);

AND2_X4 c6268(
.A1(net6517),
.A2(net6553),
.ZN(net6592)
);

AND2_X1 c6269(
.A1(net6576),
.A2(net6592),
.ZN(net6593)
);

INV_X8 c6270(
.A(net9691),
.ZN(net6594)
);

INV_X16 c6271(
.A(net6489),
.ZN(net6595)
);

SDFF_X1 c6272(
.D(net5621),
.SE(net6588),
.SI(net6595),
.CK(clk),
.Q(net6597),
.QN(net6596)
);

INV_X32 c6273(
.A(net11111),
.ZN(net6598)
);

NAND2_X1 c6274(
.A1(net6584),
.A2(net6562),
.ZN(net6599)
);

INV_X4 c6275(
.A(net9968),
.ZN(net6600)
);

NAND2_X2 c6276(
.A1(net6559),
.A2(net6557),
.ZN(net6601)
);

AOI221_X4 c6277(
.A(net4531),
.B1(net6433),
.B2(net5632),
.C1(net4524),
.C2(net6467),
.ZN(net6602)
);

NAND2_X4 c6278(
.A1(net6580),
.A2(net6599),
.ZN(net6603)
);

NOR3_X4 c6279(
.A1(net4639),
.A2(net6603),
.A3(net5611),
.ZN(net6604)
);

AND2_X2 c6280(
.A1(net6585),
.A2(net6484),
.ZN(net6605)
);

XOR2_X1 c6281(
.A(net2759),
.B(net10477),
.Z(net6606)
);

NOR3_X2 c6282(
.A1(net6542),
.A2(net6605),
.A3(net5629),
.ZN(net6607)
);

INV_X1 c6283(
.A(net10086),
.ZN(net6608)
);

NOR2_X1 c6284(
.A1(net4655),
.A2(net6559),
.ZN(net6609)
);

AND3_X4 c6285(
.A1(net6609),
.A2(net6568),
.A3(net6542),
.ZN(net6610)
);

OR2_X2 c6286(
.A1(net10464),
.A2(net11026),
.ZN(net6611)
);

NOR2_X4 c6287(
.A1(net6589),
.A2(net10631),
.ZN(net6612)
);

AOI221_X2 c6288(
.A(net5620),
.B1(net6414),
.B2(net3723),
.C1(net6550),
.C2(net6487),
.ZN(net6613)
);

NOR2_X2 c6289(
.A1(net5655),
.A2(net10805),
.ZN(net6614)
);

NAND3_X2 c6290(
.A1(net6590),
.A2(net6603),
.A3(net6557),
.ZN(net6615)
);

INV_X2 c6291(
.A(net9784),
.ZN(net6616)
);

OR3_X1 c6292(
.A1(net6555),
.A2(net6596),
.A3(net11026),
.ZN(net6617)
);

INV_X8 c6293(
.A(net10244),
.ZN(net6618)
);

XOR2_X2 c6294(
.A(net6598),
.B(net6608),
.Z(net6619)
);

MUX2_X1 c6295(
.A(net6545),
.B(net6617),
.S(net6600),
.Z(net6620)
);

OAI21_X4 c6296(
.A(net6617),
.B1(net6582),
.B2(net5644),
.ZN(net6621)
);

AOI221_X1 c6297(
.A(net6571),
.B1(net6612),
.B2(net5667),
.C1(net5617),
.C2(net5657),
.ZN(net6622)
);

MUX2_X2 c6298(
.A(net4676),
.B(net6584),
.S(net10860),
.Z(net6623)
);

SDFF_X2 c6299(
.D(net6623),
.SE(net6615),
.SI(net6621),
.CK(clk),
.Q(net6625),
.QN(net6624)
);

OAI22_X1 c6300(
.A1(net6594),
.A2(net5611),
.B1(net5632),
.B2(net6581),
.ZN(net6626)
);

DFFRS_X1 c6301(
.D(net6601),
.RN(net6625),
.SN(net6612),
.CK(clk),
.Q(net6628),
.QN(net6627)
);

NAND3_X4 c6302(
.A1(net6625),
.A2(net6608),
.A3(net11107),
.ZN(net6629)
);

OR3_X4 c6303(
.A1(net6504),
.A2(net6611),
.A3(net6629),
.ZN(net6630)
);

AND3_X2 c6304(
.A1(net6622),
.A2(net6621),
.A3(net6627),
.ZN(net6631)
);

NOR3_X1 c6305(
.A1(net5590),
.A2(net6631),
.A3(net6624),
.ZN(net6632)
);

INV_X16 c6306(
.A(net10143),
.ZN(net6633)
);

OR3_X2 c6307(
.A1(net6560),
.A2(net6618),
.A3(net4640),
.ZN(net6634)
);

XNOR2_X1 c6308(
.A(net5761),
.B(net6553),
.ZN(net6635)
);

AND4_X2 c6309(
.A1(net2821),
.A2(net5658),
.A3(net5761),
.A4(net3801),
.ZN(net6636)
);

OR2_X4 c6310(
.A1(net5633),
.A2(net10475),
.ZN(net6637)
);

OR2_X1 c6311(
.A1(net5677),
.A2(net4712),
.ZN(net6638)
);

OAI21_X2 c6312(
.A(net4748),
.B1(net6619),
.B2(net5712),
.ZN(net6639)
);

XNOR2_X2 c6313(
.A(net5750),
.B(net5761),
.ZN(net6640)
);

OAI21_X1 c6314(
.A(net3802),
.B1(net4720),
.B2(net5754),
.ZN(net6641)
);

AND2_X4 c6315(
.A1(net3781),
.A2(net5749),
.ZN(net6642)
);

AND2_X1 c6316(
.A1(net5710),
.A2(net5705),
.ZN(net6643)
);

INV_X32 c6317(
.A(net9686),
.ZN(out3)
);

NAND2_X1 c6318(
.A1(net5668),
.A2(net11192),
.ZN(net6644)
);

DFFRS_X2 c6319(
.D(net6479),
.RN(net6640),
.SN(net5687),
.CK(clk),
.Q(net6646),
.QN(net6645)
);

NAND2_X2 c6320(
.A1(net6546),
.A2(net6645),
.ZN(net6647)
);

SDFF_X1 c6321(
.D(net6639),
.SE(net6643),
.SI(net6592),
.CK(clk),
.Q(net6649),
.QN(net6648)
);

AOI21_X2 c6322(
.A(net6553),
.B1(net5544),
.B2(net3806),
.ZN(net6650)
);

NAND2_X4 c6323(
.A1(net5725),
.A2(net4720),
.ZN(net6651)
);

INV_X4 c6324(
.A(net9685),
.ZN(net6652)
);

AOI21_X1 c6325(
.A(net6592),
.B1(net5633),
.B2(net5668),
.ZN(net6653)
);

AND2_X2 c6326(
.A1(net5744),
.A2(net6646),
.ZN(net6654)
);

SDFF_X2 c6327(
.D(net6641),
.SE(net6566),
.SI(net6652),
.CK(clk),
.Q(net6656),
.QN(net6655)
);

AOI21_X4 c6328(
.A(net5705),
.B1(net6553),
.B2(net4700),
.ZN(net6657)
);

XOR2_X1 c6329(
.A(net5686),
.B(net10837),
.Z(net6658)
);

DFFRS_X1 c6330(
.D(net3806),
.RN(net4773),
.SN(net6116),
.CK(clk),
.Q(net6660),
.QN(net6659)
);

AND3_X1 c6331(
.A1(net5673),
.A2(net1833),
.A3(net5636),
.ZN(net6661)
);

SDFFS_X2 c6332(
.D(net6642),
.SE(net6583),
.SI(net6661),
.SN(net5474),
.CK(clk),
.Q(net6663),
.QN(net6662)
);

NAND3_X1 c6333(
.A1(net5698),
.A2(net6655),
.A3(net6632),
.ZN(net6664)
);

NOR3_X4 c6334(
.A1(net5519),
.A2(net3825),
.A3(net6464),
.ZN(net6665)
);

NOR3_X2 c6335(
.A1(net6658),
.A2(net5760),
.A3(net2803),
.ZN(net6666)
);

NOR2_X1 c6336(
.A1(net4759),
.A2(net4782),
.ZN(net6667)
);

AND3_X4 c6337(
.A1(net6660),
.A2(net6635),
.A3(net4712),
.ZN(net6668)
);

NAND3_X2 c6338(
.A1(net6595),
.A2(net4720),
.A3(net5710),
.ZN(net6669)
);

OR2_X2 c6339(
.A1(net6381),
.A2(net6660),
.ZN(net6670)
);

AND4_X1 c6340(
.A1(net5636),
.A2(net6660),
.A3(net4700),
.A4(net6619),
.ZN(net6671)
);

OR3_X1 c6341(
.A1(net6636),
.A2(net6608),
.A3(net5681),
.ZN(net6672)
);

MUX2_X1 c6342(
.A(net5686),
.B(net5738),
.S(net5682),
.Z(net6673)
);

AOI22_X4 c6343(
.A1(net6656),
.A2(net4792),
.B1(net6667),
.B2(net5719),
.ZN(net6674)
);

OAI21_X4 c6344(
.A(net6671),
.B1(net6667),
.B2(net10593),
.ZN(net6675)
);

INV_X1 c6345(
.A(net11111),
.ZN(net6676)
);

MUX2_X2 c6346(
.A(net4712),
.B(net6592),
.S(net5687),
.Z(net6677)
);

NAND3_X4 c6347(
.A1(net6665),
.A2(net6657),
.A3(net5578),
.ZN(net6678)
);

OR3_X4 c6348(
.A1(net5722),
.A2(net6667),
.A3(net3806),
.ZN(net6679)
);

AND3_X2 c6349(
.A1(net5688),
.A2(net6658),
.A3(net10873),
.ZN(net6680)
);

INV_X2 c6350(
.A(net9899),
.ZN(net6681)
);

NOR3_X1 c6351(
.A1(net5752),
.A2(net6619),
.A3(net6650),
.ZN(net6682)
);

OR3_X2 c6352(
.A1(net5739),
.A2(net6675),
.A3(net5578),
.ZN(net6683)
);

OAI21_X2 c6353(
.A(net6587),
.B1(net6667),
.B2(net4779),
.ZN(net6684)
);

NOR2_X4 c6354(
.A1(net3768),
.A2(net6667),
.ZN(net6685)
);

OAI21_X1 c6355(
.A(net6679),
.B1(net6643),
.B2(net6680),
.ZN(net6686)
);

NOR2_X2 c6356(
.A1(net6501),
.A2(net5755),
.ZN(net6687)
);

AOI21_X2 c6357(
.A(net6679),
.B1(net6687),
.B2(net10729),
.ZN(net6688)
);

XOR2_X2 c6358(
.A(net6548),
.B(net6656),
.Z(net6689)
);

AOI21_X1 c6359(
.A(net5689),
.B1(net6587),
.B2(net10668),
.ZN(net6690)
);

OAI221_X1 c6360(
.A(net6689),
.B1(net5636),
.B2(net6525),
.C1(net6680),
.C2(net10515),
.ZN(net6691)
);

AOI21_X4 c6361(
.A(net5712),
.B1(net6671),
.B2(net5509),
.ZN(net6692)
);

AND3_X1 c6362(
.A1(net6685),
.A2(net6673),
.A3(net4640),
.ZN(net6693)
);

NAND3_X1 c6363(
.A1(net6644),
.A2(net5755),
.A3(net6659),
.ZN(net6694)
);

NOR3_X4 c6364(
.A1(net6640),
.A2(net6674),
.A3(net4780),
.ZN(net6695)
);

NOR3_X2 c6365(
.A1(net6691),
.A2(net5724),
.A3(net6587),
.ZN(net6696)
);

AND3_X4 c6366(
.A1(net6692),
.A2(net6671),
.A3(net6648),
.ZN(net6697)
);

NAND3_X2 c6367(
.A1(net6694),
.A2(net6637),
.A3(net5519),
.ZN(net6698)
);

OR3_X1 c6368(
.A1(net5747),
.A2(net6697),
.A3(net6647),
.ZN(net6699)
);

MUX2_X1 c6369(
.A(net6619),
.B(net6697),
.S(net6680),
.Z(net6700)
);

OAI22_X4 c6370(
.A1(net2804),
.A2(net5744),
.B1(net6659),
.B2(net6679),
.ZN(net6701)
);

OAI21_X4 c6371(
.A(net6681),
.B1(net6699),
.B2(net6687),
.ZN(net6702)
);

DFFRS_X2 c6372(
.D(net6699),
.RN(net5636),
.SN(net6632),
.CK(clk),
.Q(net6704),
.QN(net6703)
);

MUX2_X2 c6373(
.A(net4780),
.B(net6658),
.S(net10721),
.Z(net6705)
);

SDFF_X1 c6374(
.D(net6647),
.SE(net6682),
.SI(net6662),
.CK(clk),
.Q(net6707),
.QN(net6706)
);

NAND3_X4 c6375(
.A1(net6613),
.A2(net6679),
.A3(net4700),
.ZN(net6708)
);

OR3_X4 c6376(
.A1(net6464),
.A2(net6690),
.A3(net6697),
.ZN(net6709)
);

AND3_X2 c6377(
.A1(net6705),
.A2(net6687),
.A3(net6693),
.ZN(net6710)
);

NOR3_X1 c6378(
.A1(net6669),
.A2(net5482),
.A3(net6687),
.ZN(net6711)
);

OR3_X2 c6379(
.A1(net6693),
.A2(net6667),
.A3(net6703),
.ZN(net6712)
);

OAI21_X2 c6380(
.A(net6712),
.B1(net5676),
.B2(net10722),
.ZN(net6713)
);

SDFF_X2 c6381(
.D(net6643),
.SE(net6710),
.SI(net6692),
.CK(clk),
.Q(net6715),
.QN(net6714)
);

OAI21_X1 c6382(
.A(net5692),
.B1(net6583),
.B2(net6595),
.ZN(net6716)
);

AOI21_X2 c6383(
.A(net6704),
.B1(net6709),
.B2(net10820),
.ZN(net6717)
);

DFFRS_X1 c6384(
.D(net6715),
.RN(net6717),
.SN(net10514),
.CK(clk),
.Q(net6719),
.QN(net6718)
);

AOI22_X2 c6385(
.A1(net6709),
.A2(net6695),
.B1(net6714),
.B2(net4773),
.ZN(net6720)
);

NAND4_X4 c6386(
.A1(net6663),
.A2(net6716),
.A3(net6681),
.A4(net6650),
.ZN(net6721)
);

OAI221_X4 c6387(
.A(net6654),
.B1(net6663),
.B2(net6721),
.C1(net6612),
.C2(net10795),
.ZN(net6722)
);

OAI211_X2 c6388(
.A(net6632),
.B(net6712),
.C1(net6679),
.C2(net10573),
.ZN(net6723)
);

OR4_X2 c6389(
.A1(net6717),
.A2(net6676),
.A3(net3777),
.A4(net6721),
.ZN(net6724)
);

OAI221_X2 c6390(
.A(net4700),
.B1(net6689),
.B2(net6658),
.C1(net1709),
.C2(net10642),
.ZN(net6725)
);

INV_X8 c6391(
.A(net3880),
.ZN(net6726)
);

INV_X16 c6392(
.A(net9625),
.ZN(net6727)
);

INV_X32 c6393(
.A(net4871),
.ZN(net6728)
);

XNOR2_X1 c6394(
.A(net5794),
.B(net4846),
.ZN(net6729)
);

INV_X4 c6395(
.A(net3912),
.ZN(net6730)
);

INV_X1 c6396(
.A(net4846),
.ZN(net6731)
);

INV_X2 c6397(
.A(net3860),
.ZN(net6732)
);

CLKGATETST_X4 c6398(
.E(net6726),
.SE(net5766),
.CK(clk),
.GCK(net6733)
);

OR2_X4 c6399(
.A1(net4830),
.A2(net5767),
.ZN(net6734)
);

INV_X8 c6400(
.A(net997),
.ZN(net6735)
);

INV_X16 c6401(
.A(net4805),
.ZN(net6736)
);

INV_X32 c6402(
.A(net1927),
.ZN(net6737)
);

INV_X4 c6403(
.A(net5784),
.ZN(net6738)
);

INV_X1 c6404(
.A(net6736),
.ZN(net6739)
);

INV_X2 c6405(
.A(net4830),
.ZN(net6740)
);

INV_X8 c6406(
.A(net5768),
.ZN(net6741)
);

INV_X16 c6407(
.A(net3899),
.ZN(net6742)
);

INV_X32 c6408(
.A(net6732),
.ZN(net6743)
);

INV_X4 c6409(
.A(net5774),
.ZN(net6744)
);

INV_X1 c6410(
.A(net4799),
.ZN(net6745)
);

OR2_X1 c6411(
.A1(net3856),
.A2(net11197),
.ZN(net6746)
);

INV_X2 c6412(
.A(net6737),
.ZN(net6747)
);

INV_X8 c6413(
.A(net2920),
.ZN(net6748)
);

XNOR2_X2 c6414(
.A(net5795),
.B(net5784),
.ZN(net6749)
);

INV_X16 c6415(
.A(net6744),
.ZN(net6750)
);

INV_X32 c6416(
.A(net9624),
.ZN(net6751)
);

INV_X4 c6417(
.A(net9710),
.ZN(net6752)
);

AND2_X4 c6418(
.A1(net6751),
.A2(net6735),
.ZN(net6753)
);

INV_X1 c6419(
.A(net9732),
.ZN(net6754)
);

INV_X2 c6420(
.A(net6753),
.ZN(net6755)
);

AND2_X1 c6421(
.A1(net6740),
.A2(net5848),
.ZN(net6756)
);

NAND2_X1 c6422(
.A1(net3912),
.A2(net5835),
.ZN(net6757)
);

NAND2_X2 c6423(
.A1(net5815),
.A2(net3880),
.ZN(net6758)
);

NAND2_X4 c6424(
.A1(net6730),
.A2(net6733),
.ZN(net6759)
);

AND2_X2 c6425(
.A1(net6746),
.A2(net4805),
.ZN(net6760)
);

INV_X8 c6426(
.A(net6759),
.ZN(net6761)
);

INV_X16 c6427(
.A(net6735),
.ZN(net6762)
);

XOR2_X1 c6428(
.A(net6762),
.B(net6759),
.Z(net6763)
);

NOR2_X1 c6429(
.A1(net6763),
.A2(net3912),
.ZN(net6764)
);

OR2_X2 c6430(
.A1(net6760),
.A2(net6761),
.ZN(net6765)
);

INV_X32 c6431(
.A(net9731),
.ZN(net6766)
);

NOR2_X4 c6432(
.A1(net4807),
.A2(net6763),
.ZN(net6767)
);

CLKGATETST_X8 c6433(
.E(net5838),
.SE(net5840),
.CK(clk),
.GCK(net6768)
);

INV_X4 c6434(
.A(net4849),
.ZN(net6769)
);

INV_X1 c6435(
.A(net9808),
.ZN(net6770)
);

INV_X2 c6436(
.A(net9706),
.ZN(net6771)
);

DFFRS_X2 c6437(
.D(net4799),
.RN(net6743),
.SN(net6726),
.CK(clk),
.Q(net6773),
.QN(net6772)
);

INV_X8 c6438(
.A(net10413),
.ZN(net6774)
);

INV_X16 c6439(
.A(net6771),
.ZN(net6775)
);

DFFR_X1 c6440(
.D(net6767),
.RN(net2952),
.CK(clk),
.Q(net6777),
.QN(net6776)
);

DFFR_X2 c6441(
.D(net6756),
.RN(net5829),
.CK(clk),
.Q(net6779),
.QN(net6778)
);

INV_X32 c6442(
.A(net6774),
.ZN(net6780)
);

NOR2_X2 c6443(
.A1(net6734),
.A2(net6777),
.ZN(net6781)
);

AOI21_X1 c6444(
.A(net6737),
.B1(net6771),
.B2(net6775),
.ZN(net6782)
);

XOR2_X2 c6445(
.A(net6743),
.B(net6781),
.Z(net6783)
);

XNOR2_X1 c6446(
.A(net6751),
.B(net6782),
.ZN(net6784)
);

OR2_X4 c6447(
.A1(net6747),
.A2(net6782),
.ZN(net6785)
);

AOI211_X1 c6448(
.A(net6777),
.B(net6775),
.C1(net6745),
.C2(net5848),
.ZN(net6786)
);

AOI21_X4 c6449(
.A(net5815),
.B1(net6782),
.B2(net5767),
.ZN(net6787)
);

DFFS_X1 c6450(
.D(net4845),
.SN(net6786),
.CK(clk),
.Q(net6789),
.QN(net6788)
);

DFFS_X2 c6451(
.D(net6769),
.SN(net6783),
.CK(clk),
.Q(net6791),
.QN(net6790)
);

OR2_X1 c6452(
.A1(net5840),
.A2(net6772),
.ZN(net6792)
);

XNOR2_X2 c6453(
.A(net6754),
.B(net6792),
.ZN(net6793)
);

SDFF_X1 c6454(
.D(net6731),
.SE(net6783),
.SI(net6763),
.CK(clk),
.Q(net6795),
.QN(net6794)
);

AND2_X4 c6455(
.A1(net6780),
.A2(net6794),
.ZN(net6796)
);

AND2_X1 c6456(
.A1(net6745),
.A2(net6780),
.ZN(net6797)
);

NAND2_X1 c6457(
.A1(net5794),
.A2(net6767),
.ZN(net6798)
);

NAND2_X2 c6458(
.A1(net5835),
.A2(net6796),
.ZN(net6799)
);

AND3_X1 c6459(
.A1(net6795),
.A2(net4810),
.A3(net10413),
.ZN(net6800)
);

NAND2_X4 c6460(
.A1(net6795),
.A2(net6776),
.ZN(net6801)
);

AND2_X2 c6461(
.A1(net6775),
.A2(net5843),
.ZN(net6802)
);

SDFF_X2 c6462(
.D(net6797),
.SE(net6749),
.SI(net6788),
.CK(clk),
.Q(net6804),
.QN(net6803)
);

OAI222_X1 c6463(
.A1(net6787),
.A2(net6750),
.B1(net6803),
.B2(net6726),
.C1(net6786),
.C2(net5848),
.ZN(net6805)
);

NAND3_X1 c6464(
.A1(net6742),
.A2(net6745),
.A3(net6793),
.ZN(net6806)
);

NOR3_X4 c6465(
.A1(net6796),
.A2(net5786),
.A3(net6799),
.ZN(net6807)
);

NOR3_X2 c6466(
.A1(net6770),
.A2(net6803),
.A3(net5767),
.ZN(net6808)
);

AND3_X4 c6467(
.A1(net6785),
.A2(net6753),
.A3(net6778),
.ZN(net6809)
);

NAND3_X2 c6468(
.A1(net6809),
.A2(net6806),
.A3(net11203),
.ZN(net6810)
);

OAI222_X4 c6469(
.A1(net6781),
.A2(net6810),
.B1(net6786),
.B2(net6788),
.C1(net5848),
.C2(net6730),
.ZN(net6811)
);

DFFRS_X1 c6470(
.D(net6738),
.RN(net6808),
.SN(net11205),
.CK(clk),
.Q(net6813),
.QN(net6812)
);

NAND4_X2 c6471(
.A1(net6808),
.A2(net6793),
.A3(net6806),
.A4(net11203),
.ZN(net6814)
);

OR3_X1 c6472(
.A1(net6810),
.A2(net6806),
.A3(net11204),
.ZN(net6815)
);

OR4_X4 c6473(
.A1(net6813),
.A2(net6800),
.A3(net11202),
.A4(net11204),
.ZN(net6816)
);

INV_X4 c6474(
.A(net6806),
.ZN(net6817)
);

INV_X1 c6475(
.A(net9583),
.ZN(net6818)
);

INV_X2 c6476(
.A(net4952),
.ZN(net6819)
);

INV_X8 c6477(
.A(net5911),
.ZN(net6820)
);

MUX2_X1 c6478(
.A(net5854),
.B(net4945),
.S(net3899),
.Z(net6821)
);

INV_X16 c6479(
.A(net4850),
.ZN(net6822)
);

INV_X32 c6480(
.A(net5937),
.ZN(net6823)
);

INV_X4 c6481(
.A(net4890),
.ZN(net6824)
);

INV_X1 c6482(
.A(net9584),
.ZN(net6825)
);

SDFFR_X1 c6483(
.D(net6812),
.RN(net5937),
.SE(net5808),
.SI(net3979),
.CK(clk),
.Q(net6827),
.QN(net6826)
);

INV_X2 c6484(
.A(net6760),
.ZN(net6828)
);

INV_X8 c6485(
.A(net10375),
.ZN(net6829)
);

INV_X16 c6486(
.A(net6819),
.ZN(net6830)
);

XOR2_X1 c6487(
.A(net6735),
.B(net6784),
.Z(net6831)
);

NOR2_X1 c6488(
.A1(net4910),
.A2(net5810),
.ZN(net6832)
);

INV_X32 c6489(
.A(net5925),
.ZN(net6833)
);

INV_X4 c6490(
.A(net6730),
.ZN(net6834)
);

INV_X1 c6491(
.A(net5913),
.ZN(net6835)
);

INV_X2 c6492(
.A(net6823),
.ZN(net6836)
);

INV_X8 c6493(
.A(net6831),
.ZN(net6837)
);

INV_X16 c6494(
.A(net6818),
.ZN(net6838)
);

INV_X32 c6495(
.A(net6822),
.ZN(net6839)
);

INV_X4 c6496(
.A(net6829),
.ZN(net6840)
);

OR2_X2 c6497(
.A1(net5786),
.A2(net5776),
.ZN(net6841)
);

INV_X1 c6498(
.A(net6820),
.ZN(net6842)
);

INV_X2 c6499(
.A(net6766),
.ZN(net6843)
);

NOR2_X4 c6500(
.A1(net4936),
.A2(net5879),
.ZN(net6844)
);

NOR2_X2 c6501(
.A1(net6841),
.A2(net5858),
.ZN(net6845)
);

OAI21_X4 c6502(
.A(net6741),
.B1(net6818),
.B2(net6816),
.ZN(net6846)
);

INV_X8 c6503(
.A(net6836),
.ZN(net6847)
);

INV_X16 c6504(
.A(net6825),
.ZN(net6848)
);

INV_X32 c6505(
.A(net6816),
.ZN(net6849)
);

MUX2_X2 c6506(
.A(net6793),
.B(net4919),
.S(net6833),
.Z(net6850)
);

XOR2_X2 c6507(
.A(net6828),
.B(net5786),
.Z(net6851)
);

INV_X4 c6508(
.A(net6773),
.ZN(net6852)
);

NAND3_X4 c6509(
.A1(net6834),
.A2(net6850),
.A3(net6846),
.ZN(net6853)
);

INV_X1 c6510(
.A(net6839),
.ZN(net6854)
);

XNOR2_X1 c6511(
.A(net3880),
.B(net4885),
.ZN(net6855)
);

INV_X2 c6512(
.A(net9767),
.ZN(net6856)
);

OR3_X4 c6513(
.A1(net6823),
.A2(net6841),
.A3(net6837),
.ZN(net6857)
);

OAI22_X2 c6514(
.A1(net6847),
.A2(net2951),
.B1(net5879),
.B2(net6848),
.ZN(net6858)
);

INV_X8 c6515(
.A(net6835),
.ZN(net6859)
);

OR2_X4 c6516(
.A1(net6853),
.A2(net6844),
.ZN(net6860)
);

INV_X16 c6517(
.A(net6821),
.ZN(net6861)
);

OR2_X1 c6518(
.A1(net997),
.A2(net10465),
.ZN(net6862)
);

INV_X32 c6519(
.A(net6834),
.ZN(net6863)
);

XNOR2_X2 c6520(
.A(net4805),
.B(net6848),
.ZN(net6864)
);

AND2_X4 c6521(
.A1(net4885),
.A2(net6836),
.ZN(net6865)
);

INV_X4 c6522(
.A(net10824),
.ZN(net6866)
);

INV_X1 c6523(
.A(net10328),
.ZN(net6867)
);

AND3_X2 c6524(
.A1(net6865),
.A2(net5861),
.A3(net6864),
.ZN(net6868)
);

INV_X2 c6525(
.A(net6856),
.ZN(net6869)
);

NOR3_X1 c6526(
.A1(net6733),
.A2(net4927),
.A3(net6866),
.ZN(net6870)
);

AND2_X1 c6527(
.A1(net6784),
.A2(net10624),
.ZN(net6871)
);

NAND2_X1 c6528(
.A1(net5855),
.A2(net6848),
.ZN(net6872)
);

NAND2_X2 c6529(
.A1(net6849),
.A2(net6843),
.ZN(net6873)
);

INV_X8 c6530(
.A(net10183),
.ZN(net6874)
);

NAND2_X4 c6531(
.A1(net6848),
.A2(net6866),
.ZN(net6875)
);

SDFFR_X2 c6532(
.D(net6874),
.RN(net6858),
.SE(net6873),
.SI(net2920),
.CK(clk),
.Q(net6877),
.QN(net6876)
);

AND2_X2 c6533(
.A1(net6873),
.A2(net11205),
.ZN(net6878)
);

INV_X16 c6534(
.A(net6827),
.ZN(net6879)
);

XOR2_X1 c6535(
.A(net6862),
.B(net6878),
.Z(net6880)
);

INV_X32 c6536(
.A(net6866),
.ZN(net6881)
);

NOR2_X1 c6537(
.A1(net6878),
.A2(net4850),
.ZN(net6882)
);

OR2_X2 c6538(
.A1(net6854),
.A2(net6880),
.ZN(net6883)
);

NOR2_X4 c6539(
.A1(net6870),
.A2(net6766),
.ZN(net6884)
);

OAI211_X4 c6540(
.A(net6871),
.B(net6877),
.C1(net6828),
.C2(net6883),
.ZN(net6885)
);

AOI221_X4 c6541(
.A(net6880),
.B1(net6836),
.B2(net6866),
.C1(net6876),
.C2(net6883),
.ZN(net6886)
);

OR3_X2 c6542(
.A1(net6863),
.A2(net5859),
.A3(net6884),
.ZN(net6887)
);

INV_X4 c6543(
.A(net9925),
.ZN(net6888)
);

AOI221_X2 c6544(
.A(net6886),
.B1(net6882),
.B2(net6831),
.C1(net6883),
.C2(net5934),
.ZN(net6889)
);

DFFRS_X2 c6545(
.D(net6887),
.RN(net4885),
.SN(net6844),
.CK(clk),
.Q(net6891),
.QN(net6890)
);

OAI21_X2 c6546(
.A(net6867),
.B1(net6890),
.B2(net6875),
.ZN(net6892)
);

OAI21_X1 c6547(
.A(net5849),
.B1(net6817),
.B2(net10466),
.ZN(net6893)
);

INV_X1 c6548(
.A(net9946),
.ZN(net6894)
);

NOR2_X2 c6549(
.A1(net5919),
.A2(net6879),
.ZN(net6895)
);

XOR2_X2 c6550(
.A(net6891),
.B(net6819),
.Z(net6896)
);

XNOR2_X1 c6551(
.A(net6882),
.B(net10640),
.ZN(net6897)
);

AOI21_X2 c6552(
.A(net6842),
.B1(net6865),
.B2(net6852),
.ZN(net6898)
);

CLKGATETST_X1 c6553(
.E(net6898),
.SE(net10554),
.CK(clk),
.GCK(net6899)
);

OR2_X4 c6554(
.A1(net6892),
.A2(net6899),
.ZN(net6900)
);

AOI221_X1 c6555(
.A(net6875),
.B1(net6894),
.B2(net6898),
.C1(net6852),
.C2(net6892),
.ZN(net6901)
);

OAI222_X2 c6556(
.A1(net6894),
.A2(net6848),
.B1(net6892),
.B2(net6900),
.C1(net6896),
.C2(net4933),
.ZN(net6902)
);

INV_X2 c6557(
.A(net5982),
.ZN(net6903)
);

INV_X8 c6558(
.A(net4838),
.ZN(net6904)
);

INV_X16 c6559(
.A(net11024),
.ZN(net6905)
);

INV_X32 c6560(
.A(net6838),
.ZN(net6906)
);

INV_X4 c6561(
.A(net10492),
.ZN(net6907)
);

OR2_X1 c6562(
.A1(net6748),
.A2(net6883),
.ZN(net6908)
);

XNOR2_X2 c6563(
.A(net6869),
.B(net6852),
.ZN(net6909)
);

AND2_X4 c6564(
.A1(net6895),
.A2(net4871),
.ZN(net6910)
);

AND2_X1 c6565(
.A1(net6872),
.A2(net6010),
.ZN(net6911)
);

INV_X1 c6566(
.A(net5998),
.ZN(net6912)
);

INV_X2 c6567(
.A(net9676),
.ZN(net6913)
);

NAND2_X1 c6568(
.A1(net5047),
.A2(net6913),
.ZN(net6914)
);

INV_X8 c6569(
.A(net11020),
.ZN(net6915)
);

INV_X16 c6570(
.A(net6912),
.ZN(net6916)
);

NAND2_X2 c6571(
.A1(net6903),
.A2(net6909),
.ZN(net6917)
);

INV_X32 c6572(
.A(net5879),
.ZN(net6918)
);

NAND2_X4 c6573(
.A1(net6918),
.A2(net10600),
.ZN(net6919)
);

AND2_X2 c6574(
.A1(net5866),
.A2(net3081),
.ZN(net6920)
);

AOI21_X1 c6575(
.A(net6920),
.B1(net6918),
.B2(net5050),
.ZN(net6921)
);

XOR2_X1 c6576(
.A(net6018),
.B(net6844),
.Z(net6922)
);

INV_X4 c6577(
.A(net5057),
.ZN(net6923)
);

AOI21_X4 c6578(
.A(net6921),
.B1(net6877),
.B2(net6904),
.ZN(net6924)
);

INV_X1 c6579(
.A(net9675),
.ZN(net6925)
);

AND3_X1 c6580(
.A1(net5050),
.A2(net6918),
.A3(net6824),
.ZN(net6926)
);

CLKGATETST_X2 c6581(
.E(net6908),
.SE(net10956),
.CK(clk),
.GCK(net6927)
);

NAND3_X1 c6582(
.A1(net2859),
.A2(net3920),
.A3(net6884),
.ZN(net6928)
);

INV_X2 c6583(
.A(net5989),
.ZN(net6929)
);

NOR2_X1 c6584(
.A1(net3956),
.A2(net6023),
.ZN(net6930)
);

OR2_X2 c6585(
.A1(net6873),
.A2(net6872),
.ZN(net6931)
);

INV_X8 c6586(
.A(net10038),
.ZN(net6932)
);

NOR2_X4 c6587(
.A1(net6884),
.A2(net3956),
.ZN(net6933)
);

NOR2_X2 c6588(
.A1(net6013),
.A2(net6930),
.ZN(net6934)
);

INV_X16 c6589(
.A(net9706),
.ZN(net6935)
);

INV_X32 c6590(
.A(net6916),
.ZN(net6936)
);

XOR2_X2 c6591(
.A(net5943),
.B(net6020),
.Z(net6937)
);

SDFF_X1 c6592(
.D(net5951),
.SE(net6883),
.SI(net5879),
.CK(clk),
.Q(net6939),
.QN(net6938)
);

XNOR2_X1 c6593(
.A(net6846),
.B(net6909),
.ZN(net6940)
);

OR2_X4 c6594(
.A1(net6939),
.A2(net6915),
.ZN(net6941)
);

NOR3_X4 c6595(
.A1(net5988),
.A2(net6900),
.A3(net2859),
.ZN(net6942)
);

INV_X4 c6596(
.A(net11129),
.ZN(net6943)
);

OR2_X1 c6597(
.A1(net6859),
.A2(net6936),
.ZN(net6944)
);

INV_X1 c6598(
.A(net6864),
.ZN(net6945)
);

NOR3_X2 c6599(
.A1(net6022),
.A2(net6911),
.A3(net6938),
.ZN(net6946)
);

AND3_X4 c6600(
.A1(net6937),
.A2(net6909),
.A3(net10956),
.ZN(net6947)
);

INV_X2 c6601(
.A(net9921),
.ZN(net6948)
);

NAND3_X2 c6602(
.A1(net6932),
.A2(net6013),
.A3(net6902),
.ZN(net6949)
);

XNOR2_X2 c6603(
.A(net6926),
.B(net10433),
.ZN(net6950)
);

AND2_X4 c6604(
.A1(net6897),
.A2(net6919),
.ZN(net6951)
);

SDFF_X2 c6605(
.D(net6911),
.SE(net6913),
.SI(net6945),
.CK(clk),
.Q(net6953),
.QN(net6952)
);

INV_X8 c6606(
.A(net6918),
.ZN(net6954)
);

INV_X16 c6607(
.A(net11054),
.ZN(net6955)
);

INV_X32 c6608(
.A(net9687),
.ZN(net6956)
);

AND2_X1 c6609(
.A1(net6944),
.A2(net6940),
.ZN(net6957)
);

NAND2_X1 c6610(
.A1(net6947),
.A2(net6955),
.ZN(net6958)
);

INV_X4 c6611(
.A(net6940),
.ZN(net6959)
);

OR3_X1 c6612(
.A1(net6727),
.A2(net6952),
.A3(net6955),
.ZN(net6960)
);

INV_X1 c6613(
.A(net6949),
.ZN(net6961)
);

NAND2_X2 c6614(
.A1(net6932),
.A2(net10635),
.ZN(net6962)
);

NAND2_X4 c6615(
.A1(net6906),
.A2(net6017),
.ZN(net6963)
);

MUX2_X1 c6616(
.A(net6961),
.B(net4032),
.S(net6930),
.Z(net6964)
);

INV_X2 c6617(
.A(net11020),
.ZN(net6965)
);

OAI21_X4 c6618(
.A(net6014),
.B1(net6939),
.B2(net5965),
.ZN(net6966)
);

MUX2_X2 c6619(
.A(net6960),
.B(net6940),
.S(net6955),
.Z(net6967)
);

AND2_X2 c6620(
.A1(net6910),
.A2(net6963),
.ZN(net6968)
);

XOR2_X1 c6621(
.A(net6958),
.B(net6879),
.Z(net6969)
);

NOR2_X1 c6622(
.A1(net6963),
.A2(net6949),
.ZN(net6970)
);

OR2_X2 c6623(
.A1(net6945),
.A2(net6018),
.ZN(net6971)
);

OAI211_X1 c6624(
.A(net6941),
.B(net6964),
.C1(net6860),
.C2(net6786),
.ZN(net6972)
);

INV_X8 c6625(
.A(net10059),
.ZN(net6973)
);

INV_X16 c6626(
.A(net10078),
.ZN(net6974)
);

NAND3_X4 c6627(
.A1(net6957),
.A2(net6960),
.A3(net6920),
.ZN(net6975)
);

INV_X32 c6628(
.A(net10039),
.ZN(net6976)
);

CLKGATETST_X4 c6629(
.E(net6968),
.SE(net6953),
.CK(clk),
.GCK(net6977)
);

INV_X4 c6630(
.A(net10198),
.ZN(net6978)
);

OR3_X4 c6631(
.A1(net6915),
.A2(net6977),
.A3(net5902),
.ZN(net6979)
);

AND3_X2 c6632(
.A1(net6934),
.A2(net6959),
.A3(net6966),
.ZN(net6980)
);

NOR2_X4 c6633(
.A1(net4980),
.A2(net6980),
.ZN(net6981)
);

INV_X1 c6634(
.A(net10000),
.ZN(net6982)
);

NOR3_X1 c6635(
.A1(net6974),
.A2(net6969),
.A3(net5899),
.ZN(net6983)
);

NOR2_X2 c6636(
.A1(net6982),
.A2(net6948),
.ZN(net6984)
);

DFFRS_X1 c6637(
.D(net6984),
.RN(net6950),
.SN(net6935),
.CK(clk),
.Q(net6986),
.QN(net6985)
);

XOR2_X2 c6638(
.A(net6959),
.B(net6986),
.Z(net6987)
);

AOI222_X1 c6639(
.A1(net6978),
.A2(net6975),
.B1(net6984),
.B2(net6985),
.C1(net6987),
.C2(net6927),
.ZN(net6988)
);

INV_X2 c6640(
.ZN(net6989)
);

XNOR2_X1 c6641(
.A(net6057),
.B(net6069),
.ZN(net6990)
);

OR2_X4 c6642(
.A1(net6925),
.A2(net6098),
.ZN(net6991)
);

OR2_X1 c6643(
.A1(net6052),
.A2(net6970),
.ZN(net6992)
);

XNOR2_X2 c6644(
.A(net6943),
.B(net11126),
.ZN(net6993)
);

AND2_X4 c6645(
.A1(net6024),
.A2(net6757),
.ZN(net6994)
);

AND2_X1 c6646(
.A1(net6089),
.A2(net6023),
.ZN(net6995)
);

NAND2_X1 c6647(
.A1(net5135),
.A2(net6902),
.ZN(net6996)
);

INV_X8 c6648(
.A(net11127),
.ZN(net6997)
);

NAND2_X2 c6649(
.A1(net5107),
.A2(net6046),
.ZN(net6998)
);

INV_X16 c6650(
.A(net6907),
.ZN(net6999)
);

CLKGATETST_X8 c6651(
.E(net6990),
.SE(net6029),
.CK(clk),
.GCK(net7000)
);

INV_X32 c6652(
.A(net3175),
.ZN(net7001)
);

NAND2_X4 c6653(
.A1(net6004),
.A2(net4141),
.ZN(net7002)
);

INV_X4 c6654(
.A(net9845),
.ZN(net7003)
);

OR3_X2 c6655(
.A1(net4985),
.A2(net6980),
.A3(net3134),
.ZN(net7004)
);

AND2_X2 c6656(
.A1(net6086),
.A2(net10921),
.ZN(net7005)
);

XOR2_X1 c6657(
.A(net6069),
.B(net6992),
.Z(net7006)
);

DFFRS_X2 c6658(
.D(net6861),
.RN(net6860),
.SN(net6023),
.CK(clk),
.Q(net7008),
.QN(net7007)
);

NOR2_X1 c6659(
.A1(net6999),
.A2(net6043),
.ZN(net7009)
);

OR2_X2 c6660(
.A1(net5079),
.A2(net6926),
.ZN(net7010)
);

NOR2_X4 c6661(
.A1(net6782),
.A2(net6905),
.ZN(net7011)
);

NOR2_X2 c6662(
.A1(net6028),
.A2(net11005),
.ZN(net7012)
);

XOR2_X2 c6663(
.A(net6860),
.B(net6726),
.Z(net7013)
);

INV_X1 c6664(
.A(net11127),
.ZN(net7014)
);

INV_X2 c6665(
.A(net9994),
.ZN(net7015)
);

OAI21_X2 c6666(
.A(net6905),
.B1(net7010),
.B2(net6943),
.ZN(net7016)
);

INV_X8 c6667(
.A(net10908),
.ZN(net7017)
);

INV_X16 c6668(
.A(net6060),
.ZN(net7018)
);

XNOR2_X1 c6669(
.A(net3180),
.B(net4099),
.ZN(net7019)
);

INV_X32 c6670(
.A(net11072),
.ZN(net7020)
);

OR2_X4 c6671(
.A1(net6980),
.A2(net5107),
.ZN(net7021)
);

OR2_X1 c6672(
.A1(net6860),
.A2(net10653),
.ZN(net7022)
);

XNOR2_X2 c6673(
.A(net6010),
.B(net6881),
.ZN(net7023)
);

AND2_X4 c6674(
.A1(net7003),
.A2(net7017),
.ZN(net7024)
);

AND2_X1 c6675(
.A1(net7014),
.A2(net6089),
.ZN(net7025)
);

NAND2_X1 c6676(
.A1(net6986),
.A2(net6038),
.ZN(net7026)
);

OAI21_X1 c6677(
.A(net6936),
.B1(net6991),
.B2(net7020),
.ZN(net7027)
);

NAND2_X2 c6678(
.A1(net5776),
.A2(net7010),
.ZN(net7028)
);

NAND2_X4 c6679(
.A1(net5995),
.A2(net6994),
.ZN(net7029)
);

AOI21_X2 c6680(
.A(net6031),
.B1(net6060),
.B2(net6933),
.ZN(net7030)
);

INV_X4 c6681(
.A(net9939),
.ZN(net7031)
);

AOI21_X1 c6682(
.A(net7018),
.B1(net6995),
.B2(net6985),
.ZN(net7032)
);

AND2_X2 c6683(
.A1(net6029),
.A2(net4985),
.ZN(net7033)
);

XOR2_X1 c6684(
.A(net5958),
.B(net6993),
.Z(net7034)
);

AOI21_X4 c6685(
.A(net7001),
.B1(net6905),
.B2(net10707),
.ZN(net7035)
);

INV_X1 c6686(
.A(net10116),
.ZN(net7036)
);

NOR2_X1 c6687(
.A1(net6935),
.A2(net979),
.ZN(net7037)
);

DFFR_X1 c6688(
.D(net6881),
.RN(net6964),
.CK(clk),
.Q(net7039),
.QN(net7038)
);

INV_X2 c6689(
.A(net9844),
.ZN(net7040)
);

OR2_X2 c6690(
.A1(net7031),
.A2(net7019),
.ZN(net7041)
);

SDFF_X1 c6691(
.D(net7040),
.SE(net7034),
.SI(net11197),
.CK(clk),
.Q(net7043),
.QN(net7042)
);

NOR2_X4 c6692(
.A1(net6922),
.A2(net6977),
.ZN(net7044)
);

NOR2_X2 c6693(
.A1(net7043),
.A2(net7000),
.ZN(net7045)
);

XOR2_X2 c6694(
.A(net7020),
.B(net10558),
.Z(net7046)
);

XNOR2_X1 c6695(
.A(net6923),
.B(net7044),
.ZN(net7047)
);

OR2_X4 c6696(
.A1(net7035),
.A2(net11082),
.ZN(net7048)
);

OR2_X1 c6697(
.A1(net7046),
.A2(net6996),
.ZN(net7049)
);

SDFFS_X1 c6698(
.D(net6054),
.SE(net7040),
.SI(net4141),
.SN(net5114),
.CK(clk),
.Q(net7051),
.QN(net7050)
);

XNOR2_X2 c6699(
.A(net7033),
.B(net7051),
.ZN(net7052)
);

AND2_X4 c6700(
.A1(net7045),
.A2(net10659),
.ZN(net7053)
);

AND3_X1 c6701(
.A1(net7037),
.A2(net6995),
.A3(net10634),
.ZN(net7054)
);

AND2_X1 c6702(
.A1(net6103),
.A2(net7035),
.ZN(net7055)
);

NAND2_X1 c6703(
.A1(net7009),
.A2(net6021),
.ZN(net7056)
);

NAND3_X1 c6704(
.A1(net6929),
.A2(net7052),
.A3(net7034),
.ZN(net7057)
);

NAND2_X2 c6705(
.A1(net6046),
.A2(net7029),
.ZN(net7058)
);

NAND2_X4 c6706(
.A1(net7050),
.A2(net10688),
.ZN(net7059)
);

AND2_X2 c6707(
.A1(net7058),
.A2(net4927),
.ZN(net7060)
);

XOR2_X1 c6708(
.A(net7059),
.B(net6089),
.Z(net7061)
);

NOR2_X1 c6709(
.A1(net6989),
.A2(net5142),
.ZN(net7062)
);

OR2_X2 c6710(
.A1(net5898),
.A2(net7056),
.ZN(net7063)
);

NOR4_X4 c6711(
.A1(net7027),
.A2(net7056),
.A3(net7035),
.A4(net6089),
.ZN(net7064)
);

NOR2_X4 c6712(
.A1(net7037),
.A2(net6989),
.ZN(net7065)
);

SDFF_X2 c6713(
.D(net7065),
.SE(net7019),
.SI(net7044),
.CK(clk),
.Q(net7067),
.QN(net7066)
);

NOR3_X4 c6714(
.A1(net6043),
.A2(net7008),
.A3(net11117),
.ZN(net7068)
);

NOR2_X2 c6715(
.A1(net4099),
.A2(net7035),
.ZN(net7069)
);

NOR3_X2 c6716(
.A1(net7045),
.A2(net7069),
.A3(net11117),
.ZN(net7070)
);

AND3_X4 c6717(
.A1(net7068),
.A2(net7036),
.A3(net10706),
.ZN(net7071)
);

XOR2_X2 c6718(
.A(net6998),
.B(net6986),
.Z(net7072)
);

XNOR2_X1 c6719(
.A(net5902),
.B(net7068),
.ZN(net7073)
);

NAND3_X2 c6720(
.A1(net7069),
.A2(net7054),
.A3(net7063),
.ZN(net7074)
);

AOI222_X4 c6721(
.A1(net7068),
.A2(net7042),
.B1(net6951),
.B2(net7035),
.C1(net5899),
.C2(net10559),
.ZN(net7075)
);

OR2_X4 c6722(
.A1(net7073),
.A2(net10780),
.ZN(net7076)
);

INV_X8 c6723(
.A(net7023),
.ZN(net7077)
);

INV_X16 c6724(
.A(net7076),
.ZN(net7078)
);

OR2_X1 c6725(
.A1(net7012),
.A2(net5211),
.ZN(net7079)
);

NOR4_X2 c6726(
.A1(net6956),
.A2(net6987),
.A3(net5211),
.A4(net6182),
.ZN(net7080)
);

XNOR2_X2 c6727(
.A(net7063),
.B(net6193),
.ZN(net7081)
);

INV_X32 c6728(
.A(net6977),
.ZN(net7082)
);

SDFFS_X2 c6729(
.D(net5994),
.SE(net5154),
.SI(net7081),
.SN(net11074),
.CK(clk),
.Q(net7084),
.QN(net7083)
);

DFFRS_X1 c6730(
.D(net6176),
.RN(net7052),
.SN(net6116),
.CK(clk),
.Q(net7086),
.QN(net7085)
);

AND2_X4 c6731(
.A1(net6141),
.A2(net6956),
.ZN(net7087)
);

AND2_X1 c6732(
.A1(net6970),
.A2(net6193),
.ZN(net7088)
);

INV_X4 c6733(
.A(net5175),
.ZN(net7089)
);

INV_X1 c6734(
.A(net10119),
.ZN(net7090)
);

NAND2_X1 c6735(
.A1(net5859),
.A2(net7081),
.ZN(net7091)
);

INV_X2 c6736(
.A(net7051),
.ZN(net7092)
);

NAND2_X2 c6737(
.A1(net6171),
.A2(net5113),
.ZN(net7093)
);

INV_X8 c6738(
.A(net7052),
.ZN(net7094)
);

INV_X16 c6739(
.A(net9558),
.ZN(net7095)
);

INV_X32 c6740(
.A(net10372),
.ZN(net7096)
);

NAND2_X4 c6741(
.A1(net7089),
.A2(net7007),
.ZN(net7097)
);

AND2_X2 c6742(
.A1(net5211),
.A2(net6177),
.ZN(net7098)
);

DFFR_X2 c6743(
.D(net7040),
.RN(net7081),
.CK(clk),
.Q(net7100),
.QN(net7099)
);

OR3_X1 c6744(
.A1(net7048),
.A2(net7084),
.A3(net5034),
.ZN(net7101)
);

XOR2_X1 c6745(
.A(net6902),
.B(net11191),
.Z(net7102)
);

INV_X4 c6746(
.A(net11097),
.ZN(net7103)
);

INV_X1 c6747(
.A(net9892),
.ZN(net7104)
);

NOR2_X1 c6748(
.A1(net6183),
.A2(net10928),
.ZN(net7105)
);

OR2_X2 c6749(
.A1(net6168),
.A2(net7084),
.ZN(net7106)
);

MUX2_X1 c6750(
.A(net7011),
.B(net6129),
.S(net7085),
.Z(net7107)
);

INV_X2 c6751(
.A(net7056),
.ZN(net7108)
);

NOR2_X4 c6752(
.A1(net7092),
.A2(net11153),
.ZN(net7109)
);

INV_X8 c6753(
.A(net10262),
.ZN(net7110)
);

INV_X16 c6754(
.A(net10319),
.ZN(net7111)
);

INV_X32 c6755(
.A(net7100),
.ZN(net7112)
);

NOR2_X2 c6756(
.A1(net7097),
.A2(net6141),
.ZN(net7113)
);

INV_X4 c6757(
.A(net6047),
.ZN(net7114)
);

XOR2_X2 c6758(
.A(net7008),
.B(net7108),
.Z(net7115)
);

INV_X1 c6759(
.A(net11035),
.ZN(net7116)
);

XNOR2_X1 c6760(
.A(net7114),
.B(net7107),
.ZN(net7117)
);

INV_X2 c6761(
.A(net7110),
.ZN(net7118)
);

OR2_X4 c6762(
.A1(net4190),
.A2(net1114),
.ZN(net7119)
);

INV_X8 c6763(
.A(net5923),
.ZN(net7120)
);

INV_X16 c6764(
.A(net7119),
.ZN(net7121)
);

INV_X32 c6765(
.A(net4222),
.ZN(net7122)
);

INV_X4 c6766(
.A(net7064),
.ZN(net7123)
);

OR2_X1 c6767(
.A1(net7105),
.A2(net7110),
.ZN(net7124)
);

DFFRS_X2 c6768(
.D(net7112),
.RN(net7108),
.SN(net7081),
.CK(clk),
.Q(net7126),
.QN(net7125)
);

XNOR2_X2 c6769(
.A(net6173),
.B(net3856),
.ZN(net7127)
);

AND2_X4 c6770(
.A1(net7111),
.A2(net6108),
.ZN(net7128)
);

AND2_X1 c6771(
.A1(net7117),
.A2(net6996),
.ZN(net7129)
);

NAND2_X1 c6772(
.A1(net6182),
.A2(net7039),
.ZN(net7130)
);

NAND2_X2 c6773(
.A1(net7127),
.A2(net6047),
.ZN(net7131)
);

OAI21_X4 c6774(
.A(net7103),
.B1(net6190),
.B2(net6977),
.ZN(net7132)
);

INV_X1 c6775(
.A(net5114),
.ZN(net7133)
);

INV_X2 c6776(
.A(net9558),
.ZN(net7134)
);

MUX2_X2 c6777(
.A(net7116),
.B(net7079),
.S(net7094),
.Z(net7135)
);

NAND3_X4 c6778(
.A1(net7128),
.A2(net7127),
.A3(net7063),
.ZN(net7136)
);

NAND2_X4 c6779(
.A1(net7133),
.A2(net6993),
.ZN(net7137)
);

AND2_X2 c6780(
.A1(net6970),
.A2(net10785),
.ZN(net7138)
);

XOR2_X1 c6781(
.A(net7077),
.B(net10507),
.Z(net7139)
);

NOR2_X1 c6782(
.A1(net6143),
.A2(net7133),
.ZN(net7140)
);

INV_X8 c6783(
.A(net9816),
.ZN(net7141)
);

INV_X16 c6784(
.A(net11021),
.ZN(net7142)
);

INV_X32 c6785(
.A(net7106),
.ZN(net7143)
);

OR2_X2 c6786(
.A1(net7121),
.A2(net5156),
.ZN(net7144)
);

SDFF_X1 c6787(
.D(net7113),
.SE(net7099),
.SI(net7079),
.CK(clk),
.Q(net7146),
.QN(net7145)
);

INV_X4 c6788(
.A(net9915),
.ZN(net7147)
);

INV_X1 c6789(
.A(net9771),
.ZN(net7148)
);

OR3_X4 c6790(
.A1(net7115),
.A2(net7138),
.A3(net5859),
.ZN(net7149)
);

NOR2_X4 c6791(
.A1(net7133),
.A2(net10570),
.ZN(net7150)
);

AND3_X2 c6792(
.A1(net7122),
.A2(net7129),
.A3(net5133),
.ZN(net7151)
);

NOR2_X2 c6793(
.A1(net7142),
.A2(net7077),
.ZN(net7152)
);

INV_X2 c6794(
.A(net10347),
.ZN(net7153)
);

SDFFRS_X1 c6795(
.D(net7136),
.RN(net7152),
.SE(net7142),
.SI(net7084),
.SN(net7081),
.CK(clk),
.Q(net7155),
.QN(net7154)
);

INV_X8 c6796(
.A(net9687),
.ZN(net7156)
);

OAI33_X1 c6797(
.A1(net7152),
.A2(net7151),
.A3(net7130),
.B1(net5848),
.B2(net5166),
.B3(net7081),
.ZN(net7157)
);

AOI211_X4 c6798(
.A(net6132),
.B(net7114),
.C1(net7133),
.C2(net11206),
.ZN(net7158)
);

XOR2_X2 c6799(
.A(net6157),
.B(net7140),
.Z(net7159)
);

NOR3_X1 c6800(
.A1(net7104),
.A2(net7156),
.A3(net7152),
.ZN(net7160)
);

XNOR2_X1 c6801(
.A(net7143),
.B(net7146),
.ZN(net7161)
);

OR3_X2 c6802(
.A1(net6191),
.A2(net7161),
.A3(net7159),
.ZN(net7162)
);

OAI21_X2 c6803(
.A(net7160),
.B1(net7154),
.B2(net7156),
.ZN(net7163)
);

OAI21_X1 c6804(
.A(net7124),
.B1(net7160),
.B2(net7126),
.ZN(net7164)
);

AOI222_X2 c6805(
.A1(net7148),
.A2(net7120),
.B1(net7164),
.B2(net7163),
.C1(net7125),
.C2(net7036),
.ZN(net7165)
);

INV_X16 c6806(
.A(net5944),
.ZN(net7166)
);

OR2_X4 c6807(
.A1(net6249),
.A2(net7147),
.ZN(net7167)
);

INV_X32 c6808(
.A(net4267),
.ZN(net7168)
);

INV_X4 c6809(
.A(net10079),
.ZN(net7169)
);

INV_X1 c6810(
.A(net9607),
.ZN(net7170)
);

OR2_X1 c6811(
.A1(net4307),
.A2(net7085),
.ZN(net7171)
);

XNOR2_X2 c6812(
.A(net6178),
.B(net5944),
.ZN(net7172)
);

INV_X2 c6813(
.A(net6266),
.ZN(net7173)
);

INV_X8 c6814(
.A(net6023),
.ZN(net7174)
);

INV_X16 c6815(
.A(net7173),
.ZN(net7175)
);

INV_X32 c6816(
.A(net6036),
.ZN(net7176)
);

AND2_X4 c6817(
.A1(net7174),
.A2(net6238),
.ZN(net7177)
);

INV_X4 c6818(
.A(net9606),
.ZN(net7178)
);

AOI21_X2 c6819(
.A(net7170),
.B1(net6210),
.B2(net6239),
.ZN(net7179)
);

INV_X1 c6820(
.A(net11059),
.ZN(net7180)
);

INV_X2 c6821(
.A(net7175),
.ZN(net7181)
);

INV_X8 c6822(
.A(net5245),
.ZN(net7182)
);

INV_X16 c6823(
.A(net7177),
.ZN(net7183)
);

INV_X32 c6824(
.A(net7146),
.ZN(net7184)
);

AOI21_X1 c6825(
.A(net3107),
.B1(net7171),
.B2(net6217),
.ZN(net7185)
);

INV_X4 c6826(
.A(net7093),
.ZN(net7186)
);

INV_X1 c6827(
.A(net7155),
.ZN(net7187)
);

AND2_X1 c6828(
.A1(net7168),
.A2(net7159),
.ZN(net7188)
);

INV_X2 c6829(
.A(net4338),
.ZN(net7189)
);

AOI21_X4 c6830(
.A(net7134),
.B1(net7080),
.B2(net7150),
.ZN(net7190)
);

INV_X8 c6831(
.A(net10302),
.ZN(net7191)
);

NAND2_X1 c6832(
.A1(net7180),
.A2(net6273),
.ZN(net7192)
);

INV_X16 c6833(
.A(net6265),
.ZN(net7193)
);

NAND2_X2 c6834(
.A1(net7156),
.A2(net7170),
.ZN(net7194)
);

NAND2_X4 c6835(
.A1(net7182),
.A2(net6265),
.ZN(net7195)
);

INV_X32 c6836(
.A(net7187),
.ZN(net7196)
);

AND2_X2 c6837(
.A1(net7107),
.A2(net6952),
.ZN(net7197)
);

INV_X4 c6838(
.A(net4025),
.ZN(net7198)
);

INV_X1 c6839(
.A(net6238),
.ZN(net7199)
);

INV_X2 c6840(
.A(net6232),
.ZN(net7200)
);

XOR2_X1 c6841(
.A(net7169),
.B(net11001),
.Z(net7201)
);

NOR2_X1 c6842(
.A1(net5288),
.A2(net7145),
.ZN(net7202)
);

INV_X8 c6843(
.A(net7167),
.ZN(net7203)
);

INV_X16 c6844(
.A(net3383),
.ZN(net7204)
);

OR2_X2 c6845(
.A1(net7204),
.A2(net7156),
.ZN(net7205)
);

INV_X32 c6846(
.A(net9827),
.ZN(net7206)
);

NOR2_X4 c6847(
.A1(net7130),
.A2(net6184),
.ZN(net7207)
);

NOR2_X2 c6848(
.A1(net7178),
.A2(net7177),
.ZN(net7208)
);

OAI221_X1 c6849(
.A(net5133),
.B1(net7155),
.B2(net7145),
.C1(net7083),
.C2(net7125),
.ZN(net7209)
);

XOR2_X2 c6850(
.A(net7080),
.B(net7126),
.Z(net7210)
);

SDFF_X2 c6851(
.D(net4302),
.SE(net6179),
.SI(net7186),
.CK(clk),
.Q(net7212),
.QN(net7211)
);

XNOR2_X1 c6852(
.A(net7188),
.B(net7177),
.ZN(net7213)
);

DFFRS_X1 c6853(
.D(net7086),
.RN(net6184),
.SN(net7185),
.CK(clk),
.Q(net7215),
.QN(net7214)
);

OR2_X4 c6854(
.A1(net7186),
.A2(net7200),
.ZN(net7216)
);

AND3_X1 c6855(
.A1(net7171),
.A2(net7081),
.A3(net7178),
.ZN(net7217)
);

INV_X4 c6856(
.A(net10507),
.ZN(net7218)
);

NAND3_X1 c6857(
.A1(net7209),
.A2(net6253),
.A3(net7189),
.ZN(net7219)
);

INV_X1 c6858(
.A(net7183),
.ZN(net7220)
);

OR2_X1 c6859(
.A1(net7083),
.A2(net11027),
.ZN(net7221)
);

XNOR2_X2 c6860(
.A(net5276),
.B(net7159),
.ZN(net7222)
);

AND2_X4 c6861(
.A1(net6993),
.A2(net6222),
.ZN(net7223)
);

AND2_X1 c6862(
.A1(net7206),
.A2(net4024),
.ZN(net7224)
);

OAI221_X4 c6863(
.A(net7184),
.B1(net5288),
.B2(net7221),
.C1(net7164),
.C2(net7125),
.ZN(net7225)
);

NOR3_X4 c6864(
.A1(net7044),
.A2(net7223),
.A3(net7199),
.ZN(net7226)
);

INV_X2 c6865(
.A(net9748),
.ZN(net7227)
);

NOR3_X2 c6866(
.A1(net7201),
.A2(net7130),
.A3(net6183),
.ZN(net7228)
);

AND3_X4 c6867(
.A1(net7223),
.A2(net7200),
.A3(net5245),
.ZN(net7229)
);

NAND2_X1 c6868(
.A1(net7218),
.A2(net10952),
.ZN(net7230)
);

NAND2_X2 c6869(
.A1(net7205),
.A2(net6987),
.ZN(net7231)
);

NAND2_X4 c6870(
.A1(net4336),
.A2(net6266),
.ZN(net7232)
);

AND2_X2 c6871(
.A1(net7223),
.A2(net10483),
.ZN(net7233)
);

XOR2_X1 c6872(
.A(net7197),
.B(net7231),
.Z(net7234)
);

NOR2_X1 c6873(
.A1(net7225),
.A2(net11098),
.ZN(net7235)
);

OR2_X2 c6874(
.A1(net7213),
.A2(net7208),
.ZN(net7236)
);

INV_X8 c6875(
.A(net10932),
.ZN(net7237)
);

NAND3_X2 c6876(
.A1(net7237),
.A2(net7036),
.A3(net7024),
.ZN(net7238)
);

OR3_X1 c6877(
.A1(net6275),
.A2(net7238),
.A3(net7175),
.ZN(net7239)
);

NOR2_X4 c6878(
.A1(net7230),
.A2(net7086),
.ZN(net7240)
);

INV_X16 c6879(
.A(net10835),
.ZN(net7241)
);

MUX2_X1 c6880(
.A(net7196),
.B(net7236),
.S(net7241),
.Z(net7242)
);

OAI21_X4 c6881(
.A(net6239),
.B1(net7238),
.B2(net7224),
.ZN(net7243)
);

NOR4_X1 c6882(
.A1(net7166),
.A2(net7233),
.A3(net7238),
.A4(net7224),
.ZN(net7244)
);

NOR2_X2 c6883(
.A1(net7228),
.A2(net7223),
.ZN(net7245)
);

MUX2_X2 c6884(
.A(net7245),
.B(net7232),
.S(net7243),
.Z(net7246)
);

AOI211_X2 c6885(
.A(net6953),
.B(net7189),
.C1(net7243),
.C2(net7223),
.ZN(net7247)
);

AOI22_X1 c6886(
.A1(net7240),
.A2(net7238),
.B1(net7243),
.B2(net7200),
.ZN(net7248)
);

OAI221_X2 c6887(
.A(net7247),
.B1(net7109),
.B2(net7238),
.C1(net6284),
.C2(net7208),
.ZN(net7249)
);

AOI221_X4 c6888(
.A(net7246),
.B1(net7024),
.B2(net7211),
.C1(net10547),
.C2(net11096),
.ZN(net7250)
);

XOR2_X2 c6889(
.A(net6098),
.B(net7164),
.Z(net7251)
);

XNOR2_X1 c6890(
.A(net5046),
.B(net6098),
.ZN(net7252)
);

OR2_X4 c6891(
.A1(net5331),
.A2(net5398),
.ZN(net7253)
);

OR2_X1 c6892(
.A1(net6350),
.A2(net2346),
.ZN(net7254)
);

INV_X32 c6893(
.A(net5994),
.ZN(net7255)
);

XNOR2_X2 c6894(
.A(net7191),
.B(net6305),
.ZN(net7256)
);

INV_X4 c6895(
.A(net6359),
.ZN(net7257)
);

AND2_X4 c6896(
.A1(net3471),
.A2(net7208),
.ZN(net7258)
);

AND2_X1 c6897(
.A1(net7159),
.A2(net7108),
.ZN(net7259)
);

NAND2_X1 c6898(
.A1(net6233),
.A2(net6273),
.ZN(net7260)
);

NAND2_X2 c6899(
.A1(net7258),
.A2(net7189),
.ZN(net7261)
);

NAND2_X4 c6900(
.A1(net6367),
.A2(net6359),
.ZN(net7262)
);

AND2_X2 c6901(
.A1(net6183),
.A2(net6226),
.ZN(net7263)
);

XOR2_X1 c6902(
.A(net7252),
.B(net6358),
.Z(net7264)
);

NOR2_X1 c6903(
.A1(net7229),
.A2(net7024),
.ZN(net7265)
);

NAND3_X4 c6904(
.A1(net7256),
.A2(net7246),
.A3(net6369),
.ZN(net7266)
);

OR2_X2 c6905(
.A1(net7222),
.A2(net7264),
.ZN(net7267)
);

INV_X1 c6906(
.A(net7259),
.ZN(net7268)
);

INV_X2 c6907(
.A(net10245),
.ZN(net7269)
);

NOR2_X4 c6908(
.A1(net7108),
.A2(net7256),
.ZN(net7270)
);

NOR2_X2 c6909(
.A1(net7024),
.A2(net7268),
.ZN(net7271)
);

INV_X8 c6910(
.A(net9666),
.ZN(net7272)
);

XOR2_X2 c6911(
.A(net7264),
.B(net7215),
.Z(net7273)
);

INV_X16 c6912(
.A(net11072),
.ZN(net7274)
);

XNOR2_X1 c6913(
.A(net7047),
.B(net11001),
.ZN(net7275)
);

OR2_X4 c6914(
.A1(net5398),
.A2(net6177),
.ZN(net7276)
);

OR2_X1 c6915(
.A1(net6305),
.A2(net6367),
.ZN(net7277)
);

OR3_X4 c6916(
.A1(net7150),
.A2(net6370),
.A3(net7264),
.ZN(net7278)
);

INV_X32 c6917(
.A(net9959),
.ZN(net7279)
);

XNOR2_X2 c6918(
.A(net7081),
.B(net6359),
.ZN(net7280)
);

AND2_X4 c6919(
.A1(net7255),
.A2(net6284),
.ZN(net7281)
);

AND2_X1 c6920(
.A1(net6302),
.A2(net7264),
.ZN(net7282)
);

INV_X4 c6921(
.A(net9801),
.ZN(net7283)
);

NAND2_X1 c6922(
.A1(net7274),
.A2(net10438),
.ZN(net7284)
);

NAND2_X2 c6923(
.A1(net6768),
.A2(net7274),
.ZN(net7285)
);

INV_X1 c6924(
.A(net10151),
.ZN(net7286)
);

NAND2_X4 c6925(
.A1(net6799),
.A2(net7270),
.ZN(net7287)
);

SDFFR_X1 c6926(
.D(net7273),
.RN(net7283),
.SE(net6288),
.SI(net6273),
.CK(clk),
.Q(net7289),
.QN(net7288)
);

AND2_X2 c6927(
.A1(net7277),
.A2(net6361),
.ZN(net7290)
);

XOR2_X1 c6928(
.A(net7286),
.B(net6359),
.Z(net7291)
);

AND3_X2 c6929(
.A1(net6344),
.A2(net7263),
.A3(net7284),
.ZN(net7292)
);

NOR2_X1 c6930(
.A1(net7261),
.A2(net7244),
.ZN(net7293)
);

OR2_X2 c6931(
.A1(net6315),
.A2(net7283),
.ZN(net7294)
);

NOR2_X4 c6932(
.A1(net6361),
.A2(net7199),
.ZN(net7295)
);

NOR2_X2 c6933(
.A1(net7279),
.A2(net7283),
.ZN(net7296)
);

INV_X2 c6934(
.A(net9822),
.ZN(net7297)
);

XOR2_X2 c6935(
.A(net7270),
.B(net7297),
.Z(net7298)
);

INV_X8 c6936(
.A(net11114),
.ZN(net7299)
);

XNOR2_X1 c6937(
.A(net7295),
.B(net7181),
.ZN(net7300)
);

OR2_X4 c6938(
.A1(net7215),
.A2(net7224),
.ZN(net7301)
);

INV_X16 c6939(
.A(net10310),
.ZN(net7302)
);

OAI222_X1 c6940(
.A1(net7296),
.A2(net7302),
.B1(net6326),
.B2(net6183),
.C1(net7268),
.C2(net5973),
.ZN(net7303)
);

OR2_X1 c6941(
.A1(net7299),
.A2(net7198),
.ZN(net7304)
);

INV_X32 c6942(
.A(net9855),
.ZN(net7305)
);

NOR3_X1 c6943(
.A1(net7287),
.A2(net7289),
.A3(net11104),
.ZN(net7306)
);

XNOR2_X2 c6944(
.A(net7306),
.B(net7302),
.ZN(net7307)
);

AND2_X4 c6945(
.A1(net7301),
.A2(net11001),
.ZN(net7308)
);

AND2_X1 c6946(
.A1(net5394),
.A2(net7264),
.ZN(net7309)
);

NAND2_X1 c6947(
.A1(net7198),
.A2(net7256),
.ZN(net7310)
);

INV_X4 c6948(
.A(net10840),
.ZN(net7311)
);

NAND2_X2 c6949(
.A1(net7285),
.A2(net7263),
.ZN(net7312)
);

NAND2_X4 c6950(
.A1(net7308),
.A2(net6098),
.ZN(net7313)
);

OR3_X2 c6951(
.A1(net7298),
.A2(net7301),
.A3(net7313),
.ZN(net7314)
);

DFFRS_X2 c6952(
.D(net5376),
.RN(net7312),
.SN(net7192),
.CK(clk),
.Q(net7316),
.QN(net7315)
);

INV_X1 c6953(
.A(net9665),
.ZN(net7317)
);

AND4_X4 c6954(
.A1(net7274),
.A2(net6222),
.A3(net6361),
.A4(net7275),
.ZN(net7318)
);

AOI221_X2 c6955(
.A(net7296),
.B1(net7312),
.B2(net7268),
.C1(net7317),
.C2(net11104),
.ZN(net7319)
);

AND2_X2 c6956(
.A1(net7292),
.A2(net7315),
.ZN(net7320)
);

XOR2_X1 c6957(
.A(net7283),
.B(net7314),
.Z(net7321)
);

OAI21_X2 c6958(
.A(net7216),
.B1(net6283),
.B2(net7319),
.ZN(net7322)
);

SDFF_X1 c6959(
.D(net7276),
.SE(net7275),
.SI(net7306),
.CK(clk),
.Q(net7324),
.QN(net7323)
);

SDFF_X2 c6960(
.D(net7319),
.SE(net7323),
.SI(net5283),
.CK(clk),
.Q(net7326),
.QN(net7325)
);

OAI222_X4 c6961(
.A1(net7320),
.A2(net7310),
.B1(net7319),
.B2(net5283),
.C1(net7325),
.C2(net7081),
.ZN(net7327)
);

OAI21_X1 c6962(
.A(net5113),
.B1(net7313),
.B2(net11131),
.ZN(net7328)
);

AOI21_X2 c6963(
.A(net5340),
.B1(net7297),
.B2(net11131),
.ZN(net7329)
);

AOI21_X1 c6964(
.A(net7329),
.B1(net7311),
.B2(net7318),
.ZN(net7330)
);

AOI21_X4 c6965(
.A(net7316),
.B1(net7319),
.B2(net7211),
.ZN(net7331)
);

AND3_X1 c6966(
.A1(net7293),
.A2(net7246),
.A3(net7317),
.ZN(net7332)
);

NAND3_X1 c6967(
.A1(net7287),
.A2(net7272),
.A3(net11131),
.ZN(net7333)
);

NOR3_X4 c6968(
.A1(net7318),
.A2(net7324),
.A3(net7333),
.ZN(net7334)
);

NAND4_X1 c6969(
.A1(net7267),
.A2(net7313),
.A3(net7268),
.A4(net10838),
.ZN(net7335)
);

OAI222_X2 c6970(
.A1(net4350),
.A2(net7324),
.B1(net5156),
.B2(net7256),
.C1(net7325),
.C2(net7288),
.ZN(net7336)
);

OR4_X1 c6971(
.A1(net7297),
.A2(net7303),
.A3(net5325),
.A4(net6316),
.ZN(net7337)
);

DFFRS_X1 c6972(
.D(net4520),
.RN(net6284),
.SN(net6927),
.CK(clk),
.Q(net7339),
.QN(net7338)
);

NOR3_X2 c6973(
.A1(net7290),
.A2(net3536),
.A3(net7101),
.ZN(net7340)
);

NOR2_X1 c6974(
.A1(net6387),
.A2(net5112),
.ZN(net7341)
);

INV_X2 c6975(
.A(net6439),
.ZN(net7342)
);

INV_X8 c6976(
.A(net7172),
.ZN(net7343)
);

INV_X16 c6977(
.A(net9594),
.ZN(net7344)
);

INV_X32 c6978(
.A(net9594),
.ZN(net7345)
);

INV_X4 c6979(
.A(net10087),
.ZN(net7346)
);

OR2_X2 c6980(
.A1(net3498),
.A2(net7181),
.ZN(net7347)
);

INV_X1 c6981(
.A(net7047),
.ZN(net7348)
);

NOR2_X4 c6982(
.A1(net7192),
.A2(net11083),
.ZN(net7349)
);

INV_X2 c6983(
.A(net11083),
.ZN(net7350)
);

DFFRS_X2 c6984(
.D(net6177),
.RN(net7158),
.SN(net6460),
.CK(clk),
.Q(net7352),
.QN(net7351)
);

INV_X8 c6985(
.A(net9810),
.ZN(net7353)
);

INV_X16 c6986(
.A(net9850),
.ZN(net7354)
);

SDFF_X1 c6987(
.D(net7158),
.SE(net6395),
.SI(net5973),
.CK(clk),
.Q(net7356),
.QN(net7355)
);

INV_X32 c6988(
.A(net10162),
.ZN(net7357)
);

INV_X4 c6989(
.A(net11021),
.ZN(net7358)
);

NOR2_X2 c6990(
.A1(net6297),
.A2(net7346),
.ZN(net7359)
);

XOR2_X2 c6991(
.A(net6399),
.B(net7355),
.Z(net7360)
);

INV_X1 c6992(
.A(net7227),
.ZN(net7361)
);

INV_X2 c6993(
.A(net11102),
.ZN(net7362)
);

INV_X8 c6994(
.A(net6418),
.ZN(net7363)
);

XNOR2_X1 c6995(
.A(net7300),
.B(net6225),
.ZN(net7364)
);

OR2_X4 c6996(
.A1(net6329),
.A2(net7345),
.ZN(net7365)
);

INV_X16 c6997(
.A(net7304),
.ZN(net7366)
);

OR2_X1 c6998(
.A1(net7365),
.A2(net5481),
.ZN(net7367)
);

XNOR2_X2 c6999(
.A(net5320),
.B(net7359),
.ZN(net7368)
);

AND2_X4 c7000(
.A1(net7350),
.A2(net6413),
.ZN(net7369)
);

AND3_X4 c7001(
.A1(net6454),
.A2(net7369),
.A3(net7131),
.ZN(net7370)
);

AND2_X1 c7002(
.A1(net7195),
.A2(net7345),
.ZN(net7371)
);

NAND2_X1 c7003(
.A1(net7368),
.A2(net6438),
.ZN(net7372)
);

NAND2_X2 c7004(
.A1(net6328),
.A2(net7364),
.ZN(net7373)
);

INV_X32 c7005(
.A(net9702),
.ZN(net7374)
);

INV_X4 c7006(
.A(net9975),
.ZN(net7375)
);

NAND2_X4 c7007(
.A1(net6442),
.A2(net7354),
.ZN(net7376)
);

AND2_X2 c7008(
.A1(net7373),
.A2(net7355),
.ZN(net7377)
);

NAND3_X2 c7009(
.A1(net7374),
.A2(net7287),
.A3(net7376),
.ZN(net7378)
);

INV_X1 c7010(
.A(net6354),
.ZN(net7379)
);

XOR2_X1 c7011(
.A(net7101),
.B(net7227),
.Z(net7380)
);

NOR2_X1 c7012(
.A1(net7265),
.A2(net7357),
.ZN(net7381)
);

OR2_X2 c7013(
.A1(net7375),
.A2(net6405),
.ZN(net7382)
);

DFFS_X1 c7014(
.D(net7225),
.SN(net7275),
.CK(clk),
.Q(net7384),
.QN(net7383)
);

NOR2_X4 c7015(
.A1(net7272),
.A2(net7351),
.ZN(net7385)
);

OR3_X1 c7016(
.A1(net7385),
.A2(net7370),
.A3(net5320),
.ZN(net7386)
);

MUX2_X1 c7017(
.A(net7358),
.B(net7386),
.S(net7360),
.Z(net7387)
);

INV_X2 c7018(
.A(net9836),
.ZN(net7388)
);

NOR2_X2 c7019(
.A1(net1542),
.A2(net6217),
.ZN(net7389)
);

OAI21_X4 c7020(
.A(net7384),
.B1(net7374),
.B2(net5320),
.ZN(net7390)
);

XOR2_X2 c7021(
.A(net7380),
.B(net6426),
.Z(net7391)
);

INV_X8 c7022(
.A(net9811),
.ZN(net7392)
);

XNOR2_X1 c7023(
.A(net7381),
.B(net6395),
.ZN(net7393)
);

DFFS_X2 c7024(
.D(net7257),
.SN(net7383),
.CK(clk),
.Q(net7395),
.QN(net7394)
);

MUX2_X2 c7025(
.A(net6434),
.B(net7389),
.S(net7391),
.Z(net7396)
);

OR2_X4 c7026(
.A1(net6354),
.A2(net11093),
.ZN(net7397)
);

OR2_X1 c7027(
.A1(net5113),
.A2(net4261),
.ZN(net7398)
);

XNOR2_X2 c7028(
.A(net4479),
.B(net7387),
.ZN(net7399)
);

SDFF_X2 c7029(
.D(net7397),
.SE(net7356),
.SI(net7363),
.CK(clk),
.Q(net7401),
.QN(net7400)
);

INV_X16 c7030(
.A(net10883),
.ZN(net7402)
);

AND2_X4 c7031(
.A1(net7402),
.A2(net7357),
.ZN(net7403)
);

INV_X32 c7032(
.A(net7345),
.ZN(net7404)
);

AOI222_X1 c7033(
.A1(net7386),
.A2(net7153),
.B1(net6354),
.B2(net7275),
.C1(net7325),
.C2(net7357),
.ZN(net7405)
);

AND2_X1 c7034(
.A1(net7403),
.A2(net7391),
.ZN(net7406)
);

NAND2_X1 c7035(
.A1(net6412),
.A2(net7386),
.ZN(net7407)
);

NAND3_X4 c7036(
.A1(net7382),
.A2(net7352),
.A3(net11083),
.ZN(net7408)
);

NAND2_X2 c7037(
.A1(net7390),
.A2(net6329),
.ZN(net7409)
);

OR3_X4 c7038(
.A1(net2569),
.A2(net6405),
.A3(net7352),
.ZN(net7410)
);

NAND2_X4 c7039(
.A1(net7409),
.A2(net6414),
.ZN(net7411)
);

AND2_X2 c7040(
.A1(net7392),
.A2(net7158),
.ZN(net7412)
);

AND3_X2 c7041(
.A1(net7301),
.A2(net5320),
.A3(net6399),
.ZN(net7413)
);

XOR2_X1 c7042(
.A(net7398),
.B(net7408),
.Z(net7414)
);

NOR2_X1 c7043(
.A1(net7412),
.A2(net7411),
.ZN(net7415)
);

OR2_X2 c7044(
.A1(net7153),
.A2(net5469),
.ZN(net7416)
);

NOR3_X1 c7045(
.A1(net3397),
.A2(net7268),
.A3(net7369),
.ZN(net7417)
);

NOR2_X4 c7046(
.A1(net7404),
.A2(net7409),
.ZN(net7418)
);

INV_X4 c7047(
.A(net10045),
.ZN(net7419)
);

NOR2_X2 c7048(
.A1(net7408),
.A2(net7398),
.ZN(net7420)
);

INV_X1 c7049(
.A(net10021),
.ZN(net7421)
);

INV_X2 c7050(
.A(net11094),
.ZN(net7422)
);

DFFRS_X1 c7051(
.D(net7414),
.RN(net7399),
.SN(net7389),
.CK(clk),
.Q(net7424),
.QN(net7423)
);

DFFRS_X2 c7052(
.D(net3536),
.RN(net7153),
.SN(net7363),
.CK(clk),
.Q(net7426),
.QN(net7425)
);

OR3_X2 c7053(
.A1(net7422),
.A2(net7419),
.A3(net7425),
.ZN(net7427)
);

OAI21_X2 c7054(
.A(net7427),
.B1(net7397),
.B2(net7423),
.ZN(net7428)
);

INV_X8 c7055(
.A(net9909),
.ZN(net7429)
);

XOR2_X2 c7056(
.A(net2553),
.B(net5544),
.Z(net7430)
);

XNOR2_X1 c7057(
.A(net7289),
.B(net4588),
.ZN(net7431)
);

INV_X16 c7058(
.A(net9554),
.ZN(net7432)
);

OR2_X4 c7059(
.A1(net3594),
.A2(net6388),
.ZN(net7433)
);

INV_X32 c7060(
.A(net9835),
.ZN(net7434)
);

INV_X4 c7061(
.A(net9903),
.ZN(net7435)
);

OAI22_X1 c7062(
.A1(net7430),
.A2(net7387),
.B1(net7109),
.B2(net5474),
.ZN(net7436)
);

OR2_X1 c7063(
.A1(net6509),
.A2(net6533),
.ZN(net7437)
);

SDFF_X1 c7064(
.D(net5555),
.SE(net6509),
.SI(net7344),
.CK(clk),
.Q(net7439),
.QN(net7438)
);

XNOR2_X2 c7065(
.A(net6527),
.B(net7289),
.ZN(net7440)
);

AND2_X4 c7066(
.A1(net7415),
.A2(net5568),
.ZN(net7441)
);

AND2_X1 c7067(
.A1(net7391),
.A2(net7338),
.ZN(net7442)
);

SDFF_X2 c7068(
.D(net4548),
.SE(net7431),
.SI(net6467),
.CK(clk),
.Q(net7444),
.QN(net7443)
);

INV_X1 c7069(
.A(net9898),
.ZN(net7445)
);

INV_X2 c7070(
.A(out0),
.ZN(net7446)
);

NAND2_X1 c7071(
.A1(net1617),
.A2(net7443),
.ZN(net7447)
);

NAND2_X2 c7072(
.A1(net4588),
.A2(net6316),
.ZN(net7448)
);

INV_X8 c7073(
.A(net11057),
.ZN(net7449)
);

NAND2_X4 c7074(
.A1(net6508),
.A2(net7372),
.ZN(net7450)
);

AND2_X2 c7075(
.A1(net7376),
.A2(net7179),
.ZN(net7451)
);

SDFFRS_X2 c7076(
.D(net6511),
.RN(net4479),
.SE(net6444),
.SI(net6133),
.SN(net3576),
.CK(clk),
.Q(net7453),
.QN(net7452)
);

SDFFR_X2 c7077(
.D(net7446),
.RN(net6477),
.SE(net5555),
.SI(net7447),
.CK(clk),
.Q(net7455),
.QN(net7454)
);

XOR2_X1 c7078(
.A(net7362),
.B(net7367),
.Z(net7456)
);

OAI21_X1 c7079(
.A(net7434),
.B1(net7438),
.B2(net7367),
.ZN(net7457)
);

INV_X16 c7080(
.A(net9837),
.ZN(net7458)
);

NOR2_X1 c7081(
.A1(net630),
.A2(net7376),
.ZN(net7459)
);

OR2_X2 c7082(
.A1(net6485),
.A2(net7289),
.ZN(net7460)
);

NOR2_X4 c7083(
.A1(net5451),
.A2(net7382),
.ZN(net7461)
);

NOR2_X2 c7084(
.A1(net7313),
.A2(net7179),
.ZN(net7462)
);

INV_X32 c7085(
.A(net10032),
.ZN(net7463)
);

XOR2_X2 c7086(
.A(net7179),
.B(net7313),
.Z(net7464)
);

AOI21_X2 c7087(
.A(net5569),
.B1(net6467),
.B2(net7445),
.ZN(net7465)
);

AND4_X2 c7088(
.A1(net6505),
.A2(net1709),
.A3(net7452),
.A4(net7447),
.ZN(net7466)
);

INV_X4 c7089(
.A(net10361),
.ZN(net7467)
);

AOI222_X4 c7090(
.A1(net5482),
.A2(net7455),
.B1(net6485),
.B2(net6529),
.C1(net7458),
.C2(net6527),
.ZN(net7468)
);

AOI21_X1 c7091(
.A(net7441),
.B1(net5451),
.B2(net7434),
.ZN(net7469)
);

XNOR2_X1 c7092(
.A(net7464),
.B(net7326),
.ZN(net7470)
);

OR2_X4 c7093(
.A1(net7382),
.A2(net7430),
.ZN(net7471)
);

OR2_X1 c7094(
.A1(net6514),
.A2(net7454),
.ZN(net7472)
);

INV_X1 c7095(
.A(net10329),
.ZN(net7473)
);

XNOR2_X2 c7096(
.A(net7465),
.B(net7413),
.ZN(net7474)
);

AND2_X4 c7097(
.A1(net7366),
.A2(net6529),
.ZN(net7475)
);

INV_X2 c7098(
.A(net10033),
.ZN(net7476)
);

AND2_X1 c7099(
.A1(net7449),
.A2(net7465),
.ZN(net7477)
);

INV_X8 c7100(
.A(net11059),
.ZN(net7478)
);

DFFRS_X1 c7101(
.D(net6544),
.RN(net7462),
.SN(net7472),
.CK(clk),
.Q(net7480),
.QN(net7479)
);

NAND2_X1 c7102(
.A1(net5481),
.A2(net7462),
.ZN(net7481)
);

NAND2_X2 c7103(
.A1(net7460),
.A2(net7471),
.ZN(net7482)
);

NAND2_X4 c7104(
.A1(net7476),
.A2(net7481),
.ZN(net7483)
);

AND2_X2 c7105(
.A1(net7440),
.A2(net7482),
.ZN(net7484)
);

XOR2_X1 c7106(
.A(net6529),
.B(net7416),
.Z(net7485)
);

NOR2_X1 c7107(
.A1(net7484),
.A2(net7483),
.ZN(net7486)
);

AOI21_X4 c7108(
.A(net7479),
.B1(net6472),
.B2(net10736),
.ZN(net7487)
);

OR2_X2 c7109(
.A1(net7462),
.A2(net7477),
.ZN(net7488)
);

NOR2_X4 c7110(
.A1(net6466),
.A2(net7478),
.ZN(net7489)
);

NOR2_X2 c7111(
.A1(net7485),
.A2(net10428),
.ZN(net7490)
);

XOR2_X2 c7112(
.A(net7477),
.B(net7357),
.Z(net7491)
);

XNOR2_X1 c7113(
.A(net7482),
.B(net7480),
.ZN(net7492)
);

OR2_X4 c7114(
.A1(net7487),
.A2(net6529),
.ZN(net7493)
);

OR2_X1 c7115(
.A1(net7388),
.A2(net7457),
.ZN(net7494)
);

AND4_X1 c7116(
.A1(net7439),
.A2(net7489),
.A3(net4540),
.A4(net7325),
.ZN(net7495)
);

AND3_X1 c7117(
.A1(net7369),
.A2(net6405),
.A3(net7471),
.ZN(net7496)
);

XNOR2_X2 c7118(
.A(net699),
.B(net7333),
.ZN(net7497)
);

AND2_X4 c7119(
.A1(net7459),
.A2(net7478),
.ZN(net7498)
);

NAND3_X1 c7120(
.A1(net7497),
.A2(net7465),
.A3(net7493),
.ZN(net7499)
);

DFFRS_X2 c7121(
.D(net4471),
.RN(net7462),
.SN(net7499),
.CK(clk),
.Q(net7501),
.QN(net7500)
);

NOR3_X4 c7122(
.A1(net7488),
.A2(out25),
.A3(net7487),
.ZN(net7502)
);

AND2_X1 c7123(
.A1(net7287),
.A2(net4534),
.ZN(net7503)
);

NOR3_X2 c7124(
.A1(net7496),
.A2(net7501),
.A3(net7494),
.ZN(net7504)
);

NAND2_X1 c7125(
.A1(net7491),
.A2(net7478),
.ZN(net7505)
);

AND3_X4 c7126(
.A1(net7307),
.A2(net7492),
.A3(net7497),
.ZN(net7506)
);

NAND2_X2 c7127(
.A1(net7505),
.A2(net7504),
.ZN(net7507)
);

NAND3_X2 c7128(
.A1(net7185),
.A2(net7507),
.A3(net7497),
.ZN(net7508)
);

OR3_X1 c7129(
.A1(net7493),
.A2(net7484),
.A3(net7497),
.ZN(net7509)
);

MUX2_X1 c7130(
.A(net7343),
.B(net7430),
.S(net7418),
.Z(net7510)
);

SDFF_X1 c7131(
.D(net7506),
.SE(net7487),
.SI(net6452),
.CK(clk),
.Q(net7512),
.QN(net7511)
);

OAI21_X4 c7132(
.A(net7498),
.B1(net7441),
.B2(net7510),
.ZN(net7513)
);

AOI22_X4 c7133(
.A1(net7435),
.A2(net7447),
.B1(net5451),
.B2(net4460),
.ZN(net7514)
);

SDFF_X2 c7134(
.D(net7510),
.SE(net7505),
.SI(net7511),
.CK(clk),
.Q(net7516),
.QN(net7515)
);

OAI33_X1 c7135(
.A1(net7485),
.A2(net7512),
.A3(net7487),
.B1(net6529),
.B2(net7489),
.B3(net7490),
.ZN(net7517)
);

MUX2_X2 c7136(
.A(net10754),
.B(net11050),
.S(net11211),
.Z(net7518)
);

INV_X16 c7137(
.A(net9553),
.ZN(net7519)
);

NAND2_X4 c7138(
.A1(net7253),
.A2(net6612),
.ZN(net7520)
);

AND2_X2 c7139(
.A1(net7437),
.A2(net6487),
.ZN(net7521)
);

XOR2_X1 c7140(
.A(net6567),
.B(net7181),
.Z(net7522)
);

NOR2_X1 c7141(
.A1(net7516),
.A2(net3698),
.ZN(net7523)
);

OR2_X2 c7142(
.A1(net2737),
.A2(net7495),
.ZN(net7524)
);

NOR2_X4 c7143(
.A1(net7432),
.A2(net6629),
.ZN(net7525)
);

INV_X32 c7144(
.A(net9716),
.ZN(net7526)
);

NOR2_X2 c7145(
.A1(net4261),
.A2(net6612),
.ZN(net7527)
);

XOR2_X2 c7146(
.A(net6606),
.B(net6586),
.Z(net7528)
);

INV_X4 c7147(
.A(net9562),
.ZN(net7529)
);

XNOR2_X1 c7148(
.A(net6487),
.B(net7458),
.ZN(net7530)
);

OR2_X4 c7149(
.A1(net7450),
.A2(net7503),
.ZN(net7531)
);

OR2_X1 c7150(
.A1(net6614),
.A2(net7527),
.ZN(net7532)
);

XNOR2_X2 c7151(
.A(net7495),
.B(net7515),
.ZN(net7533)
);

AND2_X4 c7152(
.A1(net7522),
.A2(net7526),
.ZN(net7534)
);

NAND3_X4 c7153(
.A1(net4665),
.A2(net5973),
.A3(net11211),
.ZN(net7535)
);

OR3_X4 c7154(
.A1(net7527),
.A2(net7360),
.A3(net3691),
.ZN(net7536)
);

AND2_X1 c7155(
.A1(net7418),
.A2(net4678),
.ZN(net7537)
);

AOI221_X1 c7156(
.A(net2712),
.B1(net5630),
.B2(net2674),
.C1(net6607),
.C2(net3640),
.ZN(net7538)
);

NAND2_X1 c7157(
.A1(net6572),
.A2(net6467),
.ZN(net7539)
);

NAND2_X2 c7158(
.A1(net5617),
.A2(net708),
.ZN(net7540)
);

NAND2_X4 c7159(
.A1(net4678),
.A2(net7527),
.ZN(net7541)
);

AND2_X2 c7160(
.A1(net6616),
.A2(net6487),
.ZN(net7542)
);

INV_X1 c7161(
.A(net9561),
.ZN(net7543)
);

XOR2_X1 c7162(
.A(net4461),
.B(net4640),
.Z(net7544)
);

NOR2_X1 c7163(
.A1(net6578),
.A2(net7521),
.ZN(net7545)
);

OR2_X2 c7164(
.A1(net7526),
.A2(net7530),
.ZN(net7546)
);

NOR2_X4 c7165(
.A1(net7532),
.A2(net7527),
.ZN(net7547)
);

NOR2_X2 c7166(
.A1(net7339),
.A2(net7521),
.ZN(net7548)
);

XOR2_X2 c7167(
.A(net7444),
.B(net5617),
.Z(net7549)
);

INV_X2 c7168(
.A(net9851),
.ZN(net7550)
);

XNOR2_X1 c7169(
.A(net7521),
.B(net3691),
.ZN(net7551)
);

AND3_X2 c7170(
.A1(net7481),
.A2(net7432),
.A3(net11210),
.ZN(net7552)
);

OR2_X4 c7171(
.A1(net7547),
.A2(net7450),
.ZN(net7553)
);

NOR3_X1 c7172(
.A1(net5622),
.A2(net4665),
.A3(net7520),
.ZN(net7554)
);

OR3_X2 c7173(
.A1(net7407),
.A2(net7533),
.A3(net7521),
.ZN(net7555)
);

OAI21_X2 c7174(
.A(net7533),
.B1(net7418),
.B2(net7400),
.ZN(net7556)
);

OR2_X1 c7175(
.A1(net7548),
.A2(net6607),
.ZN(net7557)
);

OAI21_X1 c7176(
.A(net7544),
.B1(net7533),
.B2(net5634),
.ZN(net7558)
);

XNOR2_X2 c7177(
.A(net7524),
.B(net7489),
.ZN(net7559)
);

DFFRS_X1 c7178(
.D(net7534),
.RN(net7552),
.SN(net5667),
.CK(clk),
.Q(net7561),
.QN(net7560)
);

DFFRS_X2 c7179(
.D(net6628),
.RN(net6572),
.SN(net6607),
.CK(clk),
.Q(net7563),
.QN(net7562)
);

AND2_X4 c7180(
.A1(net7551),
.A2(net10494),
.ZN(net7564)
);

AOI21_X2 c7181(
.A(net7401),
.B1(net5574),
.B2(net6476),
.ZN(net7565)
);

SDFF_X1 c7182(
.D(net6488),
.SE(net7548),
.SI(net5604),
.CK(clk),
.Q(net7567),
.QN(net7566)
);

AOI21_X1 c7183(
.A(net7565),
.B1(net7560),
.B2(net11062),
.ZN(net7568)
);

INV_X8 c7184(
.A(net10181),
.ZN(net7569)
);

AOI21_X4 c7185(
.A(net7531),
.B1(net7471),
.B2(net6487),
.ZN(net7570)
);

AND2_X1 c7186(
.A1(net7541),
.A2(net7528),
.ZN(net7571)
);

AND3_X1 c7187(
.A1(net6550),
.A2(net7566),
.A3(net7552),
.ZN(net7572)
);

NAND3_X1 c7188(
.A1(net6549),
.A2(net7567),
.A3(net7542),
.ZN(net7573)
);

NAND2_X1 c7189(
.A1(net4656),
.A2(net7560),
.ZN(net7574)
);

NOR3_X4 c7190(
.A1(net7551),
.A2(net7574),
.A3(net5597),
.ZN(net7575)
);

NAND2_X2 c7191(
.A1(net7451),
.A2(net7523),
.ZN(net7576)
);

NOR3_X2 c7192(
.A1(net7567),
.A2(net6554),
.A3(net7562),
.ZN(net7577)
);

NAND2_X4 c7193(
.A1(net7577),
.A2(net7536),
.ZN(net7578)
);

AND2_X2 c7194(
.A1(net7564),
.A2(net7543),
.ZN(net7579)
);

OAI221_X1 c7195(
.A(net7535),
.B1(net7520),
.B2(net7490),
.C1(net4677),
.C2(net7545),
.ZN(net7580)
);

SDFF_X2 c7196(
.D(net5515),
.SE(net7574),
.SI(net7490),
.CK(clk),
.Q(net7582),
.QN(net7581)
);

XOR2_X1 c7197(
.A(net7569),
.B(net7571),
.Z(net7583)
);

AND3_X4 c7198(
.A1(net7583),
.A2(net7489),
.A3(net10641),
.ZN(net7584)
);

NAND3_X2 c7199(
.A1(net7542),
.A2(net7528),
.A3(net6600),
.ZN(net7585)
);

NOR2_X1 c7200(
.A1(net7556),
.A2(net7578),
.ZN(net7586)
);

OR2_X2 c7201(
.A1(net7559),
.A2(net7582),
.ZN(net7587)
);

INV_X16 c7202(
.A(net9825),
.ZN(net7588)
);

NOR2_X4 c7203(
.A1(net7583),
.A2(net7582),
.ZN(net7589)
);

OR3_X1 c7204(
.A1(net7578),
.A2(net6597),
.A3(net10493),
.ZN(net7590)
);

MUX2_X1 c7205(
.A(net5616),
.B(net7589),
.S(net7490),
.Z(net7591)
);

AOI222_X2 c7206(
.A1(net7467),
.A2(net6629),
.B1(net7585),
.B2(net7566),
.C1(net7471),
.C2(net7581),
.ZN(net7592)
);

OAI21_X4 c7207(
.A(net6533),
.B1(net7545),
.B2(net10662),
.ZN(net7593)
);

INV_X32 c7208(
.A(net10942),
.ZN(net7594)
);

MUX2_X2 c7209(
.A(net7549),
.B(net7490),
.S(net7553),
.Z(net7595)
);

OAI22_X4 c7210(
.A1(net7592),
.A2(net7527),
.B1(net7585),
.B2(net10941),
.ZN(net7596)
);

SDFFRS_X1 c7211(
.D(net2759),
.RN(net7542),
.SE(net7585),
.SI(net5482),
.SN(net10925),
.CK(clk),
.Q(net7598),
.QN(net7597)
);

NOR2_X2 c7212(
.A1(net5503),
.A2(net4656),
.ZN(net7599)
);

NAND3_X4 c7213(
.A1(net5574),
.A2(net7563),
.A3(net7444),
.ZN(net7600)
);

XOR2_X2 c7214(
.A(net7593),
.B(net7590),
.Z(net7601)
);

OR3_X4 c7215(
.A1(net7599),
.A2(net7574),
.A3(net10565),
.ZN(net7602)
);

AND3_X2 c7216(
.A1(net5635),
.A2(net7563),
.A3(net7551),
.ZN(net7603)
);

XNOR2_X1 c7217(
.A(net7525),
.B(net7587),
.ZN(net7604)
);

OR2_X4 c7218(
.A1(net7603),
.A2(net10836),
.ZN(net7605)
);

OAI222_X1 c7219(
.A1(net7568),
.A2(net6564),
.B1(net7542),
.B2(net6612),
.C1(net7605),
.C2(net7585),
.ZN(net7606)
);

NOR3_X1 c7220(
.A1(net7537),
.A2(net7562),
.A3(net10879),
.ZN(net7607)
);

OR3_X2 c7221(
.A1(net5731),
.A2(net7598),
.A3(net7550),
.ZN(out19)
);

DFFRS_X1 c7222(
.D(net4782),
.RN(net6721),
.SN(net7546),
.CK(clk),
.Q(net7609),
.QN(net7608)
);

OR2_X1 c7223(
.A1(net6608),
.A2(net7546),
.ZN(net7610)
);

OAI21_X2 c7224(
.A(net3823),
.B1(net5551),
.B2(net5687),
.ZN(net7611)
);

OAI21_X1 c7225(
.A(net7457),
.B1(net6661),
.B2(net5658),
.ZN(net7612)
);

AOI21_X2 c7226(
.A(net6700),
.B1(net7588),
.B2(net6690),
.ZN(net7613)
);

AOI21_X1 c7227(
.A(net1833),
.B1(net7530),
.B2(net5720),
.ZN(net7614)
);

AOI21_X4 c7228(
.A(net4640),
.B1(net7612),
.B2(net6650),
.ZN(net7615)
);

DFFRS_X2 c7229(
.D(net5746),
.RN(net7553),
.SN(net7181),
.CK(clk),
.Q(net7617),
.QN(net7616)
);

INV_X4 c7230(
.A(net9600),
.ZN(net7618)
);

AND3_X1 c7231(
.A1(net7529),
.A2(net7445),
.A3(net7550),
.ZN(net7619)
);

NAND3_X1 c7232(
.A1(net6564),
.A2(net5667),
.A3(net3448),
.ZN(net7620)
);

NOR3_X4 c7233(
.A1(net4755),
.A2(net7609),
.A3(net6661),
.ZN(net7621)
);

SDFF_X1 c7234(
.D(net6680),
.SE(net6561),
.SI(net6721),
.CK(clk),
.Q(net7623),
.QN(net7622)
);

NOR3_X2 c7235(
.A1(net6698),
.A2(net6653),
.A3(net7597),
.ZN(net7624)
);

AND3_X4 c7236(
.A1(net6661),
.A2(net7545),
.A3(net10564),
.ZN(out8)
);

NAND3_X2 c7237(
.A1(net7621),
.A2(net7597),
.A3(net6661),
.ZN(net7625)
);

OR3_X1 c7238(
.A1(net4768),
.A2(net6680),
.A3(net5644),
.ZN(net7626)
);

MUX2_X1 c7239(
.A(net3797),
.B(net7622),
.S(net4528),
.Z(net7627)
);

OAI21_X4 c7240(
.A(net6612),
.B1(net6661),
.B2(net7581),
.ZN(out9)
);

MUX2_X2 c7241(
.A(net7530),
.B(net6561),
.S(net6683),
.Z(net7628)
);

NAND3_X4 c7242(
.A1(net7344),
.A2(net5482),
.A3(net7608),
.ZN(net7629)
);

OR3_X4 c7243(
.A1(net7550),
.A2(net7529),
.A3(out9),
.ZN(net7630)
);

AND3_X2 c7244(
.A1(net7627),
.A2(net5667),
.A3(net7494),
.ZN(net7631)
);

NOR3_X1 c7245(
.A1(net5682),
.A2(net7457),
.A3(net6652),
.ZN(net7632)
);

OR3_X2 c7246(
.A1(net6670),
.A2(net2674),
.A3(net7628),
.ZN(net7633)
);

OAI21_X2 c7247(
.A(net7623),
.B1(net6651),
.B2(net5658),
.ZN(net7634)
);

XNOR2_X2 c7248(
.A(net6664),
.B(net6684),
.ZN(net7635)
);

OAI21_X1 c7249(
.A(net7610),
.B1(net6680),
.B2(net7632),
.ZN(net7636)
);

AOI21_X2 c7250(
.A(net6405),
.B1(net7458),
.B2(net6608),
.ZN(net7637)
);

SDFFRS_X2 c7251(
.D(net7536),
.RN(net7588),
.SE(net6698),
.SI(net6648),
.SN(net6706),
.CK(clk),
.Q(net7639),
.QN(net7638)
);

SDFF_X2 c7252(
.D(net5412),
.SE(net7445),
.SI(net7545),
.CK(clk),
.Q(net7641),
.QN(net7640)
);

AOI21_X1 c7253(
.A(net3641),
.B1(net7637),
.B2(net3786),
.ZN(net7642)
);

AOI21_X4 c7254(
.A(net6649),
.B1(net4789),
.B2(net4781),
.ZN(net7643)
);

AND3_X1 c7255(
.A1(net5658),
.A2(net5723),
.A3(net7608),
.ZN(net7644)
);

NAND3_X1 c7256(
.A1(net6725),
.A2(net7640),
.A3(net10894),
.ZN(net7645)
);

NOR3_X4 c7257(
.A1(net5630),
.A2(net7638),
.A3(net10844),
.ZN(net7646)
);

OAI221_X4 c7258(
.A(net7645),
.B1(net6525),
.B2(net6700),
.C1(net7494),
.C2(net6648),
.ZN(net7647)
);

NOR3_X2 c7259(
.A1(net5672),
.A2(net4728),
.A3(net7536),
.ZN(net7648)
);

AND3_X4 c7260(
.A1(net7643),
.A2(net7546),
.A3(net6564),
.ZN(net7649)
);

NAND3_X2 c7261(
.A1(net7618),
.A2(net7628),
.A3(net3776),
.ZN(net7650)
);

OR3_X1 c7262(
.A1(net7617),
.A2(net6672),
.A3(net7640),
.ZN(net7651)
);

DFFRS_X1 c7263(
.D(net7646),
.RN(net7633),
.SN(net1833),
.CK(clk),
.Q(net7653),
.QN(net7652)
);

SDFFRS_X1 c7264(
.D(net7615),
.RN(net7344),
.SE(net1579),
.SI(out9),
.SN(net5687),
.CK(clk),
.Q(net7655),
.QN(net7654)
);

MUX2_X1 c7265(
.A(net4740),
.B(net7639),
.S(net7594),
.Z(net7656)
);

OAI21_X4 c7266(
.A(net7653),
.B1(net7632),
.B2(net10764),
.ZN(net7657)
);

MUX2_X2 c7267(
.A(net7503),
.B(net7649),
.S(net7628),
.Z(net7658)
);

NAND3_X4 c7268(
.A1(net6725),
.A2(net7653),
.A3(net6672),
.ZN(net7659)
);

OR3_X4 c7269(
.A1(net2808),
.A2(net7635),
.A3(out1),
.ZN(net7660)
);

AND3_X2 c7270(
.A1(net7641),
.A2(net7658),
.A3(net7638),
.ZN(net7661)
);

NOR3_X1 c7271(
.A1(net5644),
.A2(net7656),
.A3(net4755),
.ZN(net7662)
);

INV_X1 c7272(
.A(net9599),
.ZN(net7663)
);

DFFRS_X2 c7273(
.D(net6452),
.RN(net7653),
.SN(net7641),
.CK(clk),
.Q(net7665),
.QN(net7664)
);

AND2_X4 c7274(
.A1(net7594),
.A2(net7664),
.ZN(net7666)
);

OR3_X2 c7275(
.A1(net3777),
.A2(net7614),
.A3(net7653),
.ZN(net7667)
);

OAI21_X2 c7276(
.A(net6653),
.B1(net7619),
.B2(net4739),
.ZN(net7668)
);

OAI21_X1 c7277(
.A(net7636),
.B1(net7665),
.B2(net4528),
.ZN(net7669)
);

AOI21_X2 c7278(
.A(net6566),
.B1(net5682),
.B2(net6670),
.ZN(net7670)
);

AOI21_X1 c7279(
.A(net7626),
.B1(net3786),
.B2(net6707),
.ZN(net7671)
);

AOI21_X4 c7280(
.A(net6566),
.B1(net10887),
.B2(net10892),
.ZN(net7672)
);

AND3_X1 c7281(
.A1(net7672),
.A2(net5762),
.A3(net5745),
.ZN(net7673)
);

SDFF_X1 c7282(
.D(net6649),
.SE(net2851),
.SI(net10919),
.CK(clk),
.Q(net7675),
.QN(net7674)
);

NAND3_X1 c7283(
.A1(net4789),
.A2(net6707),
.A3(out9),
.ZN(net7676)
);

SDFF_X2 c7284(
.D(net7642),
.SE(net7655),
.SI(net7674),
.CK(clk),
.Q(net7678),
.QN(net7677)
);

NOR3_X4 c7285(
.A1(net5687),
.A2(net6650),
.A3(net10550),
.ZN(net7679)
);

AND2_X1 c7286(
.A1(net7662),
.A2(net7673),
.ZN(net7680)
);

NOR3_X2 c7287(
.A1(net7678),
.A2(net7666),
.A3(net10941),
.ZN(net7681)
);

AND3_X4 c7288(
.A1(net7630),
.A2(net7675),
.A3(net10765),
.ZN(net7682)
);

NAND3_X2 c7289(
.A1(net7680),
.A2(net7682),
.A3(net7677),
.ZN(net7683)
);

AOI22_X2 c7290(
.A1(net7620),
.A2(net7659),
.B1(net7682),
.B2(net7640),
.ZN(net7684)
);

OAI221_X2 c7291(
.A(net7670),
.B1(net7677),
.B2(net7682),
.C1(out9),
.C2(net10381),
.ZN(net7685)
);

AOI221_X4 c7292(
.A(net5687),
.B1(net7641),
.B2(net7682),
.C1(net7545),
.C2(net10381),
.ZN(net7686)
);

OR3_X1 c7293(
.A1(net7681),
.A2(net6700),
.A3(net10861),
.ZN(net7687)
);

MUX2_X1 c7294(
.A(net7675),
.B(net7657),
.S(net7652),
.Z(net7688)
);

OAI21_X4 c7295(
.A(net7628),
.B1(net6116),
.B2(net10855),
.ZN(net7689)
);

MUX2_X2 c7296(
.A(net6649),
.B(net10734),
.S(net10987),
.Z(net7690)
);

NAND3_X4 c7297(
.A1(net7663),
.A2(net7616),
.A3(net10968),
.ZN(net7691)
);

OR3_X4 c7298(
.A1(net7650),
.A2(net7652),
.A3(net10953),
.ZN(net7692)
);

DFFRS_X1 c7299(
.D(net7688),
.RN(net7674),
.SN(net11193),
.CK(clk),
.Q(net7694),
.QN(net7693)
);

SDFFS_X1 c7300(
.D(net4763),
.SE(net7668),
.SI(net7645),
.SN(net7652),
.CK(clk),
.Q(net7696),
.QN(net7695)
);

OAI222_X4 c7301(
.A1(net7609),
.A2(net7695),
.B1(net6697),
.B2(net6612),
.C1(net6721),
.C2(net10894),
.ZN(net7697)
);

AND3_X2 c7302(
.A1(net7676),
.A2(net5412),
.A3(net10919),
.ZN(net7698)
);

AOI221_X2 c7303(
.A(net4740),
.B1(net6649),
.B2(net7545),
.C1(net10895),
.C2(net10988),
.ZN(net7699)
);

NAND2_X1 c7304(
.A1(net6759),
.A2(net6779),
.ZN(net7700)
);

INV_X2 c7305(
.A(net4810),
.ZN(net7701)
);

INV_X8 c7306(
.A(net6768),
.ZN(net7702)
);

INV_X16 c7307(
.A(net6752),
.ZN(net7703)
);

NAND2_X2 c7308(
.A1(net7701),
.A2(net2884),
.ZN(net7704)
);

INV_X32 c7309(
.A(net6792),
.ZN(net7705)
);

NAND2_X4 c7310(
.A1(net6808),
.A2(net5810),
.ZN(net7706)
);

AND2_X2 c7311(
.A1(net7700),
.A2(net6740),
.ZN(net7707)
);

XOR2_X1 c7312(
.A(net5823),
.B(net6736),
.Z(net7708)
);

INV_X4 c7313(
.A(net7705),
.ZN(net7709)
);

INV_X1 c7314(
.A(net6761),
.ZN(net7710)
);

NOR3_X1 c7315(
.A1(net6729),
.A2(net6728),
.A3(net7708),
.ZN(net7711)
);

INV_X2 c7316(
.A(net9627),
.ZN(net7712)
);

INV_X8 c7317(
.A(net6753),
.ZN(net7713)
);

INV_X16 c7318(
.A(net6728),
.ZN(net7714)
);

INV_X32 c7319(
.A(net5829),
.ZN(net7715)
);

INV_X4 c7320(
.A(net4838),
.ZN(net7716)
);

INV_X1 c7321(
.A(net6804),
.ZN(net7717)
);

NOR2_X1 c7322(
.A1(net5843),
.A2(net6728),
.ZN(net7718)
);

OR2_X2 c7323(
.A1(net4841),
.A2(net6783),
.ZN(net7719)
);

NOR2_X4 c7324(
.A1(net7713),
.A2(net6790),
.ZN(net7720)
);

INV_X2 c7325(
.A(net9701),
.ZN(net7721)
);

DFFRS_X2 c7326(
.D(net6791),
.RN(net5781),
.SN(net1898),
.CK(clk),
.Q(net7723),
.QN(net7722)
);

NOR2_X2 c7327(
.A1(net2884),
.A2(net4798),
.ZN(net7724)
);

INV_X8 c7328(
.A(net10410),
.ZN(net7725)
);

XOR2_X2 c7329(
.A(net6779),
.B(net4838),
.Z(net7726)
);

INV_X16 c7330(
.A(net7703),
.ZN(net7727)
);

CLKGATETST_X1 c7331(
.E(net6729),
.SE(net6739),
.CK(clk),
.GCK(net7728)
);

INV_X32 c7332(
.A(net7725),
.ZN(net7729)
);

SDFF_X1 c7333(
.D(net7700),
.SE(net6746),
.SI(net7708),
.CK(clk),
.Q(net7731),
.QN(net7730)
);

XNOR2_X1 c7334(
.A(net7709),
.B(net7713),
.ZN(net7732)
);

OR2_X4 c7335(
.A1(net5765),
.A2(net7714),
.ZN(net7733)
);

INV_X4 c7336(
.A(net9719),
.ZN(net7734)
);

INV_X1 c7337(
.A(net9819),
.ZN(net7735)
);

OR2_X1 c7338(
.A1(net6804),
.A2(net7703),
.ZN(net7736)
);

INV_X2 c7339(
.A(net10410),
.ZN(net7737)
);

INV_X8 c7340(
.A(net7706),
.ZN(net7738)
);

INV_X16 c7341(
.A(net5795),
.ZN(net7739)
);

INV_X32 c7342(
.A(net7737),
.ZN(net7740)
);

OR3_X2 c7343(
.A1(net7725),
.A2(net7731),
.A3(net6759),
.ZN(net7741)
);

INV_X4 c7344(
.A(net7734),
.ZN(net7742)
);

INV_X1 c7345(
.A(net7706),
.ZN(net7743)
);

INV_X2 c7346(
.A(net9818),
.ZN(net7744)
);

XNOR2_X2 c7347(
.A(net7718),
.B(net6814),
.ZN(net7745)
);

AND2_X4 c7348(
.A1(net6731),
.A2(net6801),
.ZN(net7746)
);

INV_X8 c7349(
.A(net7721),
.ZN(net7747)
);

CLKGATETST_X2 c7350(
.E(net7733),
.SE(net6768),
.CK(clk),
.GCK(net7748)
);

CLKGATETST_X4 c7351(
.E(net7747),
.SE(net7745),
.CK(clk),
.GCK(net7749)
);

NAND4_X4 c7352(
.A1(net7749),
.A2(net7700),
.A3(net7729),
.A4(net6788),
.ZN(net7750)
);

AND2_X1 c7353(
.A1(net5784),
.A2(net7713),
.ZN(net7751)
);

OAI21_X2 c7354(
.A(net7720),
.B1(net7732),
.B2(net7749),
.ZN(net7752)
);

INV_X16 c7355(
.A(net7723),
.ZN(net7753)
);

INV_X32 c7356(
.A(net7753),
.ZN(net7754)
);

CLKGATETST_X8 c7357(
.E(net7748),
.SE(net5808),
.CK(clk),
.GCK(net7755)
);

INV_X4 c7358(
.A(net7741),
.ZN(net7756)
);

INV_X1 c7359(
.A(net9878),
.ZN(net7757)
);

INV_X2 c7360(
.A(net7714),
.ZN(net7758)
);

OAI21_X1 c7361(
.A(net7727),
.B1(net7747),
.B2(net7752),
.ZN(net7759)
);

DFFR_X1 c7362(
.D(net7743),
.RN(net6802),
.CK(clk),
.Q(net7761),
.QN(net7760)
);

INV_X8 c7363(
.A(net9626),
.ZN(net7762)
);

NAND2_X1 c7364(
.A1(net7729),
.A2(net7746),
.ZN(net7763)
);

NAND2_X2 c7365(
.A1(net7763),
.A2(net6757),
.ZN(net7764)
);

AOI21_X2 c7366(
.A(net7763),
.B1(net7746),
.B2(net7753),
.ZN(net7765)
);

OAI222_X2 c7367(
.A1(net7765),
.A2(net7759),
.B1(net7751),
.B2(net6763),
.C1(net7704),
.C2(net7708),
.ZN(net7766)
);

OAI211_X2 c7368(
.A(net5774),
.B(net5843),
.C1(net7754),
.C2(net7747),
.ZN(net7767)
);

DFFR_X2 c7369(
.D(net7738),
.RN(net7747),
.CK(clk),
.Q(net7769),
.QN(net7768)
);

AOI21_X1 c7370(
.A(net7769),
.B1(net7736),
.B2(net11213),
.ZN(net7770)
);

AOI21_X4 c7371(
.A(net7764),
.B1(net7742),
.B2(net7722),
.ZN(net7771)
);

DFFS_X1 c7372(
.D(net7745),
.SN(net7704),
.CK(clk),
.Q(net7773),
.QN(net7772)
);

SDFF_X2 c7373(
.D(net7771),
.SE(net7764),
.SI(net11212),
.CK(clk),
.Q(net7775),
.QN(net7774)
);

SDFFRS_X2 c7374(
.D(net7750),
.RN(net7736),
.SE(net7724),
.SI(net7730),
.SN(net7747),
.CK(clk),
.Q(net7777),
.QN(net7776)
);

AND3_X1 c7375(
.A1(net7767),
.A2(net7769),
.A3(net7747),
.ZN(net7778)
);

DFFRS_X1 c7376(
.D(net7762),
.RN(net6815),
.SN(net7778),
.CK(clk),
.Q(net7780),
.QN(net7779)
);

DFFS_X2 c7377(
.D(net7773),
.SN(net7778),
.CK(clk),
.Q(net7782),
.QN(net7781)
);

NAND2_X4 c7378(
.A1(net7748),
.A2(net7779),
.ZN(net7783)
);

CLKGATETST_X1 c7379(
.E(net7751),
.SE(net7755),
.CK(clk),
.GCK(net7784)
);

NAND3_X1 c7380(
.A1(net7737),
.A2(net7780),
.A3(net7762),
.ZN(net7785)
);

AOI222_X1 c7381(
.A1(net4865),
.A2(net7771),
.B1(net7783),
.B2(net7730),
.C1(net7747),
.C2(net937),
.ZN(net7786)
);

NOR3_X4 c7382(
.A1(net7780),
.A2(net7738),
.A3(net11214),
.ZN(net7787)
);

DFFRS_X2 c7383(
.D(net7777),
.RN(net7715),
.SN(net10568),
.CK(clk),
.Q(net7789),
.QN(net7788)
);

NOR3_X2 c7384(
.A1(net7784),
.A2(net7760),
.A3(net11215),
.ZN(net7790)
);

AND3_X4 c7385(
.A1(net7735),
.A2(net7790),
.A3(net7774),
.ZN(net7791)
);

NAND3_X2 c7386(
.A1(net7782),
.A2(net7776),
.A3(net7784),
.ZN(net7792)
);

INV_X16 c7387(
.A(net4919),
.ZN(net7793)
);

INV_X32 c7388(
.A(net6874),
.ZN(net7794)
);

INV_X4 c7389(
.A(net6817),
.ZN(net7795)
);

AND2_X2 c7390(
.A1(net3984),
.A2(net6896),
.ZN(net7796)
);

INV_X1 c7391(
.A(net9710),
.ZN(net7797)
);

INV_X2 c7392(
.A(net6746),
.ZN(net7798)
);

XOR2_X1 c7393(
.A(net6781),
.B(net7791),
.Z(net7799)
);

OR3_X1 c7394(
.A1(net7781),
.A2(net7736),
.A3(net6879),
.ZN(net7800)
);

INV_X8 c7395(
.A(net6752),
.ZN(net7801)
);

INV_X16 c7396(
.A(net9549),
.ZN(net7802)
);

INV_X32 c7397(
.A(net5861),
.ZN(net7803)
);

SDFF_X1 c7398(
.D(net7801),
.SE(net7710),
.SI(net10807),
.CK(clk),
.Q(net7805),
.QN(net7804)
);

INV_X4 c7399(
.A(net9549),
.ZN(net7806)
);

NOR2_X1 c7400(
.A1(net7773),
.A2(net5836),
.ZN(net7807)
);

INV_X1 c7401(
.A(net5941),
.ZN(net7808)
);

OR2_X2 c7402(
.A1(net7735),
.A2(net5940),
.ZN(net7809)
);

INV_X2 c7403(
.A(net937),
.ZN(net7810)
);

INV_X8 c7404(
.A(net7795),
.ZN(net7811)
);

NOR2_X4 c7405(
.A1(net7805),
.A2(net7810),
.ZN(net7812)
);

NOR2_X2 c7406(
.A1(net5933),
.A2(net6746),
.ZN(net7813)
);

INV_X16 c7407(
.A(net9767),
.ZN(net7814)
);

INV_X32 c7408(
.A(net3854),
.ZN(net7815)
);

INV_X4 c7409(
.A(net7815),
.ZN(net7816)
);

MUX2_X1 c7410(
.A(net4957),
.B(net5941),
.S(net7804),
.Z(net7817)
);

INV_X1 c7411(
.A(net10308),
.ZN(net7818)
);

INV_X2 c7412(
.A(net6840),
.ZN(net7819)
);

XOR2_X2 c7413(
.A(net7816),
.B(net5877),
.Z(net7820)
);

XNOR2_X1 c7414(
.A(net6740),
.B(net6876),
.ZN(net7821)
);

INV_X8 c7415(
.A(net10009),
.ZN(net7822)
);

INV_X16 c7416(
.A(net9912),
.ZN(net7823)
);

OAI21_X4 c7417(
.A(net7744),
.B1(net7817),
.B2(net5767),
.ZN(net7824)
);

MUX2_X2 c7418(
.A(net7808),
.B(net7810),
.S(net6736),
.Z(net7825)
);

OR2_X4 c7419(
.A1(net7798),
.A2(net7772),
.ZN(net7826)
);

INV_X32 c7420(
.A(net10334),
.ZN(net7827)
);

INV_X4 c7421(
.A(net7802),
.ZN(net7828)
);

INV_X1 c7422(
.A(net7819),
.ZN(net7829)
);

OR2_X1 c7423(
.A1(net7828),
.A2(net7796),
.ZN(net7830)
);

INV_X2 c7424(
.A(net7702),
.ZN(net7831)
);

XNOR2_X2 c7425(
.A(net7813),
.B(net5933),
.ZN(net7832)
);

NAND3_X4 c7426(
.A1(net7800),
.A2(net7702),
.A3(net7744),
.ZN(net7833)
);

INV_X8 c7427(
.A(net6736),
.ZN(net7834)
);

INV_X16 c7428(
.A(net6817),
.ZN(net7835)
);

INV_X32 c7429(
.A(net7821),
.ZN(net7836)
);

OR3_X4 c7430(
.A1(net4889),
.A2(net7793),
.A3(net7816),
.ZN(net7837)
);

INV_X4 c7431(
.A(net7809),
.ZN(net7838)
);

AND2_X4 c7432(
.A1(net7806),
.A2(net6833),
.ZN(net7839)
);

AND2_X1 c7433(
.A1(net7831),
.A2(net7837),
.ZN(net7840)
);

INV_X1 c7434(
.A(net7836),
.ZN(net7841)
);

NAND2_X1 c7435(
.A1(net7837),
.A2(net7785),
.ZN(net7842)
);

NAND2_X2 c7436(
.A1(net7797),
.A2(net6840),
.ZN(net7843)
);

AND3_X2 c7437(
.A1(net7791),
.A2(net7836),
.A3(net6896),
.ZN(net7844)
);

INV_X2 c7438(
.A(net7785),
.ZN(net7845)
);

NAND2_X4 c7439(
.A1(net7842),
.A2(net7833),
.ZN(net7846)
);

AND2_X2 c7440(
.A1(net7812),
.A2(net7841),
.ZN(net7847)
);

XOR2_X1 c7441(
.A(net6833),
.B(net7837),
.Z(net7848)
);

INV_X8 c7442(
.A(net7841),
.ZN(net7849)
);

NOR2_X1 c7443(
.A1(net7839),
.A2(net7833),
.ZN(net7850)
);

OR2_X2 c7444(
.A1(net5891),
.A2(net5869),
.ZN(net7851)
);

CLKGATETST_X2 c7445(
.E(net7825),
.SE(net7720),
.CK(clk),
.GCK(net7852)
);

NOR2_X4 c7446(
.A1(net7836),
.A2(net7851),
.ZN(net7853)
);

NOR2_X2 c7447(
.A1(net7732),
.A2(net7849),
.ZN(net7854)
);

INV_X16 c7448(
.A(net7823),
.ZN(net7855)
);

XOR2_X2 c7449(
.A(net7850),
.B(net7844),
.Z(net7856)
);

INV_X32 c7450(
.A(net7838),
.ZN(net7857)
);

XNOR2_X1 c7451(
.A(net7856),
.B(net7803),
.ZN(net7858)
);

OR2_X4 c7452(
.A1(net7845),
.A2(net7858),
.ZN(net7859)
);

NOR3_X1 c7453(
.A1(net7794),
.A2(net7857),
.A3(net6899),
.ZN(net7860)
);

INV_X4 c7454(
.A(net10148),
.ZN(net7861)
);

SDFFS_X2 c7455(
.D(net7844),
.SE(net7852),
.SI(net7849),
.SN(net7708),
.CK(clk),
.Q(net7863),
.QN(net7862)
);

OR2_X1 c7456(
.A1(net7858),
.A2(net7849),
.ZN(net7864)
);

OR4_X2 c7457(
.A1(net7852),
.A2(net7757),
.A3(net6837),
.A4(net7810),
.ZN(net7865)
);

XNOR2_X2 c7458(
.A(net7705),
.B(net7844),
.ZN(net7866)
);

SDFF_X2 c7459(
.D(net7861),
.SE(net7864),
.SI(net7837),
.CK(clk),
.Q(net7868),
.QN(net7867)
);

OR3_X2 c7460(
.A1(net7848),
.A2(net7858),
.A3(net7851),
.ZN(net7869)
);

OAI21_X2 c7461(
.A(net7803),
.B1(net7850),
.B2(net7851),
.ZN(net7870)
);

AND2_X4 c7462(
.A1(net7853),
.A2(net7717),
.ZN(net7871)
);

AND2_X1 c7463(
.A1(net7830),
.A2(net7867),
.ZN(net7872)
);

OAI21_X1 c7464(
.A(net7817),
.B1(net7857),
.B2(net7871),
.ZN(net7873)
);

AOI21_X2 c7465(
.A(net7860),
.B1(net7852),
.B2(net7833),
.ZN(net7874)
);

NAND2_X1 c7466(
.A1(net7863),
.A2(net10744),
.ZN(net7875)
);

AOI21_X1 c7467(
.A(net141),
.B1(net7875),
.B2(net7871),
.ZN(net7876)
);

SDFFRS_X1 c7468(
.D(net7871),
.RN(net7850),
.SE(net7875),
.SI(net7876),
.SN(net6786),
.CK(clk),
.Q(net7878),
.QN(net7877)
);

AOI221_X1 c7469(
.A(net7811),
.B1(net7875),
.B2(net7876),
.C1(net7877),
.C2(net6896),
.ZN(net7879)
);

INV_X1 c7470(
.A(net9741),
.ZN(net7880)
);

INV_X2 c7471(
.A(net11064),
.ZN(net7881)
);

INV_X8 c7472(
.A(net10204),
.ZN(net7882)
);

DFFRS_X1 c7473(
.D(net7834),
.RN(net7835),
.SN(net5940),
.CK(clk),
.Q(net7884),
.QN(net7883)
);

NAND2_X2 c7474(
.A1(net6976),
.A2(net7884),
.ZN(net7885)
);

INV_X16 c7475(
.A(net6919),
.ZN(net7886)
);

INV_X32 c7476(
.A(net7769),
.ZN(net7887)
);

NAND2_X4 c7477(
.A1(net7789),
.A2(net7887),
.ZN(net7888)
);

INV_X4 c7478(
.A(net5965),
.ZN(net7889)
);

INV_X1 c7479(
.A(net7832),
.ZN(net7890)
);

INV_X2 c7480(
.A(net10869),
.ZN(net7891)
);

AND2_X2 c7481(
.A1(net6814),
.A2(net5026),
.ZN(net7892)
);

XOR2_X1 c7482(
.A(net6928),
.B(net7801),
.Z(net7893)
);

INV_X8 c7483(
.A(net9664),
.ZN(net7894)
);

INV_X16 c7484(
.A(net7790),
.ZN(net7895)
);

INV_X32 c7485(
.A(net10146),
.ZN(net7896)
);

NOR2_X1 c7486(
.A1(net7896),
.A2(net6969),
.ZN(net7897)
);

OR2_X2 c7487(
.A1(net6019),
.A2(net7887),
.ZN(net7898)
);

NOR2_X4 c7488(
.A1(net6784),
.A2(net7788),
.ZN(net7899)
);

AOI21_X4 c7489(
.A(net7829),
.B1(net5836),
.B2(net7883),
.ZN(net7900)
);

NOR2_X2 c7490(
.A1(net5985),
.A2(net7768),
.ZN(net7901)
);

XOR2_X2 c7491(
.A(net6969),
.B(net4934),
.Z(net7902)
);

XNOR2_X1 c7492(
.A(net7827),
.B(net5935),
.ZN(net7903)
);

INV_X4 c7493(
.A(net7889),
.ZN(net7904)
);

OR2_X4 c7494(
.A1(net7870),
.A2(net7888),
.ZN(net7905)
);

AND3_X1 c7495(
.A1(net7901),
.A2(net7892),
.A3(net6927),
.ZN(net7906)
);

INV_X1 c7496(
.A(net9877),
.ZN(net7907)
);

OR2_X1 c7497(
.A1(net3920),
.A2(net7903),
.ZN(net7908)
);

INV_X2 c7498(
.A(net9718),
.ZN(net7909)
);

INV_X8 c7499(
.A(net7872),
.ZN(net7910)
);

INV_X16 c7500(
.A(net10217),
.ZN(net7911)
);

XNOR2_X2 c7501(
.A(net7904),
.B(net7893),
.ZN(net7912)
);

AND2_X4 c7502(
.A1(net7857),
.A2(net7884),
.ZN(net7913)
);

INV_X32 c7503(
.A(net10060),
.ZN(net7914)
);

INV_X4 c7504(
.A(net10423),
.ZN(net7915)
);

AND2_X1 c7505(
.A1(net7880),
.A2(net6852),
.ZN(net7916)
);

NAND2_X1 c7506(
.A1(net7900),
.A2(net6966),
.ZN(net7917)
);

NAND3_X1 c7507(
.A1(net6844),
.A2(net7827),
.A3(net6966),
.ZN(net7918)
);

NOR3_X4 c7508(
.A1(net5033),
.A2(net7908),
.A3(net10491),
.ZN(net7919)
);

NAND2_X2 c7509(
.A1(net6900),
.A2(net7880),
.ZN(net7920)
);

INV_X1 c7510(
.A(net10423),
.ZN(net7921)
);

NOR3_X2 c7511(
.A1(net7898),
.A2(net7920),
.A3(net7876),
.ZN(net7922)
);

INV_X2 c7512(
.A(net7895),
.ZN(net7923)
);

AND3_X4 c7513(
.A1(net7907),
.A2(net7908),
.A3(net11053),
.ZN(net7924)
);

INV_X8 c7514(
.A(net10187),
.ZN(net7925)
);

INV_X16 c7515(
.A(net6962),
.ZN(net7926)
);

INV_X32 c7516(
.A(net11019),
.ZN(net7927)
);

NAND2_X4 c7517(
.A1(net6868),
.A2(net6844),
.ZN(net7928)
);

AND2_X2 c7518(
.A1(net6802),
.A2(net7790),
.ZN(net7929)
);

INV_X4 c7519(
.A(net7909),
.ZN(net7930)
);

NAND3_X2 c7520(
.A1(net6913),
.A2(net7922),
.A3(net7731),
.ZN(net7931)
);

XOR2_X1 c7521(
.A(net7810),
.B(net11136),
.Z(net7932)
);

INV_X1 c7522(
.A(net9664),
.ZN(net7933)
);

NOR2_X1 c7523(
.A1(net5977),
.A2(net7758),
.ZN(net7934)
);

OR3_X1 c7524(
.A1(net7770),
.A2(net6951),
.A3(net10954),
.ZN(net7935)
);

OR2_X2 c7525(
.A1(net6762),
.A2(net7925),
.ZN(net7936)
);

NOR2_X4 c7526(
.A1(net7742),
.A2(net7927),
.ZN(net7937)
);

INV_X2 c7527(
.A(net7913),
.ZN(net7938)
);

MUX2_X1 c7528(
.A(net7927),
.B(net7917),
.S(net10389),
.Z(net7939)
);

NOR2_X2 c7529(
.A1(net7897),
.A2(net7927),
.ZN(net7940)
);

AOI211_X1 c7530(
.A(net7938),
.B(net7936),
.C1(net7874),
.C2(net7768),
.ZN(net7941)
);

OAI21_X4 c7531(
.A(net7892),
.B1(net7835),
.B2(net6919),
.ZN(net7942)
);

MUX2_X2 c7532(
.A(net7916),
.B(net7892),
.S(net6908),
.Z(net7943)
);

XOR2_X2 c7533(
.A(net7851),
.B(net7887),
.Z(net7944)
);

XNOR2_X1 c7534(
.A(net7930),
.B(net11053),
.ZN(net7945)
);

INV_X8 c7535(
.A(net7939),
.ZN(net7946)
);

OR2_X4 c7536(
.A1(net7930),
.A2(net10434),
.ZN(net7947)
);

OR2_X1 c7537(
.A1(net7933),
.A2(net10954),
.ZN(net7948)
);

DFFRS_X2 c7538(
.D(net7919),
.RN(net7920),
.SN(net7922),
.CK(clk),
.Q(net7950),
.QN(net7949)
);

XNOR2_X2 c7539(
.A(net7907),
.B(net7886),
.ZN(net7951)
);

NAND3_X4 c7540(
.A1(net5972),
.A2(net7951),
.A3(net7941),
.ZN(net7952)
);

OAI221_X1 c7541(
.A(net7887),
.B1(net7929),
.B2(net4934),
.C1(net7888),
.C2(net7768),
.ZN(net7953)
);

INV_X16 c7542(
.A(net10203),
.ZN(net7954)
);

OR3_X4 c7543(
.A1(net7900),
.A2(net7886),
.A3(net11063),
.ZN(net7955)
);

AND3_X2 c7544(
.A1(net7947),
.A2(net7944),
.A3(net7937),
.ZN(net7956)
);

SDFFR_X1 c7545(
.D(net7892),
.RN(net7949),
.SE(net6955),
.SI(net10581),
.CK(clk),
.Q(net7958),
.QN(net7957)
);

NOR3_X1 c7546(
.A1(net7953),
.A2(net7950),
.A3(net5045),
.ZN(net7959)
);

INV_X32 c7547(
.A(net11064),
.ZN(net7960)
);

AND2_X4 c7548(
.A1(net7955),
.A2(net7960),
.ZN(net7961)
);

NAND4_X2 c7549(
.A1(net7899),
.A2(net7960),
.A3(net7961),
.A4(net5025),
.ZN(net7962)
);

OR3_X2 c7550(
.A1(net7757),
.A2(net7769),
.A3(net10921),
.ZN(net7963)
);

OAI221_X4 c7551(
.A(net7881),
.B1(net7962),
.B2(net7950),
.C1(net7963),
.C2(net7730),
.ZN(net7964)
);

OAI221_X2 c7552(
.A(net7954),
.B1(net7940),
.B2(net7961),
.C1(net7964),
.C2(net7888),
.ZN(net7965)
);

AND2_X1 c7553(
.A1(net7874),
.A2(net7072),
.ZN(net7966)
);

NAND2_X1 c7554(
.A1(net6943),
.A2(net6933),
.ZN(net7967)
);

NAND2_X2 c7555(
.A1(net7833),
.A2(net7894),
.ZN(net7968)
);

NAND2_X4 c7556(
.A1(net7968),
.A2(net7925),
.ZN(net7969)
);

AND2_X2 c7557(
.A1(net7770),
.A2(net6943),
.ZN(net7970)
);

XOR2_X1 c7558(
.A(net6757),
.B(net7814),
.Z(net7971)
);

NOR2_X1 c7559(
.A1(net3153),
.A2(net6027),
.ZN(net7972)
);

OR2_X2 c7560(
.A1(net7969),
.A2(net7886),
.ZN(net7973)
);

NOR2_X4 c7561(
.A1(net7967),
.A2(net7970),
.ZN(net7974)
);

NOR2_X2 c7562(
.A1(net4945),
.A2(net7062),
.ZN(net7975)
);

XOR2_X2 c7563(
.A(net7932),
.B(net6757),
.Z(net7976)
);

INV_X4 c7564(
.A(net9995),
.ZN(net7977)
);

XNOR2_X1 c7565(
.A(net7972),
.B(net7976),
.ZN(net7978)
);

OR2_X4 c7566(
.A1(net7977),
.A2(net7957),
.ZN(net7979)
);

INV_X1 c7567(
.A(net7025),
.ZN(net7980)
);

OAI21_X2 c7568(
.A(net6852),
.B1(net7966),
.B2(net7807),
.ZN(net7981)
);

OR2_X1 c7569(
.A1(net7971),
.A2(net7979),
.ZN(net7982)
);

INV_X2 c7570(
.A(net10958),
.ZN(net7983)
);

XNOR2_X2 c7571(
.A(net6883),
.B(net7927),
.ZN(net7984)
);

AND2_X4 c7572(
.A1(net7846),
.A2(net7917),
.ZN(net7985)
);

AND2_X1 c7573(
.A1(net7979),
.A2(net7967),
.ZN(net7986)
);

NAND2_X1 c7574(
.A1(net7976),
.A2(net7920),
.ZN(net7987)
);

CLKGATETST_X4 c7575(
.E(net7004),
.SE(net7025),
.CK(clk),
.GCK(net7988)
);

INV_X8 c7576(
.A(net7981),
.ZN(net7989)
);

INV_X16 c7577(
.A(net7882),
.ZN(net7990)
);

OR4_X4 c7578(
.A1(net7925),
.A2(net7066),
.A3(net7847),
.A4(net7053),
.ZN(net7991)
);

NAND2_X2 c7579(
.A1(net7973),
.A2(net7903),
.ZN(net7992)
);

NAND2_X4 c7580(
.A1(net7988),
.A2(net7990),
.ZN(net7993)
);

AND2_X2 c7581(
.A1(net6926),
.A2(net7951),
.ZN(net7994)
);

XOR2_X1 c7582(
.A(net7974),
.B(net7903),
.Z(net7995)
);

NOR2_X1 c7583(
.A1(net7958),
.A2(net7979),
.ZN(net7996)
);

OR2_X2 c7584(
.A1(net7980),
.A2(net7956),
.ZN(net7997)
);

NOR2_X4 c7585(
.A1(net7970),
.A2(net7000),
.ZN(net7998)
);

NOR2_X2 c7586(
.A1(net7989),
.A2(net7000),
.ZN(net7999)
);

INV_X32 c7587(
.A(net7999),
.ZN(net8000)
);

OAI21_X1 c7588(
.A(net6879),
.B1(net7874),
.B2(net7996),
.ZN(net8001)
);

XOR2_X2 c7589(
.A(net8001),
.B(net6926),
.Z(net8002)
);

AOI21_X2 c7590(
.A(net4934),
.B1(net7988),
.B2(net7968),
.ZN(net8003)
);

INV_X4 c7591(
.A(net9938),
.ZN(net8004)
);

XNOR2_X1 c7592(
.A(net7923),
.B(net7990),
.ZN(net8005)
);

INV_X1 c7593(
.A(net10182),
.ZN(net8006)
);

OR2_X4 c7594(
.A1(net7993),
.A2(net7997),
.ZN(net8007)
);

SDFF_X1 c7595(
.D(net7825),
.SE(net6955),
.SI(net7968),
.CK(clk),
.Q(net8009),
.QN(net8008)
);

OR2_X1 c7596(
.A1(net6955),
.A2(net7941),
.ZN(net8010)
);

SDFF_X2 c7597(
.D(net8007),
.SE(net6879),
.SI(net7918),
.CK(clk),
.Q(net8012),
.QN(net8011)
);

OAI22_X2 c7598(
.A1(net7067),
.A2(net8006),
.B1(net7967),
.B2(net8003),
.ZN(net8013)
);

XNOR2_X2 c7599(
.A(net7940),
.B(net7025),
.ZN(net8014)
);

AND2_X4 c7600(
.A1(net7903),
.A2(net6091),
.ZN(net8015)
);

CLKGATETST_X8 c7601(
.E(net7034),
.SE(net10390),
.CK(clk),
.GCK(net8016)
);

AND2_X1 c7602(
.A1(net7975),
.A2(net8014),
.ZN(net8017)
);

NAND2_X1 c7603(
.A1(net7847),
.A2(net7917),
.ZN(net8018)
);

INV_X2 c7604(
.A(net9776),
.ZN(net8019)
);

OAI211_X4 c7605(
.A(net8019),
.B(net5142),
.C1(net5934),
.C2(net8016),
.ZN(net8020)
);

NAND2_X2 c7606(
.A1(net8012),
.A2(net7997),
.ZN(net8021)
);

NAND2_X4 c7607(
.A1(net5142),
.A2(net5046),
.ZN(net8022)
);

AND2_X2 c7608(
.A1(net7994),
.A2(net8014),
.ZN(net8023)
);

XOR2_X1 c7609(
.A(net7991),
.B(net8011),
.Z(net8024)
);

INV_X8 c7610(
.A(net10075),
.ZN(net8025)
);

NOR2_X1 c7611(
.A1(net7843),
.A2(net4945),
.ZN(net8026)
);

OAI211_X1 c7612(
.A(net7978),
.B(net8024),
.C1(net5072),
.C2(net7964),
.ZN(net8027)
);

AOI21_X1 c7613(
.A(net5973),
.B1(net8008),
.B2(net11027),
.ZN(net8028)
);

OR2_X2 c7614(
.A1(net8028),
.A2(net8020),
.ZN(net8029)
);

NOR2_X4 c7615(
.A1(net7921),
.A2(net7990),
.ZN(net8030)
);

SDFFRS_X2 c7616(
.D(net7775),
.RN(net6883),
.SE(net7034),
.SI(net7968),
.SN(net7996),
.CK(clk),
.Q(net8032),
.QN(net8031)
);

INV_X16 c7617(
.A(net11072),
.ZN(net8033)
);

NOR2_X2 c7618(
.A1(net8033),
.A2(net8031),
.ZN(net8034)
);

DFFRS_X1 c7619(
.D(net8006),
.RN(net7034),
.SN(net8020),
.CK(clk),
.Q(net8036),
.QN(net8035)
);

AOI21_X4 c7620(
.A(net5836),
.B1(net7796),
.B2(net8014),
.ZN(net8037)
);

XOR2_X2 c7621(
.A(net8005),
.B(net8036),
.Z(net8038)
);

AND3_X1 c7622(
.A1(net7062),
.A2(net7979),
.A3(net8025),
.ZN(net8039)
);

NAND3_X1 c7623(
.A1(net7984),
.A2(net8037),
.A3(net8035),
.ZN(net8040)
);

AOI222_X4 c7624(
.A1(net8026),
.A2(net8036),
.B1(net5142),
.B2(net7996),
.C1(net7810),
.C2(net10914),
.ZN(net8041)
);

XNOR2_X1 c7625(
.A(net8025),
.B(net8039),
.ZN(net8042)
);

NOR4_X4 c7626(
.A1(net8009),
.A2(net8033),
.A3(net8007),
.A4(net8031),
.ZN(net8043)
);

NOR3_X4 c7627(
.A1(net8042),
.A2(net8039),
.A3(net11098),
.ZN(net8044)
);

INV_X32 c7628(
.A(net10958),
.ZN(net8045)
);

NOR3_X2 c7629(
.A1(net6951),
.A2(net7770),
.A3(net10914),
.ZN(net8046)
);

AND3_X4 c7630(
.A1(net8038),
.A2(net8020),
.A3(net10848),
.ZN(net8047)
);

NOR4_X2 c7631(
.A1(net8037),
.A2(net8034),
.A3(net6991),
.A4(net10849),
.ZN(net8048)
);

OR2_X4 c7632(
.A1(net8018),
.A2(net8047),
.ZN(net8049)
);

NAND3_X2 c7633(
.A1(net8041),
.A2(net8049),
.A3(net8037),
.ZN(net8050)
);

OAI33_X1 c7634(
.A1(net8016),
.A2(net8017),
.A3(net8014),
.B1(net8020),
.B2(net7996),
.B3(net11081),
.ZN(net8051)
);

OR3_X1 c7635(
.A1(net8049),
.A2(net7049),
.A3(net8017),
.ZN(net8052)
);

OR2_X1 c7636(
.A1(net8045),
.A2(net6799),
.ZN(net8053)
);

XNOR2_X2 c7637(
.A(net6108),
.B(net7908),
.ZN(net8054)
);

MUX2_X1 c7638(
.A(net8039),
.B(net7118),
.S(net7822),
.Z(net8055)
);

AND2_X4 c7639(
.A1(net7005),
.A2(net8020),
.ZN(net8056)
);

AOI211_X4 c7640(
.A(net6902),
.B(net5072),
.C1(net6129),
.C2(net6160),
.ZN(net8057)
);

INV_X4 c7641(
.A(net8020),
.ZN(net8058)
);

AND2_X1 c7642(
.A1(net7865),
.A2(net8057),
.ZN(net8059)
);

INV_X1 c7643(
.A(net11115),
.ZN(net8060)
);

NAND2_X1 c7644(
.A1(net7132),
.A2(net8045),
.ZN(net8061)
);

INV_X2 c7645(
.A(net9570),
.ZN(net8062)
);

OAI21_X4 c7646(
.A(net8048),
.B1(net7084),
.B2(net11001),
.ZN(net8063)
);

NAND2_X2 c7647(
.A1(net8039),
.A2(net10623),
.ZN(net8064)
);

NAND2_X4 c7648(
.A1(net7890),
.A2(net8053),
.ZN(net8065)
);

AND2_X2 c7649(
.A1(net6160),
.A2(net10653),
.ZN(net8066)
);

XOR2_X1 c7650(
.A(net8062),
.B(net6086),
.Z(net8067)
);

NOR2_X1 c7651(
.A1(net7090),
.A2(net7087),
.ZN(net8068)
);

OR2_X2 c7652(
.A1(net2244),
.A2(net7990),
.ZN(net8069)
);

INV_X8 c7653(
.A(net8068),
.ZN(net8070)
);

NOR2_X4 c7654(
.A1(net8066),
.A2(net7863),
.ZN(net8071)
);

INV_X16 c7655(
.A(net10101),
.ZN(net8072)
);

NOR2_X2 c7656(
.A1(net8060),
.A2(net7822),
.ZN(net8073)
);

MUX2_X2 c7657(
.A(net7078),
.B(net8015),
.S(net7796),
.Z(net8074)
);

INV_X32 c7658(
.A(net5072),
.ZN(net8075)
);

INV_X4 c7659(
.A(net9817),
.ZN(net8076)
);

INV_X1 c7660(
.A(net11055),
.ZN(net8077)
);

XOR2_X2 c7661(
.A(net6129),
.B(net7951),
.Z(net8078)
);

XNOR2_X1 c7662(
.A(net4261),
.B(net10566),
.ZN(net8079)
);

INV_X2 c7663(
.A(net10290),
.ZN(net8080)
);

OR2_X4 c7664(
.A1(net7164),
.A2(net10700),
.ZN(net8081)
);

OR2_X1 c7665(
.A1(net8067),
.A2(net7807),
.ZN(net8082)
);

DFFR_X1 c7666(
.D(net7948),
.RN(net7165),
.CK(clk),
.Q(net8084),
.QN(net8083)
);

XNOR2_X2 c7667(
.A(net7000),
.B(net8083),
.ZN(net8085)
);

AND2_X4 c7668(
.A1(net7997),
.A2(net7118),
.ZN(net8086)
);

NAND3_X4 c7669(
.A1(net8071),
.A2(net5166),
.A3(net7088),
.ZN(net8087)
);

AND2_X1 c7670(
.A1(net8079),
.A2(net2244),
.ZN(net8088)
);

NAND2_X1 c7671(
.A1(net7946),
.A2(net7163),
.ZN(net8089)
);

OR3_X4 c7672(
.A1(net8074),
.A2(net6086),
.A3(net8082),
.ZN(net8090)
);

NAND2_X2 c7673(
.A1(net8088),
.A2(net7141),
.ZN(net8091)
);

INV_X8 c7674(
.A(net10267),
.ZN(net8092)
);

INV_X16 c7675(
.A(net11035),
.ZN(net8093)
);

NAND2_X4 c7676(
.A1(net7137),
.A2(net8074),
.ZN(net8094)
);

AND3_X2 c7677(
.A1(net8082),
.A2(net8032),
.A3(net8034),
.ZN(net8095)
);

DFFR_X2 c7678(
.D(net8064),
.RN(net7126),
.CK(clk),
.Q(net8097),
.QN(net8096)
);

AND2_X2 c7679(
.A1(net7163),
.A2(net7147),
.ZN(out13)
);

XOR2_X1 c7680(
.A(net8085),
.B(net4840),
.Z(net8098)
);

NOR2_X1 c7681(
.A1(net5214),
.A2(net2244),
.ZN(net8099)
);

OR2_X2 c7682(
.A1(net8093),
.A2(net8099),
.ZN(net8100)
);

NOR2_X4 c7683(
.A1(net7990),
.A2(net8097),
.ZN(net8101)
);

NOR2_X2 c7684(
.A1(net8092),
.A2(net6902),
.ZN(net8102)
);

INV_X32 c7685(
.A(net9914),
.ZN(net8103)
);

DFFS_X1 c7686(
.D(net8086),
.SN(net7818),
.CK(clk),
.Q(net8105),
.QN(net8104)
);

INV_X4 c7687(
.A(net10269),
.ZN(net8106)
);

AOI221_X4 c7688(
.A(net4223),
.B1(net7930),
.B2(net8103),
.C1(net8053),
.C2(net8070),
.ZN(net8107)
);

DFFRS_X2 c7689(
.D(net7708),
.RN(net8100),
.SN(net8099),
.CK(clk),
.Q(net8109),
.QN(net8108)
);

NOR3_X1 c7690(
.A1(net8080),
.A2(net8075),
.A3(net8053),
.ZN(net8110)
);

AOI221_X2 c7691(
.A(net8103),
.B1(net7077),
.B2(net8082),
.C1(out13),
.C2(net7996),
.ZN(net8111)
);

INV_X1 c7692(
.A(net9770),
.ZN(net8112)
);

XOR2_X2 c7693(
.A(net8098),
.B(net8060),
.Z(net8113)
);

XNOR2_X1 c7694(
.A(net8089),
.B(net7087),
.ZN(net8114)
);

INV_X2 c7695(
.A(net10016),
.ZN(net8115)
);

OR2_X4 c7696(
.A1(net8109),
.A2(net8061),
.ZN(net8116)
);

OR3_X2 c7697(
.A1(net7118),
.A2(net8114),
.A3(net8108),
.ZN(net8117)
);

OR2_X1 c7698(
.A1(net8102),
.A2(net7163),
.ZN(net8118)
);

XNOR2_X2 c7699(
.A(net8118),
.B(net8109),
.ZN(net8119)
);

OAI21_X2 c7700(
.A(net7995),
.B1(net8119),
.B2(net6908),
.ZN(net8120)
);

INV_X8 c7701(
.A(net9775),
.ZN(net8121)
);

INV_X16 c7702(
.A(net9569),
.ZN(net8122)
);

OAI21_X1 c7703(
.A(net8107),
.B1(net8102),
.B2(net8116),
.ZN(net8123)
);

AOI21_X2 c7704(
.A(net8072),
.B1(net7985),
.B2(net8101),
.ZN(net8124)
);

AOI21_X1 c7705(
.A(net5154),
.B1(net8117),
.B2(net8054),
.ZN(net8125)
);

AND2_X4 c7706(
.A1(net8115),
.A2(net2244),
.ZN(net8126)
);

AOI21_X4 c7707(
.A(net8113),
.B1(net8106),
.B2(net8098),
.ZN(net8127)
);

AND2_X1 c7708(
.A1(net8122),
.A2(net10386),
.ZN(net8128)
);

AND3_X1 c7709(
.A1(net8101),
.A2(net7140),
.A3(net8127),
.ZN(net8129)
);

NAND3_X1 c7710(
.A1(net7141),
.A2(net8103),
.A3(net8127),
.ZN(net8130)
);

AOI222_X2 c7711(
.A1(net8099),
.A2(net8094),
.B1(net8130),
.B2(net8119),
.C1(net7126),
.C2(net7164),
.ZN(net8131)
);

NOR3_X4 c7712(
.A1(net7866),
.A2(net8123),
.A3(net11218),
.ZN(net8132)
);

NOR3_X2 c7713(
.A1(net8124),
.A2(net8128),
.A3(net8127),
.ZN(net8133)
);

AND3_X4 c7714(
.A1(net8130),
.A2(net8122),
.A3(net8132),
.ZN(net8134)
);

NAND3_X2 c7715(
.A1(net8112),
.A2(net7141),
.A3(net10385),
.ZN(net8135)
);

SDFF_X1 c7716(
.D(net8058),
.SE(net8103),
.SI(net8091),
.CK(clk),
.Q(net8137),
.QN(net8136)
);

OR3_X1 c7717(
.A1(net8095),
.A2(net8137),
.A3(net7995),
.ZN(net8138)
);

OAI222_X1 c7718(
.A1(net8122),
.A2(net8127),
.B1(net8102),
.B2(net8136),
.C1(net7164),
.C2(out13),
.ZN(net8139)
);

INV_X32 c7719(
.A(net5167),
.ZN(net8140)
);

NAND2_X1 c7720(
.A1(net7945),
.A2(net7053),
.ZN(net8141)
);

NAND2_X2 c7721(
.A1(net6213),
.A2(net10586),
.ZN(net8142)
);

NAND2_X4 c7722(
.A1(net7203),
.A2(net7036),
.ZN(net8143)
);

INV_X4 c7723(
.A(net6210),
.ZN(net8144)
);

INV_X1 c7724(
.A(net9632),
.ZN(net8145)
);

AND2_X2 c7725(
.A1(net5935),
.A2(net6213),
.ZN(net8146)
);

XOR2_X1 c7726(
.A(net7926),
.B(net6177),
.Z(net8147)
);

NOR4_X1 c7727(
.A1(net7053),
.A2(net5818),
.A3(net7193),
.A4(net8111),
.ZN(net8148)
);

INV_X2 c7728(
.A(net9960),
.ZN(net8149)
);

NOR2_X1 c7729(
.A1(net7193),
.A2(net7036),
.ZN(net8150)
);

INV_X8 c7730(
.A(net8129),
.ZN(net8151)
);

DFFS_X2 c7731(
.D(net7250),
.SN(net6248),
.CK(clk),
.Q(net8153),
.QN(net8152)
);

OAI222_X4 c7732(
.A1(net8036),
.A2(net7818),
.B1(net7221),
.B2(net7810),
.C1(net7083),
.C2(net7930),
.ZN(net8154)
);

INV_X16 c7733(
.A(net7937),
.ZN(net8155)
);

OR2_X2 c7734(
.A1(net8084),
.A2(net7221),
.ZN(net8156)
);

MUX2_X1 c7735(
.A(net7241),
.B(net7164),
.S(net11046),
.Z(net8157)
);

NOR2_X4 c7736(
.A1(net8149),
.A2(net8146),
.ZN(net8158)
);

INV_X32 c7737(
.A(net9828),
.ZN(net8159)
);

INV_X4 c7738(
.A(net7194),
.ZN(net8160)
);

NOR2_X2 c7739(
.A1(net6248),
.A2(net7036),
.ZN(net8161)
);

INV_X1 c7740(
.A(net9798),
.ZN(net8162)
);

XOR2_X2 c7741(
.A(net7911),
.B(net7189),
.Z(net8163)
);

XNOR2_X1 c7742(
.A(net7917),
.B(net8003),
.ZN(net8164)
);

OR2_X4 c7743(
.A1(net6213),
.A2(net5848),
.ZN(net8165)
);

OR2_X1 c7744(
.A1(net8015),
.A2(net6086),
.ZN(net8166)
);

XNOR2_X2 c7745(
.A(net7248),
.B(net7965),
.ZN(net8167)
);

AND2_X4 c7746(
.A1(net8162),
.A2(net7053),
.ZN(net8168)
);

INV_X2 c7747(
.A(net10158),
.ZN(net8169)
);

INV_X8 c7748(
.A(net9847),
.ZN(net8170)
);

AND2_X1 c7749(
.A1(net8143),
.A2(net7965),
.ZN(net8171)
);

SDFF_X2 c7750(
.D(net8157),
.SE(net7248),
.SI(net8168),
.CK(clk),
.Q(net8173),
.QN(net8172)
);

SDFFR_X2 c7751(
.D(net8167),
.RN(net7908),
.SE(net8031),
.SI(net7083),
.CK(clk),
.Q(net8175),
.QN(net8174)
);

INV_X16 c7752(
.A(net11098),
.ZN(net8176)
);

INV_X32 c7753(
.A(net9799),
.ZN(net8177)
);

CLKGATETST_X1 c7754(
.E(net8158),
.SE(net8061),
.CK(clk),
.GCK(net8178)
);

NAND2_X1 c7755(
.A1(net1380),
.A2(net8160),
.ZN(net8179)
);

NAND2_X2 c7756(
.A1(net8166),
.A2(net8144),
.ZN(net8180)
);

INV_X4 c7757(
.A(net11059),
.ZN(net8181)
);

INV_X1 c7758(
.A(net7126),
.ZN(net8182)
);

INV_X2 c7759(
.A(net11059),
.ZN(net8183)
);

INV_X8 c7760(
.A(net8077),
.ZN(net8184)
);

NAND2_X4 c7761(
.A1(net8173),
.A2(net8182),
.ZN(net8185)
);

AND2_X2 c7762(
.A1(net5837),
.A2(net8160),
.ZN(net8186)
);

XOR2_X1 c7763(
.A(net7036),
.B(net7945),
.Z(net8187)
);

NOR2_X1 c7764(
.A1(net6899),
.A2(net8174),
.ZN(net8188)
);

OR2_X2 c7765(
.A1(net8151),
.A2(net8178),
.ZN(net8189)
);

INV_X16 c7766(
.A(net7233),
.ZN(net8190)
);

NOR2_X4 c7767(
.A1(net7084),
.A2(out13),
.ZN(net8191)
);

AOI211_X2 c7768(
.A(net7220),
.B(net8146),
.C1(net8182),
.C2(net8187),
.ZN(net8192)
);

NOR2_X2 c7769(
.A1(net7077),
.A2(net8057),
.ZN(net8193)
);

XOR2_X2 c7770(
.A(net8190),
.B(net11046),
.Z(net8194)
);

XNOR2_X1 c7771(
.A(net8185),
.B(net7164),
.ZN(net8195)
);

INV_X32 c7772(
.A(net10040),
.ZN(net8196)
);

AOI221_X1 c7773(
.A(net7239),
.B1(net8144),
.B2(net8166),
.C1(net7200),
.C2(net8182),
.ZN(net8197)
);

OR2_X4 c7774(
.A1(net8196),
.A2(net8172),
.ZN(net8198)
);

OAI21_X4 c7775(
.A(net8175),
.B1(net8034),
.B2(net8198),
.ZN(net8199)
);

MUX2_X2 c7776(
.A(net8146),
.B(net8196),
.S(net8104),
.Z(net8200)
);

AOI22_X1 c7777(
.A1(net8192),
.A2(net8187),
.B1(net8197),
.B2(net7096),
.ZN(net8201)
);

INV_X4 c7778(
.A(net9727),
.ZN(net8202)
);

INV_X1 c7779(
.A(net10932),
.ZN(net8203)
);

OR2_X1 c7780(
.A1(net8179),
.A2(net6028),
.ZN(net8204)
);

NAND3_X4 c7781(
.A1(net8183),
.A2(net8190),
.A3(net7053),
.ZN(net8205)
);

XNOR2_X2 c7782(
.A(net8057),
.B(net11219),
.ZN(net8206)
);

OR3_X4 c7783(
.A1(net7140),
.A2(net8164),
.A3(net8084),
.ZN(net8207)
);

DFFRS_X1 c7784(
.D(net8170),
.RN(net8204),
.SN(net8192),
.CK(clk),
.Q(net8209),
.QN(net8208)
);

AND2_X4 c7785(
.A1(net8194),
.A2(net8207),
.ZN(net8210)
);

INV_X2 c7786(
.A(net10052),
.ZN(net8211)
);

AND2_X1 c7787(
.A1(net8166),
.A2(net10453),
.ZN(net8212)
);

AND3_X2 c7788(
.A1(net8141),
.A2(net8202),
.A3(net8208),
.ZN(net8213)
);

INV_X8 c7789(
.A(net9631),
.ZN(net8214)
);

NAND2_X1 c7790(
.A1(net8191),
.A2(net7053),
.ZN(net8215)
);

AND4_X4 c7791(
.A1(net8212),
.A2(net8190),
.A3(net8179),
.A4(net7200),
.ZN(net8216)
);

NOR3_X1 c7792(
.A1(net8203),
.A2(net8210),
.A3(net8212),
.ZN(net8217)
);

OR3_X2 c7793(
.A1(net8188),
.A2(net8202),
.A3(net8205),
.ZN(net8218)
);

NAND2_X2 c7794(
.A1(net8218),
.A2(net10791),
.ZN(net8219)
);

NAND4_X1 c7795(
.A1(net8215),
.A2(net8206),
.A3(net8218),
.A4(out13),
.ZN(net8220)
);

OAI21_X2 c7796(
.A(net8177),
.B1(net8179),
.B2(net11096),
.ZN(net8221)
);

OAI21_X1 c7797(
.A(net8217),
.B1(net8214),
.B2(net11096),
.ZN(net8222)
);

OAI222_X2 c7798(
.A1(net8180),
.A2(net8221),
.B1(net8218),
.B2(net8197),
.C1(net7125),
.C2(net8178),
.ZN(net8223)
);

DFFRS_X2 c7799(
.D(net8159),
.RN(net8121),
.SN(net8223),
.CK(clk),
.Q(net8225),
.QN(net8224)
);

OAI221_X1 c7800(
.A(net8144),
.B1(net8217),
.B2(net8224),
.C1(net8218),
.C2(net10453),
.ZN(net8226)
);

OR4_X1 c7801(
.A1(net8211),
.A2(net8221),
.A3(net8217),
.A4(net8224),
.ZN(net8227)
);

NAND2_X4 c7802(
.A1(net7260),
.A2(net7224),
.ZN(net8228)
);

AND2_X2 c7803(
.A1(net6332),
.A2(net6987),
.ZN(net8229)
);

INV_X16 c7804(
.A(net9581),
.ZN(net8230)
);

XOR2_X1 c7805(
.A(net7224),
.B(net8187),
.Z(net8231)
);

NOR2_X1 c7806(
.A1(net548),
.A2(net8168),
.ZN(net8232)
);

AOI21_X2 c7807(
.A(net8205),
.B1(net8197),
.B2(net7275),
.ZN(net8233)
);

AOI21_X1 c7808(
.A(net8164),
.B1(net7208),
.B2(net8032),
.ZN(net8234)
);

OR2_X2 c7809(
.A1(net6373),
.A2(net10967),
.ZN(net8235)
);

INV_X32 c7810(
.A(net10349),
.ZN(net8236)
);

INV_X4 c7811(
.A(net10277),
.ZN(net8237)
);

NOR2_X4 c7812(
.A1(net8237),
.A2(net7212),
.ZN(net8238)
);

NOR2_X2 c7813(
.A1(net7241),
.A2(net7038),
.ZN(net8239)
);

AOI21_X4 c7814(
.A(net7983),
.B1(net7317),
.B2(net6373),
.ZN(net8240)
);

XOR2_X2 c7815(
.A(net8197),
.B(net7930),
.Z(net8241)
);

AND3_X1 c7816(
.A1(net8123),
.A2(net7275),
.A3(net5166),
.ZN(net8242)
);

XNOR2_X1 c7817(
.A(net7305),
.B(net7254),
.ZN(net8243)
);

NAND3_X1 c7818(
.A1(net8193),
.A2(net8238),
.A3(net7241),
.ZN(net8244)
);

OR2_X4 c7819(
.A1(net7330),
.A2(net7317),
.ZN(net8245)
);

INV_X1 c7820(
.A(net10122),
.ZN(net8246)
);

INV_X2 c7821(
.A(net11073),
.ZN(net8247)
);

OR2_X1 c7822(
.A1(net8187),
.A2(net10679),
.ZN(net8248)
);

XNOR2_X2 c7823(
.A(net7321),
.B(net5363),
.ZN(net8249)
);

NOR3_X4 c7824(
.A1(net6086),
.A2(net8238),
.A3(net7918),
.ZN(net8250)
);

CLKGATETST_X2 c7825(
.E(net8234),
.SE(net8233),
.CK(clk),
.GCK(net8251)
);

NOR3_X2 c7826(
.A1(net8059),
.A2(net7284),
.A3(net8232),
.ZN(net8252)
);

AND2_X4 c7827(
.A1(net6307),
.A2(net8242),
.ZN(net8253)
);

AND2_X1 c7828(
.A1(net8199),
.A2(net7284),
.ZN(net8254)
);

INV_X8 c7829(
.A(net11057),
.ZN(net8255)
);

INV_X16 c7830(
.A(net9841),
.ZN(net8256)
);

NAND2_X1 c7831(
.A1(net8247),
.A2(net8246),
.ZN(net8257)
);

INV_X32 c7832(
.A(net9752),
.ZN(net8258)
);

AND3_X4 c7833(
.A1(net8081),
.A2(net8258),
.A3(net8255),
.ZN(net8259)
);

NAND2_X2 c7834(
.A1(net5364),
.A2(net8219),
.ZN(net8260)
);

NAND3_X2 c7835(
.A1(net7291),
.A2(net7224),
.A3(net11095),
.ZN(net8261)
);

NAND2_X4 c7836(
.A1(net7908),
.A2(net8248),
.ZN(net8262)
);

INV_X4 c7837(
.A(net11006),
.ZN(net8263)
);

AND2_X2 c7838(
.A1(net8161),
.A2(net8254),
.ZN(net8264)
);

XOR2_X1 c7839(
.A(net7294),
.B(net7983),
.Z(net8265)
);

NOR2_X1 c7840(
.A1(net7208),
.A2(net8257),
.ZN(net8266)
);

OR3_X1 c7841(
.A1(net8061),
.A2(net8232),
.A3(net10895),
.ZN(net8267)
);

MUX2_X1 c7842(
.A(net8140),
.B(net7039),
.S(net8123),
.Z(net8268)
);

OAI21_X4 c7843(
.A(net8265),
.B1(net7268),
.B2(net8232),
.ZN(net8269)
);

OR2_X2 c7844(
.A1(net8154),
.A2(net6282),
.ZN(net8270)
);

NOR2_X4 c7845(
.A1(net7334),
.A2(net5033),
.ZN(net8271)
);

MUX2_X2 c7846(
.A(net6358),
.B(net7208),
.S(net3402),
.Z(net8272)
);

SDFFRS_X1 c7847(
.D(net8163),
.RN(net8233),
.SE(net8178),
.SI(net6356),
.SN(net6786),
.CK(clk),
.Q(net8274),
.QN(net8273)
);

NOR2_X2 c7848(
.A1(net6373),
.A2(net8240),
.ZN(net8275)
);

CLKGATETST_X4 c7849(
.E(net8270),
.SE(net8275),
.CK(clk),
.GCK(net8276)
);

AOI222_X1 c7850(
.A1(net8256),
.A2(net8245),
.B1(net7284),
.B2(net8197),
.C1(net8187),
.C2(net7325),
.ZN(net8277)
);

NAND3_X4 c7851(
.A1(net8272),
.A2(net5364),
.A3(net7226),
.ZN(net8278)
);

OR3_X4 c7852(
.A1(net6160),
.A2(net8014),
.A3(net8251),
.ZN(net8279)
);

XOR2_X2 c7853(
.A(net3448),
.B(net10571),
.Z(net8280)
);

XNOR2_X1 c7854(
.A(net8168),
.B(net8121),
.ZN(net8281)
);

AND3_X2 c7855(
.A1(net5389),
.A2(net8240),
.A3(net7131),
.ZN(net8282)
);

NOR3_X1 c7856(
.A1(net8276),
.A2(net8279),
.A3(net11131),
.ZN(net8283)
);

OR2_X4 c7857(
.A1(net8204),
.A2(net10906),
.ZN(net8284)
);

OR2_X1 c7858(
.A1(net8184),
.A2(net11221),
.ZN(net8285)
);

INV_X1 c7859(
.A(net9854),
.ZN(net8286)
);

XNOR2_X2 c7860(
.A(net4127),
.B(net8275),
.ZN(net8287)
);

AOI222_X4 c7861(
.A1(net8251),
.A2(net8284),
.B1(net8254),
.B2(net8232),
.C1(net8197),
.C2(net8111),
.ZN(net8288)
);

AND2_X4 c7862(
.A1(net8243),
.A2(net8255),
.ZN(net8289)
);

OR3_X2 c7863(
.A1(net8061),
.A2(net7038),
.A3(net11222),
.ZN(net8290)
);

OAI21_X2 c7864(
.A(net8264),
.B1(net8238),
.B2(net8240),
.ZN(net8291)
);

INV_X2 c7865(
.A(net10035),
.ZN(net8292)
);

AND2_X1 c7866(
.A1(net8289),
.A2(net7226),
.ZN(net8293)
);

NAND2_X1 c7867(
.A1(net8285),
.A2(net8263),
.ZN(net8294)
);

OAI21_X1 c7868(
.A(net8267),
.B1(net7241),
.B2(net6160),
.ZN(net8295)
);

SDFF_X1 c7869(
.D(net8290),
.SE(net7309),
.SI(net8278),
.CK(clk),
.Q(net8297),
.QN(net8296)
);

AOI21_X2 c7870(
.A(net8271),
.B1(net8267),
.B2(net7211),
.ZN(net8298)
);

AOI21_X1 c7871(
.A(net7254),
.B1(net7241),
.B2(net10545),
.ZN(net8299)
);

AOI21_X4 c7872(
.A(net8294),
.B1(net8238),
.B2(net8296),
.ZN(net8300)
);

SDFF_X2 c7873(
.D(net8287),
.SE(net8293),
.SI(net11221),
.CK(clk),
.Q(net8302),
.QN(net8301)
);

AND3_X1 c7874(
.A1(net7284),
.A2(net8295),
.A3(net8300),
.ZN(net8303)
);

NAND3_X1 c7875(
.A1(net8145),
.A2(net8297),
.A3(net8294),
.ZN(net8304)
);

NOR3_X4 c7876(
.A1(net8034),
.A2(net5035),
.A3(net8059),
.ZN(net8305)
);

NOR3_X2 c7877(
.A1(net7254),
.A2(net8290),
.A3(net11220),
.ZN(net8306)
);

INV_X8 c7878(
.A(net9580),
.ZN(net8307)
);

OAI221_X4 c7879(
.A(net8303),
.B1(net8304),
.B2(net8306),
.C1(net8278),
.C2(net7164),
.ZN(net8308)
);

NAND2_X2 c7880(
.A1(net8307),
.A2(net11095),
.ZN(net8309)
);

NAND2_X4 c7881(
.A1(net8295),
.A2(net8300),
.ZN(net8310)
);

AND3_X4 c7882(
.A1(net6927),
.A2(net6344),
.A3(net8297),
.ZN(net8311)
);

NAND3_X2 c7883(
.A1(net8310),
.A2(net8311),
.A3(net11095),
.ZN(net8312)
);

DFFRS_X1 c7884(
.D(net8275),
.RN(net8311),
.SN(net8312),
.CK(clk),
.Q(net8314),
.QN(net8313)
);

INV_X16 c7885(
.A(net11061),
.ZN(net8315)
);

AND2_X2 c7886(
.A1(net5444),
.A2(net6447),
.ZN(net8316)
);

INV_X32 c7887(
.A(net7164),
.ZN(net8317)
);

INV_X4 c7888(
.A(net10311),
.ZN(net8318)
);

XOR2_X1 c7889(
.A(net5035),
.B(net10967),
.Z(net8319)
);

NOR2_X1 c7890(
.A1(net8258),
.A2(net8209),
.ZN(net8320)
);

INV_X1 c7891(
.A(net9805),
.ZN(net8321)
);

OR2_X2 c7892(
.A1(net5407),
.A2(net8286),
.ZN(net8322)
);

INV_X2 c7893(
.A(net10791),
.ZN(net8323)
);

INV_X8 c7894(
.A(net11022),
.ZN(net8324)
);

INV_X16 c7895(
.A(net7275),
.ZN(net8325)
);

INV_X32 c7896(
.A(net11209),
.ZN(net8326)
);

INV_X4 c7897(
.A(net9743),
.ZN(net8327)
);

NOR2_X4 c7898(
.A1(net6400),
.A2(net8320),
.ZN(net8328)
);

INV_X1 c7899(
.A(net9961),
.ZN(net8329)
);

INV_X2 c7900(
.A(net11135),
.ZN(net8330)
);

NOR2_X2 c7901(
.A1(net8325),
.A2(net7342),
.ZN(net8331)
);

XOR2_X2 c7902(
.A(net8323),
.B(net5444),
.Z(net8332)
);

INV_X8 c7903(
.A(net11135),
.ZN(net8333)
);

XNOR2_X1 c7904(
.A(net8209),
.B(net8327),
.ZN(net8334)
);

OR2_X4 c7905(
.A1(net8321),
.A2(net7226),
.ZN(net8335)
);

INV_X16 c7906(
.A(net10364),
.ZN(net8336)
);

OR2_X1 c7907(
.A1(net7370),
.A2(net8254),
.ZN(net8337)
);

OAI22_X1 c7908(
.A1(net8315),
.A2(net8316),
.B1(net8182),
.B2(net8224),
.ZN(net8338)
);

XNOR2_X2 c7909(
.A(net8239),
.B(net8235),
.ZN(net8339)
);

AND2_X4 c7910(
.A1(net8327),
.A2(net10683),
.ZN(net8340)
);

AND2_X1 c7911(
.A1(net7363),
.A2(net8326),
.ZN(net8341)
);

NAND2_X1 c7912(
.A1(net8309),
.A2(net10774),
.ZN(net8342)
);

NAND2_X2 c7913(
.A1(net6301),
.A2(net7275),
.ZN(net8343)
);

NAND2_X4 c7914(
.A1(net7342),
.A2(net7378),
.ZN(net8344)
);

AND2_X2 c7915(
.A1(net6218),
.A2(net7226),
.ZN(net8345)
);

XOR2_X1 c7916(
.A(net8333),
.B(net5425),
.Z(net8346)
);

INV_X32 c7917(
.A(net10165),
.ZN(net8347)
);

INV_X4 c7918(
.A(net9785),
.ZN(net8348)
);

NOR2_X1 c7919(
.A1(net7131),
.A2(net8341),
.ZN(net8349)
);

OR2_X2 c7920(
.A1(net8032),
.A2(net7353),
.ZN(net8350)
);

OR3_X1 c7921(
.A1(net8336),
.A2(net8346),
.A3(net8337),
.ZN(net8351)
);

NOR2_X4 c7922(
.A1(net8324),
.A2(net8327),
.ZN(net8352)
);

NOR2_X2 c7923(
.A1(net7268),
.A2(net8299),
.ZN(net8353)
);

MUX2_X1 c7924(
.A(net8327),
.B(net8326),
.S(net2570),
.Z(net8354)
);

XOR2_X2 c7925(
.A(net8346),
.B(net7930),
.Z(net8355)
);

XNOR2_X1 c7926(
.A(net8344),
.B(net10449),
.ZN(net8356)
);

OR2_X4 c7927(
.A1(net8318),
.A2(net8345),
.ZN(net8357)
);

AND4_X2 c7928(
.A1(net7406),
.A2(net8345),
.A3(net6395),
.A4(net11209),
.ZN(net8358)
);

OR2_X1 c7929(
.A1(net7356),
.A2(net7226),
.ZN(net8359)
);

INV_X1 c7930(
.A(net8351),
.ZN(net8360)
);

XNOR2_X2 c7931(
.A(net8338),
.B(net8357),
.ZN(net8361)
);

AND2_X4 c7932(
.A1(net8343),
.A2(net8316),
.ZN(net8362)
);

AND2_X1 c7933(
.A1(net7038),
.A2(net10967),
.ZN(net8363)
);

INV_X2 c7934(
.A(net8363),
.ZN(net8364)
);

NAND2_X1 c7935(
.A1(net7822),
.A2(out13),
.ZN(net8365)
);

INV_X8 c7936(
.A(net8362),
.ZN(net8366)
);

NAND2_X2 c7937(
.A1(net7930),
.A2(net8346),
.ZN(net8367)
);

AND4_X1 c7938(
.A1(net8236),
.A2(net8344),
.A3(net8367),
.A4(net7355),
.ZN(net8368)
);

OAI21_X4 c7939(
.A(net6370),
.B1(net8366),
.B2(net8349),
.ZN(net8369)
);

NAND2_X4 c7940(
.A1(net8359),
.A2(net7226),
.ZN(net8370)
);

INV_X16 c7941(
.A(net9849),
.ZN(net8371)
);

AND2_X2 c7942(
.A1(net8250),
.A2(net8214),
.ZN(net8372)
);

DFFRS_X2 c7943(
.D(net8339),
.RN(net8353),
.SN(net8279),
.CK(clk),
.Q(net8374),
.QN(net8373)
);

XOR2_X1 c7944(
.A(net5425),
.B(net8372),
.Z(net8375)
);

NOR2_X1 c7945(
.A1(net8330),
.A2(net8355),
.ZN(net8376)
);

MUX2_X2 c7946(
.A(net5283),
.B(net8357),
.S(net8353),
.Z(net8377)
);

OR2_X2 c7947(
.A1(net6326),
.A2(net7387),
.ZN(net8378)
);

NOR2_X4 c7948(
.A1(net8326),
.A2(net8366),
.ZN(net8379)
);

NAND3_X4 c7949(
.A1(net8367),
.A2(net8349),
.A3(net8342),
.ZN(net8380)
);

NOR2_X2 c7950(
.A1(net8350),
.A2(net8189),
.ZN(net8381)
);

XOR2_X2 c7951(
.A(net8355),
.B(net7356),
.Z(net8382)
);

SDFFS_X1 c7952(
.D(net8366),
.SE(net8379),
.SI(net8370),
.SN(net7363),
.CK(clk),
.Q(net8384),
.QN(net8383)
);

OR3_X4 c7953(
.A1(net8352),
.A2(net8365),
.A3(net8329),
.ZN(net8385)
);

AND3_X2 c7954(
.A1(net8380),
.A2(net8385),
.A3(net8383),
.ZN(net8386)
);

INV_X32 c7955(
.A(net11094),
.ZN(net8387)
);

NOR3_X1 c7956(
.A1(net8384),
.A2(net8347),
.A3(net8380),
.ZN(net8388)
);

AOI22_X4 c7957(
.A1(net8268),
.A2(net8381),
.B1(net8386),
.B2(net7357),
.ZN(net8389)
);

OR3_X2 c7958(
.A1(net7377),
.A2(net8365),
.A3(net8384),
.ZN(net8390)
);

SDFF_X1 c7959(
.D(net8360),
.SE(net6337),
.SI(net8385),
.CK(clk),
.Q(net8392),
.QN(net8391)
);

SDFF_X2 c7960(
.D(net2570),
.SE(net8392),
.SI(net8111),
.CK(clk),
.Q(net8394),
.QN(net8393)
);

OAI21_X2 c7961(
.A(net8375),
.B1(net8394),
.B2(net8391),
.ZN(net8395)
);

OAI21_X1 c7962(
.A(net7269),
.B1(net8387),
.B2(net8393),
.ZN(net8396)
);

OAI33_X1 c7963(
.A1(net8364),
.A2(net8383),
.A3(net8248),
.B1(net5474),
.B2(net6369),
.B3(net10819),
.ZN(net8397)
);

SDFFRS_X2 c7964(
.D(net8320),
.RN(net8388),
.SE(net8379),
.SI(net7268),
.SN(net11224),
.CK(clk),
.Q(net8399),
.QN(net8398)
);

OAI22_X4 c7965(
.A1(net8356),
.A2(net8350),
.B1(net8391),
.B2(net11224),
.ZN(net8400)
);

AOI22_X2 c7966(
.A1(net8386),
.A2(net8348),
.B1(net10544),
.B2(net11224),
.ZN(net8401)
);

AOI21_X2 c7967(
.A(net8385),
.B1(net10724),
.B2(net10952),
.ZN(net8402)
);

INV_X4 c7968(
.A(net11050),
.ZN(net8403)
);

NAND4_X4 c7969(
.A1(net6460),
.A2(net8248),
.A3(net7500),
.A4(net7471),
.ZN(net8404)
);

AOI21_X1 c7970(
.A(net6253),
.B1(net7447),
.B2(net8316),
.ZN(net8405)
);

INV_X1 c7971(
.A(net11092),
.ZN(net8406)
);

XNOR2_X1 c7972(
.A(net8254),
.B(net6342),
.ZN(net8407)
);

OR2_X4 c7973(
.A1(net7518),
.A2(net7475),
.ZN(net8408)
);

OR2_X1 c7974(
.A1(net8266),
.A2(net8407),
.ZN(net8409)
);

XNOR2_X2 c7975(
.A(net7501),
.B(net11225),
.ZN(net8410)
);

AOI21_X4 c7976(
.A(net8382),
.B1(net8409),
.B2(net7353),
.ZN(net8411)
);

AND2_X4 c7977(
.A1(net8406),
.A2(net8331),
.ZN(net8412)
);

AND3_X1 c7978(
.A1(net5544),
.A2(net6476),
.A3(net7367),
.ZN(net8413)
);

AND2_X1 c7979(
.A1(net7378),
.A2(net8313),
.ZN(net8414)
);

NAND2_X1 c7980(
.A1(net8348),
.A2(net8372),
.ZN(net8415)
);

NAND3_X1 c7981(
.A1(net8342),
.A2(net8309),
.A3(net7509),
.ZN(net8416)
);

NOR3_X4 c7982(
.A1(net7512),
.A2(net8409),
.A3(net7326),
.ZN(net8417)
);

INV_X2 c7983(
.A(net9904),
.ZN(net8418)
);

INV_X8 c7984(
.A(net9918),
.ZN(net8419)
);

DFFRS_X1 c7985(
.D(net7502),
.RN(net8408),
.SN(net8407),
.CK(clk),
.Q(net8421),
.QN(net8420)
);

NAND2_X2 c7986(
.A1(net7442),
.A2(net8409),
.ZN(net8422)
);

NAND2_X4 c7987(
.A1(net8417),
.A2(net10427),
.ZN(net8423)
);

NOR3_X2 c7988(
.A1(net8414),
.A2(net8373),
.A3(net7473),
.ZN(net8424)
);

AND3_X4 c7989(
.A1(net1709),
.A2(net8422),
.A3(net11221),
.ZN(net8425)
);

NAND3_X2 c7990(
.A1(net8402),
.A2(net5551),
.A3(net11223),
.ZN(net8426)
);

INV_X16 c7991(
.A(net9806),
.ZN(net8427)
);

INV_X32 c7992(
.A(net9744),
.ZN(net8428)
);

AND2_X2 c7993(
.A1(net8340),
.A2(net8407),
.ZN(net8429)
);

OR3_X1 c7994(
.A1(net6342),
.A2(net8411),
.A3(net8420),
.ZN(net8430)
);

INV_X4 c7995(
.A(net9902),
.ZN(net8431)
);

DFFRS_X2 c7996(
.D(net7483),
.RN(net8430),
.SN(net8423),
.CK(clk),
.Q(net8433),
.QN(net8432)
);

XOR2_X1 c7997(
.A(net6472),
.B(net8225),
.Z(net8434)
);

NOR2_X1 c7998(
.A1(net7367),
.A2(net8429),
.ZN(net8435)
);

SDFF_X1 c7999(
.D(net8427),
.SE(net8424),
.SI(net8429),
.CK(clk),
.Q(net8437),
.QN(net8436)
);

INV_X1 c8000(
.A(net9692),
.ZN(net8438)
);

MUX2_X1 c8001(
.A(net7455),
.B(net8434),
.S(net7429),
.Z(net8439)
);

OR2_X2 c8002(
.A1(net6316),
.A2(net8419),
.ZN(net8440)
);

NOR2_X4 c8003(
.A1(net7426),
.A2(net8418),
.ZN(net8441)
);

OAI21_X4 c8004(
.A(net8431),
.B1(net6342),
.B2(net7458),
.ZN(net8442)
);

MUX2_X2 c8005(
.A(net7433),
.B(net6518),
.S(net8316),
.Z(net8443)
);

NOR2_X2 c8006(
.A1(net7039),
.A2(net7447),
.ZN(net8444)
);

SDFF_X2 c8007(
.D(net7429),
.SE(net8434),
.SI(net8379),
.CK(clk),
.Q(net8446),
.QN(net8445)
);

NAND3_X4 c8008(
.A1(net4329),
.A2(net8419),
.A3(net7326),
.ZN(net8447)
);

XOR2_X2 c8009(
.A(net8413),
.B(net7453),
.Z(net8448)
);

OR3_X4 c8010(
.A1(net8442),
.A2(net8316),
.A3(net8443),
.ZN(net8449)
);

OAI211_X2 c8011(
.A(net8438),
.B(net4540),
.C1(net8436),
.C2(net11220),
.ZN(net8450)
);

INV_X2 c8012(
.A(net11119),
.ZN(net8451)
);

XNOR2_X1 c8013(
.A(net8444),
.B(net8446),
.ZN(net8452)
);

OR2_X4 c8014(
.A1(net8452),
.A2(net8342),
.ZN(net8453)
);

AND3_X2 c8015(
.A1(net8440),
.A2(net8429),
.A3(net8443),
.ZN(net8454)
);

OR4_X2 c8016(
.A1(net8402),
.A2(net8453),
.A3(net8443),
.A4(net8418),
.ZN(net8455)
);

NOR3_X1 c8017(
.A1(net4540),
.A2(net8432),
.A3(net2674),
.ZN(net8456)
);

SDFFRS_X1 c8018(
.D(net8329),
.RN(net7822),
.SE(net8454),
.SI(net8429),
.SN(net8278),
.CK(clk),
.Q(net8458),
.QN(net8457)
);

OR3_X2 c8019(
.A1(net8276),
.A2(net8456),
.A3(net8445),
.ZN(net8459)
);

AOI211_X1 c8020(
.A(net8421),
.B(net6342),
.C1(net5474),
.C2(net10450),
.ZN(net8460)
);

OAI21_X2 c8021(
.A(net8281),
.B1(net8451),
.B2(net8454),
.ZN(net8461)
);

OAI21_X1 c8022(
.A(net8189),
.B1(net8458),
.B2(net7361),
.ZN(net8462)
);

DFFRS_X1 c8023(
.D(net8379),
.RN(net8453),
.SN(net7500),
.CK(clk),
.Q(net8464),
.QN(net8463)
);

OAI221_X2 c8024(
.A(net8449),
.B1(net8379),
.B2(net8393),
.C1(net10910),
.C2(net11210),
.ZN(net8465)
);

AOI21_X2 c8025(
.A(net6469),
.B1(net7353),
.B2(net10886),
.ZN(net8466)
);

DFFRS_X2 c8026(
.D(net8441),
.RN(net8456),
.SN(net7724),
.CK(clk),
.Q(net8468),
.QN(net8467)
);

AOI21_X1 c8027(
.A(net7354),
.B1(net6469),
.B2(net8463),
.ZN(net8469)
);

AOI21_X4 c8028(
.A(net8468),
.B1(net8429),
.B2(net8450),
.ZN(net8470)
);

AOI221_X4 c8029(
.A(net5549),
.B1(net8278),
.B2(net8457),
.C1(net7918),
.C2(net8255),
.ZN(net8471)
);

AND3_X1 c8030(
.A1(net7353),
.A2(net8464),
.A3(net10961),
.ZN(net8472)
);

OR2_X1 c8031(
.A1(net8451),
.A2(net8266),
.ZN(net8473)
);

NAND3_X1 c8032(
.A1(net8464),
.A2(net4534),
.A3(net10549),
.ZN(net8474)
);

NOR3_X4 c8033(
.A1(net6518),
.A2(net8423),
.A3(net5315),
.ZN(net8475)
);

NOR3_X2 c8034(
.A1(net8472),
.A2(net8278),
.A3(net8470),
.ZN(net8476)
);

SDFF_X1 c8035(
.D(net8337),
.SE(net7492),
.SI(net8111),
.CK(clk),
.Q(net8478),
.QN(net8477)
);

AND3_X4 c8036(
.A1(net8461),
.A2(net8415),
.A3(net8429),
.ZN(net8479)
);

NAND4_X2 c8037(
.A1(net8433),
.A2(net8447),
.A3(net3565),
.A4(net8457),
.ZN(net8480)
);

INV_X8 c8038(
.A(net11092),
.ZN(net8481)
);

NAND3_X2 c8039(
.A1(net8437),
.A2(net8313),
.A3(net10417),
.ZN(net8482)
);

XNOR2_X2 c8040(
.A(net10839),
.B(net10911),
.ZN(net8483)
);

SDFF_X2 c8041(
.D(net8403),
.SE(net8480),
.SI(net8378),
.CK(clk),
.Q(net8485),
.QN(net8484)
);

AND2_X4 c8042(
.A1(net8428),
.A2(net10416),
.ZN(net8486)
);

OR3_X1 c8043(
.A1(net8473),
.A2(net8481),
.A3(net8482),
.ZN(net8487)
);

MUX2_X1 c8044(
.A(net8487),
.B(net8482),
.S(net8441),
.Z(net8488)
);

OAI21_X4 c8045(
.A(net8483),
.B1(net8418),
.B2(net10723),
.ZN(net8489)
);

MUX2_X2 c8046(
.A(net8466),
.B(net8483),
.S(net10922),
.Z(net8490)
);

NAND3_X4 c8047(
.A1(net7361),
.A2(net8489),
.A3(net8488),
.ZN(net8491)
);

OR3_X4 c8048(
.A1(net8484),
.A2(net10588),
.A3(net10881),
.ZN(net8492)
);

DFFRS_X1 c8049(
.D(net7499),
.RN(net8486),
.SN(net8467),
.CK(clk),
.Q(net8494),
.QN(net8493)
);

AOI222_X2 c8050(
.A1(net8485),
.A2(net8492),
.B1(net8494),
.B2(net8457),
.C1(net8255),
.C2(net8420),
.ZN(net8495)
);

AND2_X1 c8051(
.A1(net8299),
.A2(net8454),
.ZN(net8496)
);

NAND2_X1 c8052(
.A1(net8396),
.A2(net2712),
.ZN(net8497)
);

NAND2_X2 c8053(
.A1(net3576),
.A2(out25),
.ZN(net8498)
);

AND3_X2 c8054(
.A1(net828),
.A2(net8392),
.A3(net7271),
.ZN(net8499)
);

DFFRS_X2 c8055(
.D(net8279),
.RN(net8232),
.SN(net5315),
.CK(clk),
.Q(net8501),
.QN(net8500)
);

NAND2_X4 c8056(
.A1(net5613),
.A2(net7539),
.ZN(net8502)
);

NOR3_X1 c8057(
.A1(net8248),
.A2(net4689),
.A3(net6607),
.ZN(net8503)
);

SDFF_X1 c8058(
.D(net8422),
.SE(net7586),
.SI(net5411),
.CK(clk),
.Q(net8505),
.QN(net8504)
);

OR3_X2 c8059(
.A1(net7539),
.A2(net6600),
.A3(net7585),
.ZN(net8506)
);

OAI21_X2 c8060(
.A(net8506),
.B1(net8458),
.B2(net2570),
.ZN(net8507)
);

AOI221_X2 c8061(
.A(net7471),
.B1(net8504),
.B2(net7539),
.C1(net6426),
.C2(net7489),
.ZN(net8508)
);

SDFF_X2 c8062(
.D(net8214),
.SE(net7271),
.SI(net8394),
.CK(clk),
.Q(net8510),
.QN(net8509)
);

AND2_X2 c8063(
.A1(net5381),
.A2(net1708),
.ZN(net8511)
);

OAI21_X1 c8064(
.A(net7576),
.B1(net7471),
.B2(net7552),
.ZN(net8512)
);

AOI21_X2 c8065(
.A(net3691),
.B1(out25),
.B2(net3403),
.ZN(net8513)
);

XOR2_X1 c8066(
.A(net8374),
.B(net8450),
.Z(net8514)
);

AOI21_X1 c8067(
.A(net8508),
.B1(net5632),
.B2(net11225),
.ZN(net8515)
);

INV_X16 c8068(
.A(net11050),
.ZN(net8516)
);

DFFRS_X1 c8069(
.D(net7600),
.RN(net8500),
.SN(net8511),
.CK(clk),
.Q(net8518),
.QN(net8517)
);

DFFRS_X2 c8070(
.D(net7472),
.RN(net7602),
.SN(net7605),
.CK(clk),
.Q(net8520),
.QN(net8519)
);

AOI21_X4 c8071(
.A(net6607),
.B1(net8491),
.B2(net7585),
.ZN(net8521)
);

AOI221_X1 c8072(
.A(net7607),
.B1(net8422),
.B2(net8474),
.C1(net8232),
.C2(net8509),
.ZN(net8522)
);

SDFF_X1 c8073(
.D(net7453),
.SE(net8418),
.SI(net8415),
.CK(clk),
.Q(net8524),
.QN(net8523)
);

OR4_X4 c8074(
.A1(net6597),
.A2(net4476),
.A3(net7271),
.A4(net8509),
.ZN(net8525)
);

AND3_X1 c8075(
.A1(net3698),
.A2(net8517),
.A3(net8520),
.ZN(net8526)
);

NAND3_X1 c8076(
.A1(net8506),
.A2(net5381),
.A3(net10948),
.ZN(net8527)
);

SDFF_X2 c8077(
.D(net5411),
.SE(net5632),
.SI(net3691),
.CK(clk),
.Q(net8529),
.QN(net8528)
);

NOR3_X4 c8078(
.A1(net8371),
.A2(net8422),
.A3(net3698),
.ZN(net8530)
);

NOR2_X1 c8079(
.A1(net7604),
.A2(net8182),
.ZN(net8531)
);

NOR3_X2 c8080(
.A1(net7360),
.A2(net8505),
.A3(net8529),
.ZN(net8532)
);

AND3_X4 c8081(
.A1(net8385),
.A2(net7123),
.A3(net10656),
.ZN(net8533)
);

NAND3_X2 c8082(
.A1(net7552),
.A2(net8511),
.A3(net8474),
.ZN(net8534)
);

OR3_X1 c8083(
.A1(net7585),
.A2(net8469),
.A3(net8385),
.ZN(net8535)
);

MUX2_X1 c8084(
.A(net8418),
.B(net8520),
.S(net8524),
.Z(net8536)
);

OR2_X2 c8085(
.A1(net7573),
.A2(net11103),
.ZN(net8537)
);

OAI21_X4 c8086(
.A(net6476),
.B1(net8394),
.B2(net6477),
.ZN(net8538)
);

MUX2_X2 c8087(
.A(net6426),
.B(net8537),
.S(net8520),
.Z(net8539)
);

INV_X32 c8088(
.A(net9616),
.ZN(net8540)
);

NAND3_X4 c8089(
.A1(net8539),
.A2(net8537),
.A3(net8470),
.ZN(net8541)
);

OR3_X4 c8090(
.A1(net8497),
.A2(net7452),
.A3(net8536),
.ZN(net8542)
);

INV_X4 c8091(
.A(net9715),
.ZN(net8543)
);

OAI222_X1 c8092(
.A1(net5613),
.A2(net7489),
.B1(net8511),
.B2(net8519),
.C1(net10832),
.C2(net10970),
.ZN(net8544)
);

AND3_X2 c8093(
.A1(net6634),
.A2(net8518),
.A3(net2737),
.ZN(net8545)
);

NOR3_X1 c8094(
.A1(net8235),
.A2(net8510),
.A3(net8497),
.ZN(net8546)
);

OR3_X2 c8095(
.A1(net8398),
.A2(net8497),
.A3(net10541),
.ZN(net8547)
);

OAI21_X2 c8096(
.A(net4528),
.B1(net3698),
.B2(net8509),
.ZN(net8548)
);

DFFRS_X1 c8097(
.D(net8540),
.RN(net7605),
.SN(net10742),
.CK(clk),
.Q(net8550),
.QN(net8549)
);

OAI21_X1 c8098(
.A(net8510),
.B1(net6597),
.B2(net8519),
.ZN(net8551)
);

AOI21_X2 c8099(
.A(net4689),
.B1(net8514),
.B2(net8536),
.ZN(net8552)
);

AOI21_X1 c8100(
.A(net6586),
.B1(net6633),
.B2(net10618),
.ZN(net8553)
);

AOI21_X4 c8101(
.A(net8456),
.B1(net8533),
.B2(net8548),
.ZN(net8554)
);

AND3_X1 c8102(
.A1(net7540),
.A2(net8543),
.A3(net8524),
.ZN(net8555)
);

OAI221_X1 c8103(
.A(net6600),
.B1(net8543),
.B2(net8497),
.C1(net7586),
.C2(net6467),
.ZN(net8556)
);

NAND3_X1 c8104(
.A1(net6467),
.A2(net8550),
.A3(net8497),
.ZN(net8557)
);

NOR3_X4 c8105(
.A1(net6477),
.A2(net8531),
.A3(net8548),
.ZN(net8558)
);

OAI22_X2 c8106(
.A1(net8509),
.A2(net8528),
.B1(net10924),
.B2(net10929),
.ZN(net8559)
);

NOR3_X2 c8107(
.A1(net8559),
.A2(net8552),
.A3(net8548),
.ZN(net8560)
);

NOR2_X4 c8108(
.A1(net8553),
.A2(net8560),
.ZN(net8561)
);

AND3_X4 c8109(
.A1(net8232),
.A2(net8520),
.A3(net6633),
.ZN(net8562)
);

NAND3_X2 c8110(
.A1(net8548),
.A2(net8536),
.A3(net8513),
.ZN(net8563)
);

OR3_X1 c8111(
.A1(net7586),
.A2(net8556),
.A3(net8562),
.ZN(net8564)
);

OAI211_X4 c8112(
.A(net6600),
.B(net8510),
.C1(net10618),
.C2(net11103),
.ZN(net8565)
);

MUX2_X1 c8113(
.A(net8470),
.B(net8564),
.S(net8510),
.Z(net8566)
);

OAI21_X4 c8114(
.A(net8454),
.B1(net8563),
.B2(net8561),
.ZN(net8567)
);

NOR2_X2 c8115(
.A1(net8562),
.A2(net10702),
.ZN(net8568)
);

MUX2_X2 c8116(
.A(net8309),
.B(net8537),
.S(net8548),
.Z(net8569)
);

XOR2_X2 c8117(
.A(net8569),
.B(net8541),
.Z(net8570)
);

NAND3_X4 c8118(
.A1(net8249),
.A2(net8570),
.A3(net8392),
.ZN(net8571)
);

OR3_X4 c8119(
.A1(net8557),
.A2(net8448),
.A3(net8549),
.ZN(net8572)
);

DFFRS_X2 c8120(
.D(net7387),
.RN(net8458),
.SN(net8567),
.CK(clk),
.Q(net8574),
.QN(net8573)
);

AND3_X2 c8121(
.A1(net8551),
.A2(net8478),
.A3(net10725),
.ZN(net8575)
);

NOR3_X1 c8122(
.A1(net8561),
.A2(net8497),
.A3(net10541),
.ZN(net8576)
);

OR3_X2 c8123(
.A1(net8415),
.A2(net8546),
.A3(net8545),
.ZN(net8577)
);

SDFF_X1 c8124(
.D(net7579),
.SE(net7605),
.SI(net11107),
.CK(clk),
.Q(net8579),
.QN(net8578)
);

OAI21_X2 c8125(
.A(net8555),
.B1(net8575),
.B2(net8551),
.ZN(net8580)
);

OAI21_X1 c8126(
.A(net8580),
.B1(net6633),
.B2(net3691),
.ZN(net8581)
);

INV_X1 c8127(
.A(net9615),
.ZN(net8582)
);

AOI21_X2 c8128(
.A(net7585),
.B1(net10550),
.B2(net10655),
.ZN(net8583)
);

AOI21_X1 c8129(
.A(net7424),
.B1(net8545),
.B2(net8583),
.ZN(net8584)
);

AOI21_X4 c8130(
.A(net8565),
.B1(net7605),
.B2(net8572),
.ZN(net8585)
);

AND3_X1 c8131(
.A1(net8532),
.A2(net8581),
.A3(net8548),
.ZN(net8586)
);

NAND3_X1 c8132(
.A1(net8450),
.A2(net8529),
.A3(net10966),
.ZN(net8587)
);

NOR3_X4 c8133(
.A1(net8586),
.A2(net8511),
.A3(net10877),
.ZN(net8588)
);

OAI211_X1 c8160(
.A(net6690),
.B(net4728),
.C1(out3),
.C2(net5719),
.ZN(net8589)
);

SDFF_X2 c8161(
.D(net8511),
.SE(net8314),
.SI(net8629),
.CK(clk),
.Q(net8591),
.QN(net8590)
);

NOR4_X4 c8162(
.A1(net7690),
.A2(net8579),
.A3(net6697),
.A4(net8634),
.ZN(net8592)
);

NOR3_X2 c8163(
.A1(net7458),
.A2(net8591),
.A3(net8631),
.ZN(net8593)
);

INV_X2 c8164(
.A(net11237),
.ZN(out6)
);

NOR4_X2 c8165(
.A1(net6525),
.A2(net6719),
.A3(net5723),
.A4(net8511),
.ZN(net8594)
);

AOI211_X4 c8166(
.A(net7632),
.B(net7699),
.C1(net8622),
.C2(net10982),
.ZN(net8595)
);

NOR4_X1 c8167(
.A1(net7666),
.A2(net7545),
.A3(net8631),
.A4(net10382),
.ZN(net8596)
);

AND3_X4 c8168(
.A1(net8591),
.A2(net8622),
.A3(net10991),
.ZN(net8597)
);

NAND3_X2 c8169(
.A1(net8595),
.A2(net8597),
.A3(net8542),
.ZN(net8598)
);

OR3_X1 c8170(
.A1(net5723),
.A2(net7682),
.A3(net8622),
.ZN(net8599)
);

MUX2_X1 c8171(
.A(net8469),
.B(net8597),
.S(net8635),
.Z(net8600)
);

SDFFS_X2 c8172(
.D(net8630),
.SE(net8628),
.SI(net6718),
.SN(net8637),
.CK(clk),
.Q(net8602),
.QN(net8601)
);

OAI21_X4 c8173(
.A(net8478),
.B1(net8579),
.B2(net7699),
.ZN(net8603)
);

MUX2_X2 c8174(
.A(net5670),
.B(net7494),
.S(net8637),
.Z(net8604)
);

NAND3_X4 c8175(
.A1(net5509),
.A2(net7494),
.A3(net8624),
.ZN(out20)
);

OAI221_X4 c8176(
.A(net8599),
.B1(net8635),
.B2(net8590),
.C1(net8622),
.C2(net8511),
.ZN(net8605)
);

OR3_X4 c8177(
.A1(net6561),
.A2(net8637),
.A3(net5743),
.ZN(net8606)
);

AND3_X2 c8178(
.A1(net8474),
.A2(net8642),
.A3(net8589),
.ZN(net8607)
);

NOR3_X1 c8179(
.A1(net8621),
.A2(net8601),
.A3(net10981),
.ZN(out21)
);

OR3_X2 c8180(
.A1(net8638),
.A2(net7639),
.A3(net8639),
.ZN(net8608)
);

OAI21_X2 c8181(
.A(net8622),
.B1(net8593),
.B2(net8591),
.ZN(net8609)
);

OAI21_X1 c8182(
.A(net8589),
.B1(net8602),
.B2(net7458),
.ZN(out11)
);

AOI21_X2 c8183(
.A(net2851),
.B1(net7678),
.B2(net10768),
.ZN(net8610)
);

DFFRS_X1 c8184(
.D(net8491),
.RN(net8607),
.SN(net10991),
.CK(clk),
.Q(out17),
.QN(net8611)
);

OAI221_X2 c8185(
.A(net8627),
.B1(net7651),
.B2(net8477),
.C1(net6721),
.ZN(net11000)
);

OAI222_X4 c8186(
.A1(net8629),
.A2(net8592),
.B1(net8590),
.B2(net8611),
.C1(out25),
.C2(net7545),
.ZN(net8613)
);

AOI211_X2 c8187(
.A(net8603),
.B(out17),
.C1(out1),
.C2(out23),
.ZN(net8614)
);

AOI221_X4 c8188(
.A(net4727),
.B1(net8611),
.B2(net8637),
.C1(net10832),
.C2(net10888),
.ZN(net8615)
);

OAI222_X2 c8189(
.A1(net6697),
.A2(net8608),
.B1(net8637),
.B2(out17),
.C1(net5632),
.C2(net8574),
.ZN(net8616)
);

AOI222_X1 c8190(
.A1(net7598),
.A2(net8596),
.B1(net8634),
.B2(net7682),
.C1(net8622),
.C2(net11011),
.ZN(net8617)
);

AOI21_X1 c8191(
.A(net8631),
.B1(net5720),
.B2(net10382),
.ZN(out18)
);

AOI21_X4 c8192(
.A(out18),
.B1(net10892),
.B2(net11061),
.ZN(net8618)
);

AND3_X1 c8193(
.A1(net6650),
.A2(net7694),
.A3(net5632),
.ZN(net8619)
);

DFFRS_X2 c8194(
.D(net7644),
.RN(net7699),
.SN(out16),
.CK(clk),
.Q(net8621),
.QN(net8620)
);

NAND3_X1 c8195(
.A1(net4728),
.A2(net7666),
.A3(net8488),
.ZN(out24)
);

NOR3_X4 c8196(
.A1(net7588),
.A2(net7625),
.A3(net8620),
.ZN(net8622)
);

NOR3_X2 c8197(
.A1(net7545),
.A2(net8542),
.A3(net5720),
.ZN(net8623)
);

SDFF_X1 c8198(
.D(net7612),
.SE(net5632),
.SI(net2851),
.CK(clk),
.Q(net8625),
.QN(net8624)
);

AND3_X4 c8199(
.A1(net6646),
.A2(out9),
.A3(net6561),
.ZN(net8626)
);

NAND3_X2 c8200(
.A1(net8626),
.A2(net4789),
.A3(net8477),
.ZN(net8627)
);

AOI22_X1 c8201(
.A1(net7667),
.A2(net8625),
.B1(net8542),
.B2(out9),
.ZN(net8628)
);

OR3_X1 c8202(
.A1(net7639),
.A2(net8623),
.A3(net8622),
.ZN(net8629)
);

MUX2_X1 c8203(
.A(net7582),
.B(net7632),
.S(net5632),
.Z(net8630)
);

OAI21_X4 c8204(
.A(net5743),
.B1(net6690),
.B2(net7545),
.ZN(net8631)
);

AND4_X4 c8205(
.A1(net6684),
.A2(net6561),
.A3(net8631),
.A4(net10769),
.ZN(out22)
);

MUX2_X2 c8206(
.A(net2849),
.B(net6721),
.S(net7699),
.Z(net8632)
);

NAND4_X1 c8207(
.A1(net8498),
.A2(net7678),
.A3(net7682),
.A4(net6561),
.ZN(net8633)
);

SDFF_X2 c8208(
.D(net7696),
.SE(net7553),
.SI(net7693),
.CK(clk),
.Q(net8635),
.QN(net8634)
);

NAND3_X4 c8209(
.A1(net6652),
.A2(net6525),
.A3(net8578),
.ZN(out14)
);

OR3_X4 c8210(
.A1(net8488),
.A2(net8511),
.A3(net4727),
.ZN(net8636)
);

AND3_X2 c8211(
.A1(net7691),
.A2(net8631),
.A3(net7632),
.ZN(net8637)
);

NOR3_X1 c8212(
.A1(net5720),
.A2(net4789),
.A3(net10720),
.ZN(net8638)
);

DFFRS_X1 c8213(
.D(net8633),
.RN(net8635),
.SN(net7494),
.CK(clk),
.Q(net8640),
.QN(net8639)
);

OR3_X2 c8214(
.A1(net7651),
.A2(net8640),
.A3(net8637),
.ZN(net8641)
);

OAI21_X2 c8215(
.A(net8314),
.B1(net7588),
.B2(net10943),
.ZN(out12)
);

INV_X8 c8216(
.A(net11236),
.ZN(net8642)
);

INV_X16 c8217(
.A(net7783),
.ZN(net8643)
);

INV_X32 c8218(
.A(net9660),
.ZN(net8644)
);

XNOR2_X1 c8219(
.A(net4798),
.B(net7747),
.ZN(net8645)
);

INV_X4 c8220(
.A(net8643),
.ZN(net8646)
);

INV_X1 c8221(
.A(net7759),
.ZN(net8647)
);

INV_X2 c8222(
.A(net8644),
.ZN(net8648)
);

INV_X8 c8223(
.A(net6815),
.ZN(net8649)
);

INV_X16 c8224(
.A(net7783),
.ZN(net8650)
);

OR2_X4 c8225(
.A1(net5818),
.A2(net6789),
.ZN(net8651)
);

INV_X32 c8226(
.A(net6755),
.ZN(net8652)
);

INV_X4 c8227(
.A(net7755),
.ZN(net8653)
);

INV_X1 c8228(
.A(net8644),
.ZN(net8654)
);

OAI21_X1 c8229(
.A(net4865),
.B1(net8650),
.B2(net7712),
.ZN(net8655)
);

OR2_X1 c8230(
.A1(net6799),
.A2(net7783),
.ZN(net8656)
);

INV_X2 c8231(
.A(net5837),
.ZN(net8657)
);

INV_X8 c8232(
.A(net8657),
.ZN(net8658)
);

INV_X16 c8233(
.A(net8650),
.ZN(net8659)
);

INV_X32 c8234(
.A(net9660),
.ZN(net8660)
);

INV_X4 c8235(
.A(net7740),
.ZN(net8661)
);

INV_X1 c8236(
.A(net8650),
.ZN(net8662)
);

INV_X2 c8237(
.A(net8648),
.ZN(net8663)
);

INV_X8 c8238(
.A(net7747),
.ZN(net8664)
);

INV_X16 c8239(
.A(net7792),
.ZN(net8665)
);

XNOR2_X2 c8240(
.A(net8652),
.B(net7731),
.ZN(net8666)
);

AND2_X4 c8241(
.A1(net8657),
.A2(net8666),
.ZN(net8667)
);

INV_X32 c8242(
.A(net8667),
.ZN(net8668)
);

INV_X4 c8243(
.A(net8666),
.ZN(net8669)
);

INV_X1 c8244(
.A(net8647),
.ZN(net8670)
);

INV_X2 c8245(
.A(net7761),
.ZN(net8671)
);

CLKGATETST_X8 c8246(
.E(net5808),
.SE(net8655),
.CK(clk),
.GCK(net8672)
);

INV_X8 c8247(
.A(net5767),
.ZN(net8673)
);

INV_X16 c8248(
.A(net8659),
.ZN(net8674)
);

INV_X32 c8249(
.A(net6809),
.ZN(net8675)
);

INV_X4 c8250(
.A(net8646),
.ZN(net8676)
);

INV_X1 c8251(
.A(net7739),
.ZN(net8677)
);

INV_X2 c8252(
.A(net9720),
.ZN(net8678)
);

INV_X8 c8253(
.A(net8672),
.ZN(net8679)
);

INV_X16 c8254(
.A(net8669),
.ZN(net8680)
);

INV_X32 c8255(
.A(net8678),
.ZN(net8681)
);

AND2_X1 c8256(
.A1(net8677),
.A2(net8665),
.ZN(net8682)
);

NAND2_X1 c8257(
.A1(net8676),
.A2(net8666),
.ZN(net8683)
);

NAND2_X2 c8258(
.A1(net8671),
.A2(net8651),
.ZN(net8684)
);

NAND2_X4 c8259(
.A1(net8659),
.A2(net8681),
.ZN(net8685)
);

AND2_X2 c8260(
.A1(net8683),
.A2(net8653),
.ZN(net8686)
);

INV_X4 c8261(
.A(net8682),
.ZN(net8687)
);

XOR2_X1 c8262(
.A(net7754),
.B(net8671),
.Z(net8688)
);

INV_X1 c8263(
.A(net7784),
.ZN(net8689)
);

NOR2_X1 c8264(
.A1(net8674),
.A2(net7783),
.ZN(net8690)
);

INV_X2 c8265(
.A(net8681),
.ZN(net8691)
);

OR2_X2 c8266(
.A1(net8660),
.A2(net8688),
.ZN(net8692)
);

INV_X8 c8267(
.A(net8691),
.ZN(net8693)
);

NOR2_X4 c8268(
.A1(net8674),
.A2(net8654),
.ZN(net8694)
);

NOR2_X2 c8269(
.A1(net8694),
.A2(net8681),
.ZN(net8695)
);

INV_X16 c8270(
.A(net8663),
.ZN(net8696)
);

XOR2_X2 c8271(
.A(net8686),
.B(net8682),
.Z(net8697)
);

XNOR2_X1 c8272(
.A(net8668),
.B(net8697),
.ZN(net8698)
);

OR2_X4 c8273(
.A1(net6789),
.A2(net8687),
.ZN(net8699)
);

AOI21_X2 c8274(
.A(net8661),
.B1(net8678),
.B2(net8687),
.ZN(net8700)
);

OR2_X1 c8275(
.A1(net8645),
.A2(net8697),
.ZN(net8701)
);

XNOR2_X2 c8276(
.A(net8665),
.B(net8651),
.ZN(net8702)
);

AND2_X4 c8277(
.A1(net8688),
.A2(net8678),
.ZN(net8703)
);

AND2_X1 c8278(
.A1(net8703),
.A2(net8692),
.ZN(net8704)
);

NAND2_X1 c8279(
.A1(net8679),
.A2(net6789),
.ZN(net8705)
);

NAND2_X2 c8280(
.A1(net8683),
.A2(net8691),
.ZN(net8706)
);

NAND2_X4 c8281(
.A1(net8704),
.A2(net8705),
.ZN(net8707)
);

OR4_X1 c8282(
.A1(net8695),
.A2(net8703),
.A3(net8705),
.A4(net8670),
.ZN(net8708)
);

AND2_X2 c8283(
.A1(net8656),
.A2(net8707),
.ZN(net8709)
);

OAI22_X1 c8284(
.A1(net8709),
.A2(net8707),
.B1(net7784),
.B2(net8705),
.ZN(net8710)
);

SDFFR_X1 c8285(
.D(net8698),
.RN(net7761),
.SE(net7728),
.SI(net8687),
.CK(clk),
.Q(net8712),
.QN(net8711)
);

AOI21_X1 c8286(
.A(net8675),
.B1(net8711),
.B2(net5822),
.ZN(net8713)
);

AOI21_X4 c8287(
.A(net8706),
.B1(net8700),
.B2(net8692),
.ZN(net8714)
);

DFFRS_X2 c8288(
.D(net8672),
.RN(net8707),
.SN(net8708),
.CK(clk),
.Q(net8716),
.QN(net8715)
);

SDFF_X1 c8289(
.D(net8699),
.SE(net8698),
.SI(net8707),
.CK(clk),
.Q(net8718),
.QN(net8717)
);

XOR2_X1 c8290(
.A(net7755),
.B(net8709),
.Z(net8719)
);

NOR2_X1 c8291(
.A1(net7740),
.A2(net8703),
.ZN(net8720)
);

AND4_X2 c8292(
.A1(net8696),
.A2(net8715),
.A3(net8701),
.A4(net8714),
.ZN(net8721)
);

AND4_X1 c8293(
.A1(net8690),
.A2(net8679),
.A3(net8645),
.A4(net8687),
.ZN(net8722)
);

OR2_X2 c8294(
.A1(net8722),
.A2(net8720),
.ZN(net8723)
);

AND3_X1 c8295(
.A1(net8662),
.A2(net8654),
.A3(net8714),
.ZN(net8724)
);

AOI22_X4 c8296(
.A1(net8724),
.A2(net8678),
.B1(net8707),
.ZN(net8725)
);

SDFF_X2 c8297(
.D(net8700),
.SE(net8699),
.SI(net8724),
.CK(clk),
.Q(net8727),
.QN(net8726)
);

OAI22_X4 c8298(
.A1(net8724),
.A2(net8706),
.B1(net8666),
.B2(net10411),
.ZN(net8728)
);

AOI222_X4 c8299(
.A1(net8724),
.A2(net8726),
.B1(net8670),
.B2(net8666),
.C1(net7730),
.C2(net10622),
.ZN(net8729)
);

NOR2_X4 c8300(
.A1(net7826),
.A2(net8689),
.ZN(net8730)
);

NOR2_X2 c8301(
.A1(net7736),
.A2(net6826),
.ZN(net8731)
);

XOR2_X2 c8302(
.A(net8714),
.B(net8664),
.Z(net8732)
);

INV_X32 c8303(
.A(net9678),
.ZN(net8733)
);

XNOR2_X1 c8304(
.A(net8719),
.B(net7854),
.ZN(net8734)
);

OR2_X4 c8305(
.A1(net8692),
.A2(net8714),
.ZN(net8735)
);

OR2_X1 c8306(
.A1(net8712),
.A2(net6843),
.ZN(net8736)
);

INV_X4 c8307(
.A(net3920),
.ZN(net8737)
);

XNOR2_X2 c8308(
.A(net7728),
.B(net5869),
.ZN(net8738)
);

AND2_X4 c8309(
.A1(net8707),
.A2(net8671),
.ZN(net8739)
);

AND2_X1 c8310(
.A1(net5810),
.A2(net8647),
.ZN(net8740)
);

INV_X1 c8311(
.A(net8652),
.ZN(net8741)
);

NAND2_X1 c8312(
.A1(net8736),
.A2(net6896),
.ZN(net8742)
);

INV_X2 c8313(
.A(net7777),
.ZN(net8743)
);

NAND2_X2 c8314(
.A1(net8713),
.A2(net6824),
.ZN(net8744)
);

INV_X8 c8315(
.A(net8664),
.ZN(net8745)
);

NAND2_X4 c8316(
.A1(net6755),
.A2(net3920),
.ZN(net8746)
);

AND2_X2 c8317(
.A1(net8710),
.A2(net11226),
.ZN(net8747)
);

INV_X16 c8318(
.A(net7878),
.ZN(net8748)
);

XOR2_X1 c8319(
.A(net7712),
.B(net8670),
.Z(net8749)
);

NOR2_X1 c8320(
.A1(net8723),
.A2(net6799),
.ZN(net8750)
);

OR2_X2 c8321(
.A1(net8727),
.A2(net11227),
.ZN(net8751)
);

NOR2_X4 c8322(
.A1(net8716),
.A2(net8731),
.ZN(net8752)
);

INV_X32 c8323(
.A(net8747),
.ZN(net8753)
);

NOR2_X2 c8324(
.A1(net8743),
.A2(net7776),
.ZN(net8754)
);

INV_X4 c8325(
.A(net8742),
.ZN(net8755)
);

NAND3_X1 c8326(
.A1(net8753),
.A2(net5822),
.A3(net8752),
.ZN(net8756)
);

XOR2_X2 c8327(
.A(net7854),
.B(net7736),
.Z(net8757)
);

INV_X1 c8328(
.A(net8680),
.ZN(net8758)
);

XNOR2_X1 c8329(
.A(net6827),
.B(net7801),
.ZN(net8759)
);

INV_X2 c8330(
.A(net8689),
.ZN(net8760)
);

INV_X8 c8331(
.A(net9677),
.ZN(net8761)
);

OR2_X4 c8332(
.A1(net8654),
.A2(net8738),
.ZN(net8762)
);

OR2_X1 c8333(
.A1(net8750),
.A2(net8673),
.ZN(net8763)
);

DFFRS_X1 c8334(
.D(net8701),
.RN(net8760),
.SN(net8714),
.CK(clk),
.Q(net8765),
.QN(net8764)
);

NOR3_X4 c8335(
.A1(net8748),
.A2(net6899),
.A3(net7854),
.ZN(net8766)
);

XNOR2_X2 c8336(
.A(net8755),
.B(net8760),
.ZN(net8767)
);

AND2_X4 c8337(
.A1(net7868),
.A2(net10517),
.ZN(net8768)
);

AND2_X1 c8338(
.A1(net8647),
.A2(net8684),
.ZN(net8769)
);

NOR3_X2 c8339(
.A1(net7752),
.A2(net8759),
.A3(net8741),
.ZN(net8770)
);

INV_X16 c8340(
.A(net9926),
.ZN(net8771)
);

NAND2_X1 c8341(
.A1(net8734),
.A2(net8761),
.ZN(net8772)
);

INV_X32 c8342(
.A(net8757),
.ZN(net8773)
);

DFFR_X1 c8343(
.D(net8772),
.RN(net8757),
.CK(clk),
.Q(net8775),
.QN(net8774)
);

NAND2_X2 c8344(
.A1(net8759),
.A2(net8751),
.ZN(net8776)
);

INV_X4 c8345(
.A(net8745),
.ZN(net8777)
);

AND3_X4 c8346(
.A1(net8697),
.A2(net8746),
.A3(net8664),
.ZN(net8778)
);

NAND2_X4 c8347(
.A1(net8671),
.A2(net8664),
.ZN(net8779)
);

AND2_X2 c8348(
.A1(net8776),
.A2(net8759),
.ZN(net8780)
);

INV_X1 c8349(
.A(net10333),
.ZN(net8781)
);

DFFR_X2 c8350(
.D(net8673),
.RN(net8701),
.CK(clk),
.Q(net8783),
.QN(net8782)
);

XOR2_X1 c8351(
.A(net8766),
.B(net8777),
.Z(net8784)
);

NOR2_X1 c8352(
.A1(net7717),
.A2(net8755),
.ZN(net8785)
);

NAND3_X2 c8353(
.A1(net8691),
.A2(net8757),
.A3(net8746),
.ZN(net8786)
);

OR2_X2 c8354(
.A1(net8775),
.A2(net8770),
.ZN(net8787)
);

OR3_X1 c8355(
.A1(net8653),
.A2(net8784),
.A3(net6843),
.ZN(net8788)
);

AOI221_X2 c8356(
.A(net8739),
.B1(net8761),
.B2(net8782),
.C1(net8760),
.C2(net8771),
.ZN(net8789)
);

MUX2_X1 c8357(
.A(net8693),
.B(net8773),
.S(net7807),
.Z(net8790)
);

OAI21_X4 c8358(
.A(net8767),
.B1(net8783),
.B2(net8784),
.ZN(net8791)
);

DFFRS_X2 c8359(
.D(net8786),
.RN(net8710),
.SN(net7712),
.CK(clk),
.Q(net8793),
.QN(net8792)
);

MUX2_X2 c8360(
.A(net8727),
.B(net8775),
.S(net8782),
.Z(net8794)
);

NOR2_X4 c8361(
.A1(net7855),
.A2(net8687),
.ZN(net8795)
);

NAND3_X4 c8362(
.A1(net8770),
.A2(net8793),
.A3(net8761),
.ZN(net8796)
);

OR3_X4 c8363(
.A1(net8795),
.A2(net8794),
.A3(net8792),
.ZN(net8797)
);

AND3_X2 c8364(
.A1(net6801),
.A2(net8796),
.A3(net7878),
.ZN(net8798)
);

NOR3_X1 c8365(
.A1(net6837),
.A2(net5935),
.A3(net8751),
.ZN(net8799)
);

NOR2_X2 c8366(
.A1(net8798),
.A2(net8793),
.ZN(net8800)
);

OR3_X2 c8367(
.A1(net8702),
.A2(net8784),
.A3(net8714),
.ZN(net8801)
);

OAI21_X2 c8368(
.A(net8800),
.B1(net8784),
.B2(net10807),
.ZN(net8802)
);

XOR2_X2 c8369(
.A(net8783),
.B(net8797),
.Z(net8803)
);

OAI21_X1 c8370(
.A(net5767),
.B1(net8708),
.B2(net8800),
.ZN(net8804)
);

XNOR2_X1 c8371(
.A(net8763),
.B(net8730),
.ZN(net8805)
);

AOI21_X2 c8372(
.A(net8803),
.B1(net8785),
.B2(net8697),
.ZN(net8806)
);

SDFF_X1 c8373(
.D(net8773),
.SE(net8805),
.SI(net10843),
.CK(clk),
.Q(net8808),
.QN(net8807)
);

AOI21_X1 c8374(
.A(net8806),
.B1(net8805),
.B2(net8779),
.ZN(net8809)
);

AOI21_X4 c8375(
.A(net8780),
.B1(net8801),
.B2(net7752),
.ZN(net8810)
);

SDFFRS_X2 c8376(
.D(net8799),
.RN(net7867),
.SE(net8797),
.SI(net7796),
.SN(net8649),
.CK(clk),
.Q(net8812),
.QN(net8811)
);

OR2_X4 c8377(
.A1(net8785),
.A2(net8774),
.ZN(net8813)
);

OAI33_X1 c8378(
.A1(net8752),
.A2(net8813),
.A3(net8812),
.B1(net8794),
.B2(net8771),
.B3(net7810),
.ZN(net8814)
);

AND3_X1 c8379(
.A1(net8778),
.A2(net4840),
.A3(net10639),
.ZN(net8815)
);

NAND3_X1 c8380(
.A1(net8800),
.A2(net7841),
.A3(net8808),
.ZN(net8816)
);

SDFFR_X2 c8381(
.D(net8735),
.RN(net8806),
.SE(net7796),
.SI(net10621),
.CK(clk),
.Q(net8818),
.QN(net8817)
);

AOI22_X2 c8382(
.A1(net8817),
.A2(net8811),
.B1(net10516),
.B2(net10600),
.ZN(net8819)
);

OR2_X1 c8383(
.A1(net6966),
.A2(net6899),
.ZN(net8820)
);

XNOR2_X2 c8384(
.A(net7801),
.B(net8684),
.ZN(net8821)
);

AND2_X4 c8385(
.A1(net6877),
.A2(net8797),
.ZN(net8822)
);

AND2_X1 c8386(
.A1(net8771),
.A2(net10585),
.ZN(net8823)
);

NOR3_X4 c8387(
.A1(net7840),
.A2(net8808),
.A3(net8670),
.ZN(net8824)
);

NAND2_X1 c8388(
.A1(net8821),
.A2(net7929),
.ZN(net8825)
);

INV_X2 c8389(
.A(net11051),
.ZN(net8826)
);

INV_X8 c8390(
.A(net8718),
.ZN(net8827)
);

INV_X16 c8391(
.A(net9999),
.ZN(net8828)
);

NAND2_X2 c8392(
.A1(net8735),
.A2(net7914),
.ZN(net8829)
);

NAND2_X4 c8393(
.A1(net8826),
.A2(net6975),
.ZN(net8830)
);

AND2_X2 c8394(
.A1(net7746),
.A2(net5035),
.ZN(net8831)
);

AOI221_X1 c8395(
.A(net8746),
.B1(net8805),
.B2(net7961),
.C1(net7918),
.C2(net8771),
.ZN(net8832)
);

XOR2_X1 c8396(
.A(net8737),
.B(net6020),
.Z(net8833)
);

NOR2_X1 c8397(
.A1(net8740),
.A2(net8812),
.ZN(net8834)
);

OR2_X2 c8398(
.A1(net7914),
.A2(net8827),
.ZN(net8835)
);

NOR2_X4 c8399(
.A1(net8779),
.A2(net8824),
.ZN(net8836)
);

NOR2_X2 c8400(
.A1(net8818),
.A2(net8831),
.ZN(net8837)
);

XOR2_X2 c8401(
.A(net6967),
.B(net8684),
.Z(net8838)
);

XNOR2_X1 c8402(
.A(net8761),
.B(net8670),
.ZN(net8839)
);

INV_X32 c8403(
.A(net10216),
.ZN(net8840)
);

OR2_X4 c8404(
.A1(net7704),
.A2(net8787),
.ZN(net8841)
);

SDFF_X2 c8405(
.D(net8839),
.SE(net7818),
.SI(net8746),
.CK(clk),
.Q(net8843),
.QN(net8842)
);

OR2_X1 c8406(
.A1(net6808),
.A2(net8840),
.ZN(net8844)
);

NOR3_X2 c8407(
.A1(net7868),
.A2(net8831),
.A3(net8835),
.ZN(net8845)
);

XNOR2_X2 c8408(
.A(net8797),
.B(net10474),
.ZN(net8846)
);

INV_X4 c8409(
.A(net10147),
.ZN(net8847)
);

INV_X1 c8410(
.A(net10159),
.ZN(net8848)
);

AND2_X4 c8411(
.A1(net5053),
.A2(net8846),
.ZN(net8849)
);

AND2_X1 c8412(
.A1(net6975),
.A2(net8761),
.ZN(net8850)
);

NAND2_X1 c8413(
.A1(net8655),
.A2(net8781),
.ZN(net8851)
);

AND3_X4 c8414(
.A1(net8733),
.A2(net7963),
.A3(net6824),
.ZN(net8852)
);

NAND2_X2 c8415(
.A1(net8781),
.A2(net8843),
.ZN(net8853)
);

NAND3_X2 c8416(
.A1(net8850),
.A2(net8717),
.A3(net7704),
.ZN(net8854)
);

OR3_X1 c8417(
.A1(net7835),
.A2(net7886),
.A3(net8853),
.ZN(net8855)
);

NAND2_X4 c8418(
.A1(net8687),
.A2(net8851),
.ZN(net8856)
);

AND2_X2 c8419(
.A1(net8807),
.A2(net10954),
.ZN(net8857)
);

INV_X2 c8420(
.A(net9998),
.ZN(net8858)
);

XOR2_X1 c8421(
.A(net8684),
.B(net8789),
.Z(net8859)
);

INV_X8 c8422(
.A(net9586),
.ZN(net8860)
);

NOR2_X1 c8423(
.A1(net6914),
.A2(net6933),
.ZN(net8861)
);

OAI221_X1 c8424(
.A(net8754),
.B1(net3920),
.B2(net8820),
.C1(net8811),
.C2(net10954),
.ZN(net8862)
);

SDFFS_X1 c8425(
.D(net7849),
.SE(net8833),
.SI(net8835),
.SN(net8831),
.CK(clk),
.Q(net8864),
.QN(net8863)
);

DFFRS_X1 c8426(
.D(net8857),
.RN(net8825),
.SN(net8861),
.CK(clk),
.Q(net8866),
.QN(net8865)
);

SDFFS_X2 c8427(
.D(net8791),
.SE(net8861),
.SI(net8794),
.SN(net8811),
.CK(clk),
.Q(net8868),
.QN(net8867)
);

OR2_X2 c8428(
.A1(net8835),
.A2(net7963),
.ZN(net8869)
);

OAI221_X4 c8429(
.A(net8790),
.B1(net8855),
.B2(net8819),
.C1(net7810),
.C2(net8760),
.ZN(net8870)
);

NOR2_X4 c8430(
.A1(net8833),
.A2(net11003),
.ZN(net8871)
);

NOR2_X2 c8431(
.A1(net8794),
.A2(net8867),
.ZN(net8872)
);

MUX2_X1 c8432(
.A(net6824),
.B(net8649),
.S(net8731),
.Z(net8873)
);

NAND4_X4 c8433(
.A1(net8708),
.A2(net7888),
.A3(net8825),
.A4(net8685),
.ZN(net8874)
);

OAI221_X2 c8434(
.A(net8847),
.B1(net8845),
.B2(net8863),
.C1(net6021),
.C2(net8651),
.ZN(net8875)
);

OAI21_X4 c8435(
.A(net8864),
.B1(net8831),
.B2(net8833),
.ZN(net8876)
);

DFFS_X1 c8436(
.D(net8670),
.SN(net7910),
.CK(clk),
.Q(net8878),
.QN(net8877)
);

XOR2_X2 c8437(
.A(net8705),
.B(net10893),
.Z(net8879)
);

XNOR2_X1 c8438(
.A(net8830),
.B(net8846),
.ZN(net8880)
);

INV_X16 c8439(
.A(net11051),
.ZN(net8881)
);

OR2_X4 c8440(
.A1(net8768),
.A2(net7961),
.ZN(net8882)
);

OR2_X1 c8441(
.A1(net8844),
.A2(net7888),
.ZN(net8883)
);

INV_X32 c8442(
.A(net10316),
.ZN(net8884)
);

XNOR2_X2 c8443(
.A(net8858),
.B(net8866),
.ZN(net8885)
);

AND2_X4 c8444(
.A1(net8885),
.A2(net5973),
.ZN(net8886)
);

AND2_X1 c8445(
.A1(net7888),
.A2(net8845),
.ZN(net8887)
);

NAND2_X1 c8446(
.A1(net8851),
.A2(net8797),
.ZN(net8888)
);

NAND2_X2 c8447(
.A1(net8888),
.A2(net10829),
.ZN(net8889)
);

NAND2_X4 c8448(
.A1(net8848),
.A2(net8808),
.ZN(net8890)
);

MUX2_X2 c8449(
.A(net8856),
.B(net8864),
.S(net8888),
.Z(net8891)
);

AND2_X2 c8450(
.A1(net8888),
.A2(net8818),
.ZN(net8892)
);

XOR2_X1 c8451(
.A(net7961),
.B(net11003),
.Z(net8893)
);

INV_X4 c8452(
.A(net9585),
.ZN(net8894)
);

NAND3_X4 c8453(
.A1(net8744),
.A2(net8868),
.A3(net8833),
.ZN(net8895)
);

OR3_X4 c8454(
.A1(net8894),
.A2(net8852),
.A3(net8885),
.ZN(net8896)
);

INV_X1 c8455(
.A(net10063),
.ZN(net8897)
);

NOR2_X1 c8456(
.A1(net8862),
.A2(net8885),
.ZN(net8898)
);

AND3_X2 c8457(
.A1(net6933),
.A2(net7835),
.A3(net11063),
.ZN(net8899)
);

OR2_X2 c8458(
.A1(net8879),
.A2(net8881),
.ZN(net8900)
);

NOR3_X1 c8459(
.A1(net6979),
.A2(net8863),
.A3(net10474),
.ZN(net8901)
);

NOR2_X4 c8460(
.A1(net8901),
.A2(net8892),
.ZN(net8902)
);

NOR2_X2 c8461(
.A1(net8769),
.A2(net6927),
.ZN(net8903)
);

OR3_X2 c8462(
.A1(net8887),
.A2(net8898),
.A3(net8865),
.ZN(net8904)
);

SDFFR_X1 c8463(
.D(net7963),
.RN(net8893),
.SE(net8769),
.SI(net8883),
.CK(clk),
.Q(net8906),
.QN(net8905)
);

SDFFRS_X1 c8464(
.D(net8902),
.RN(net8900),
.SE(net8903),
.SI(net8885),
.SN(net7724),
.CK(clk),
.Q(net8908),
.QN(net8907)
);

XOR2_X2 c8465(
.A(net8869),
.B(net8907),
.Z(net8909)
);

INV_X2 c8466(
.A(net11019),
.ZN(net8910)
);

XNOR2_X1 c8467(
.A(net6896),
.B(net8897),
.ZN(net8911)
);

INV_X8 c8468(
.A(net10957),
.ZN(net8912)
);

OR2_X4 c8469(
.A1(net6991),
.A2(net8003),
.ZN(net8913)
);

OAI21_X2 c8470(
.A(net7894),
.B1(net8658),
.B2(net7731),
.ZN(net8914)
);

OAI21_X1 c8471(
.A(net8022),
.B1(net8861),
.B2(net10956),
.ZN(net8915)
);

INV_X16 c8472(
.A(net11061),
.ZN(net8916)
);

OR2_X1 c8473(
.A1(net8915),
.A2(net11130),
.ZN(net8917)
);

INV_X32 c8474(
.A(net10240),
.ZN(net8918)
);

AOI21_X2 c8475(
.A(net8787),
.B1(net8884),
.B2(net8843),
.ZN(net8919)
);

XNOR2_X2 c8476(
.A(net7841),
.B(net7992),
.ZN(net8920)
);

AOI21_X1 c8477(
.A(net8047),
.B1(net8897),
.B2(net8831),
.ZN(net8921)
);

AND2_X4 c8478(
.A1(net7885),
.A2(net6991),
.ZN(net8922)
);

AND2_X1 c8479(
.A1(net7998),
.A2(net7982),
.ZN(net8923)
);

AOI21_X4 c8480(
.A(net4080),
.B1(net8923),
.B2(net8845),
.ZN(net8924)
);

NAND2_X1 c8481(
.A1(net5869),
.A2(net8751),
.ZN(net8925)
);

NAND2_X2 c8482(
.A1(net6091),
.A2(net8919),
.ZN(net8926)
);

AND3_X1 c8483(
.A1(net7072),
.A2(net6843),
.A3(net8651),
.ZN(net8927)
);

NAND2_X4 c8484(
.A1(net7814),
.A2(net11137),
.ZN(net8928)
);

AND2_X2 c8485(
.A1(net7071),
.A2(net7951),
.ZN(net8929)
);

NAND3_X1 c8486(
.A1(net7891),
.A2(net8649),
.A3(net10789),
.ZN(net8930)
);

DFFRS_X2 c8487(
.D(net7034),
.RN(net8845),
.SN(net8751),
.CK(clk),
.Q(net8932),
.QN(net8931)
);

DFFS_X2 c8488(
.D(net6021),
.SN(net8899),
.CK(clk),
.Q(net8934),
.QN(net8933)
);

NOR3_X4 c8489(
.A1(net8758),
.A2(net8738),
.A3(net7793),
.ZN(net8935)
);

NOR3_X2 c8490(
.A1(net7986),
.A2(net8846),
.A3(net8705),
.ZN(net8936)
);

XOR2_X1 c8491(
.A(net6951),
.B(net10901),
.Z(net8937)
);

SDFF_X1 c8492(
.D(net8914),
.SE(net8017),
.SI(net8819),
.CK(clk),
.Q(net8939),
.QN(net8938)
);

AND3_X4 c8493(
.A1(net8927),
.A2(net7918),
.A3(net7841),
.ZN(net8940)
);

NAND3_X2 c8494(
.A1(net8823),
.A2(net8928),
.A3(net8771),
.ZN(net8941)
);

NOR2_X1 c8495(
.A1(net8878),
.A2(net8905),
.ZN(net8942)
);

CLKGATETST_X1 c8496(
.E(net8017),
.SE(net8912),
.CK(clk),
.GCK(net8943)
);

SDFF_X2 c8497(
.D(net8788),
.SE(net8003),
.SI(net8927),
.CK(clk),
.Q(net8945),
.QN(net8944)
);

OR2_X2 c8498(
.A1(net7049),
.A2(net5869),
.ZN(net8946)
);

OR3_X1 c8499(
.A1(net7956),
.A2(net8877),
.A3(net8838),
.ZN(net8947)
);

NOR2_X4 c8500(
.A1(net7982),
.A2(net8658),
.ZN(net8948)
);

NOR2_X2 c8501(
.A1(net8940),
.A2(net7886),
.ZN(net8949)
);

INV_X4 c8502(
.A(net10241),
.ZN(net8950)
);

XOR2_X2 c8503(
.A(net8878),
.B(net10802),
.Z(net8951)
);

XNOR2_X1 c8504(
.A(net8951),
.B(net8908),
.ZN(net8952)
);

OR2_X4 c8505(
.A1(net8868),
.A2(net8903),
.ZN(net8953)
);

OR2_X1 c8506(
.A1(net8651),
.A2(net8866),
.ZN(net8954)
);

XNOR2_X2 c8507(
.A(net6951),
.B(net8949),
.ZN(net8955)
);

AND2_X4 c8508(
.A1(net8909),
.A2(net8915),
.ZN(net8956)
);

DFFRS_X1 c8509(
.D(net7731),
.RN(net8944),
.SN(net8926),
.CK(clk),
.Q(net8958),
.QN(net8957)
);

MUX2_X1 c8510(
.A(net8922),
.B(net6991),
.S(net8765),
.Z(net8959)
);

AND2_X1 c8511(
.A1(net8016),
.A2(net10867),
.ZN(net8960)
);

INV_X1 c8512(
.A(net10282),
.ZN(net8961)
);

CLKGATETST_X2 c8513(
.E(net8947),
.SE(net8658),
.CK(clk),
.GCK(net8962)
);

NAND2_X1 c8514(
.A1(net8958),
.A2(net8860),
.ZN(net8963)
);

OAI21_X4 c8515(
.A(net8920),
.B1(net8730),
.B2(net7049),
.ZN(net8964)
);

MUX2_X2 c8516(
.A(net8943),
.B(net8897),
.S(net8840),
.Z(net8965)
);

NAND2_X2 c8517(
.A1(net6933),
.A2(net8962),
.ZN(net8966)
);

NAND2_X4 c8518(
.A1(net8966),
.A2(net8840),
.ZN(net8967)
);

AND2_X2 c8519(
.A1(net8890),
.A2(net8758),
.ZN(net8968)
);

XOR2_X1 c8520(
.A(net8964),
.B(net8967),
.Z(net8969)
);

NOR2_X1 c8521(
.A1(net8965),
.A2(net8685),
.ZN(net8970)
);

NAND3_X4 c8522(
.A1(net7891),
.A2(net8022),
.A3(net8788),
.ZN(net8971)
);

OR3_X4 c8523(
.A1(net8917),
.A2(net8765),
.A3(net8915),
.ZN(net8972)
);

INV_X2 c8524(
.A(net10957),
.ZN(net8973)
);

OR2_X2 c8525(
.A1(net8831),
.A2(net10790),
.ZN(net8974)
);

OAI211_X2 c8526(
.A(net8966),
.B(net8943),
.C1(net8037),
.C2(net11097),
.ZN(net8975)
);

NOR2_X4 c8527(
.A1(net8963),
.A2(net6997),
.ZN(net8976)
);

NOR2_X2 c8528(
.A1(net8961),
.A2(net10777),
.ZN(net8977)
);

DFFRS_X2 c8529(
.D(net8977),
.RN(net8926),
.SN(net8973),
.CK(clk),
.Q(net8979),
.QN(net8978)
);

AND3_X2 c8530(
.A1(net8651),
.A2(net8914),
.A3(net10689),
.ZN(net8980)
);

NOR3_X1 c8531(
.A1(net7885),
.A2(net8963),
.A3(net11082),
.ZN(net8981)
);

OR3_X2 c8532(
.A1(net8949),
.A2(net8960),
.A3(net8975),
.ZN(net8982)
);

XOR2_X2 c8533(
.A(net8945),
.B(net8974),
.Z(net8983)
);

SDFF_X1 c8534(
.D(net8738),
.SE(net8957),
.SI(net8883),
.CK(clk),
.Q(net8985),
.QN(net8984)
);

SDFF_X2 c8535(
.D(net8730),
.SE(net8968),
.SI(net8985),
.CK(clk),
.Q(net8987),
.QN(net8986)
);

OAI21_X2 c8536(
.A(net8973),
.B1(net8958),
.B2(net8984),
.ZN(net8988)
);

OAI21_X1 c8537(
.A(net8925),
.B1(net8983),
.B2(net8985),
.ZN(net8989)
);

AOI21_X2 c8538(
.A(net7021),
.B1(net8985),
.B2(net7985),
.ZN(net8990)
);

AOI21_X1 c8539(
.A(net8974),
.B1(net10683),
.B2(net10714),
.ZN(net8991)
);

AOI21_X4 c8540(
.A(net8981),
.B1(net8966),
.B2(net8919),
.ZN(net8992)
);

AND3_X1 c8541(
.A1(net8845),
.A2(net8942),
.A3(net10956),
.ZN(net8993)
);

NAND3_X1 c8542(
.A1(net8976),
.A2(net8987),
.A3(net10751),
.ZN(net8994)
);

DFFRS_X1 c8543(
.D(net8993),
.RN(net10843),
.SN(net11136),
.CK(clk),
.Q(net8996),
.QN(net8995)
);

NOR3_X4 c8544(
.A1(net8935),
.A2(net8992),
.A3(net8995),
.ZN(net8997)
);

OR4_X2 c8545(
.A1(net8959),
.A2(net8970),
.A3(net8920),
.A4(net8811),
.ZN(net8998)
);

XNOR2_X1 c8546(
.A(net8010),
.B(net10581),
.ZN(net8999)
);

AOI221_X4 c8547(
.A(net8999),
.B1(net8994),
.B2(net8988),
.C1(net8984),
.C2(net7996),
.ZN(net9000)
);

NOR3_X2 c8548(
.A1(net8984),
.A2(net10473),
.A3(net10566),
.ZN(net9001)
);

AND3_X4 c8549(
.A1(net7951),
.A2(net8979),
.A3(net8938),
.ZN(net9002)
);

NAND3_X2 c8550(
.A1(net8135),
.A2(net8926),
.A3(net8975),
.ZN(net9003)
);

INV_X8 c8551(
.A(net11017),
.ZN(net9004)
);

OR2_X4 c8552(
.A1(net6843),
.A2(net8908),
.ZN(net9005)
);

OR2_X1 c8553(
.A1(net8053),
.A2(net8893),
.ZN(net9006)
);

XNOR2_X2 c8554(
.A(net8070),
.B(net8962),
.ZN(net9007)
);

OR3_X1 c8555(
.A1(net8828),
.A2(net9006),
.A3(net8986),
.ZN(net9008)
);

AND2_X4 c8556(
.A1(net8934),
.A2(net8859),
.ZN(net9009)
);

MUX2_X1 c8557(
.A(net8941),
.B(net8987),
.S(net8891),
.Z(net9010)
);

OAI21_X4 c8558(
.A(net7814),
.B1(net8889),
.B2(net9006),
.ZN(net9011)
);

AOI222_X2 c8559(
.A1(net8838),
.A2(net5166),
.B1(net9005),
.B2(net8926),
.C1(net8950),
.C2(net8978),
.ZN(net9012)
);

MUX2_X2 c8560(
.A(net7941),
.B(net8912),
.S(net8030),
.Z(net9013)
);

NAND3_X4 c8561(
.A1(net8893),
.A2(net9008),
.A3(net8954),
.ZN(net9014)
);

AND2_X1 c8562(
.A1(net8685),
.A2(net9014),
.ZN(net9015)
);

CLKGATETST_X4 c8563(
.E(net8784),
.SE(net8926),
.CK(clk),
.GCK(net9016)
);

OR3_X4 c8564(
.A1(net7793),
.A2(net9016),
.A3(net8865),
.ZN(net9017)
);

INV_X16 c8565(
.A(net10313),
.ZN(net9018)
);

AND3_X2 c8566(
.A1(net8929),
.A2(net7941),
.A3(net8126),
.ZN(net9019)
);

NAND2_X1 c8567(
.A1(net8950),
.A2(net8911),
.ZN(net9020)
);

NOR3_X1 c8568(
.A1(net8891),
.A2(net8685),
.A3(net8136),
.ZN(net9021)
);

INV_X32 c8569(
.A(net10371),
.ZN(net9022)
);

NAND2_X2 c8570(
.A1(net7964),
.A2(net8846),
.ZN(net9023)
);

OR3_X2 c8571(
.A1(net8952),
.A2(net8995),
.A3(net10828),
.ZN(net9024)
);

NAND2_X4 c8572(
.A1(net8954),
.A2(net8819),
.ZN(net9025)
);

AND2_X2 c8573(
.A1(net8882),
.A2(net8980),
.ZN(net9026)
);

OAI21_X2 c8574(
.A(net9023),
.B1(net8137),
.B2(net8037),
.ZN(net9027)
);

OAI21_X1 c8575(
.A(net8133),
.B1(net8784),
.B2(net11216),
.ZN(net9028)
);

AOI21_X2 c8576(
.A(net8137),
.B1(net8705),
.B2(net5934),
.ZN(net9029)
);

AOI21_X1 c8577(
.A(net6096),
.B1(net8992),
.B2(net7096),
.ZN(net9030)
);

XOR2_X1 c8578(
.A(net7992),
.B(net8016),
.Z(net9031)
);

AOI21_X4 c8579(
.A(net8906),
.B1(net9000),
.B2(net10794),
.ZN(net9032)
);

DFFRS_X2 c8580(
.D(net8866),
.RN(net9001),
.SN(net7088),
.CK(clk),
.Q(net9034),
.QN(net9033)
);

NOR2_X1 c8581(
.A1(net10801),
.A2(net11217),
.ZN(net9035)
);

AND3_X1 c8582(
.A1(net8056),
.A2(net9004),
.A3(net8921),
.ZN(net9036)
);

OAI222_X1 c8583(
.A1(net7985),
.A2(net8921),
.B1(net9005),
.B2(net9035),
.C1(net9019),
.C2(net8117),
.ZN(net9037)
);

NAND3_X1 c8584(
.A1(net8073),
.A2(net8649),
.A3(net8921),
.ZN(net9038)
);

OR2_X2 c8585(
.A1(net7966),
.A2(net8932),
.ZN(net9039)
);

NOR3_X4 c8586(
.A1(net8903),
.A2(net9029),
.A3(net8741),
.ZN(net9040)
);

NOR3_X2 c8587(
.A1(net8078),
.A2(net7796),
.A3(net8096),
.ZN(net9041)
);

AND3_X4 c8588(
.A1(net9025),
.A2(net9004),
.A3(net8126),
.ZN(net9042)
);

SDFF_X1 c8589(
.D(net9016),
.SE(net9014),
.SI(net8126),
.CK(clk),
.Q(net9044),
.QN(net9043)
);

SDFF_X2 c8590(
.D(net7810),
.SE(net9026),
.SI(net7088),
.CK(clk),
.Q(net9046),
.QN(net9045)
);

DFFRS_X1 c8591(
.D(net8968),
.RN(net9045),
.SN(net10750),
.CK(clk),
.Q(net9048),
.QN(net9047)
);

NAND3_X2 c8592(
.A1(net9041),
.A2(net9026),
.A3(net7964),
.ZN(net9049)
);

OR3_X1 c8593(
.A1(net7088),
.A2(net9027),
.A3(net8685),
.ZN(net9050)
);

MUX2_X1 c8594(
.A(net8916),
.B(net9029),
.S(net8014),
.Z(net9051)
);

OAI21_X4 c8595(
.A(net8853),
.B1(net9031),
.B2(net6096),
.ZN(net9052)
);

MUX2_X2 c8596(
.A(net8649),
.B(net8731),
.S(net9021),
.Z(net9053)
);

NAND3_X4 c8597(
.A1(net8837),
.A2(net8139),
.A3(net8913),
.ZN(net9054)
);

DFFRS_X2 c8598(
.D(net8906),
.RN(net9021),
.SN(net11207),
.CK(clk),
.Q(net9056),
.QN(net9055)
);

OR3_X4 c8599(
.A1(net9052),
.A2(net8852),
.A3(net9033),
.ZN(net9057)
);

AND3_X2 c8600(
.A1(net8126),
.A2(net9051),
.A3(net9033),
.ZN(net9058)
);

NOR3_X1 c8601(
.A1(net8030),
.A2(net8852),
.A3(net9047),
.ZN(net9059)
);

SDFF_X1 c8602(
.D(net8846),
.SE(net9010),
.SI(net8939),
.CK(clk),
.Q(net9061),
.QN(net9060)
);

OR3_X2 c8603(
.A1(net9013),
.A2(net9008),
.A3(net10900),
.ZN(net9062)
);

SDFF_X2 c8604(
.D(net9021),
.SE(net9031),
.SI(net8933),
.CK(clk),
.Q(net9064),
.QN(net9063)
);

INV_X4 c8605(
.A(net11017),
.ZN(net9065)
);

INV_X1 c8606(
.A(net10015),
.ZN(net9066)
);

OAI21_X2 c8607(
.A(net8819),
.B1(net9018),
.B2(net11207),
.ZN(net9067)
);

AOI221_X2 c8608(
.A(net8117),
.B1(net8070),
.B2(net9035),
.C1(net9043),
.C2(net8932),
.ZN(net9068)
);

OAI222_X4 c8609(
.A1(net8016),
.A2(net9061),
.B1(net9059),
.B2(net8975),
.C1(net8988),
.C2(net9019),
.ZN(net9069)
);

DFFRS_X1 c8610(
.D(net8956),
.RN(net7886),
.SN(net9059),
.CK(clk),
.Q(net9071),
.QN(net9070)
);

INV_X2 c8611(
.A(net9726),
.ZN(net9072)
);

OAI21_X1 c8612(
.A(net8658),
.B1(net8993),
.B2(net11052),
.ZN(net9073)
);

AOI21_X2 c8613(
.A(net9058),
.B1(net9062),
.B2(net9060),
.ZN(net9074)
);

DFFRS_X2 c8614(
.D(net8968),
.RN(net9071),
.SN(net8104),
.CK(clk),
.Q(net9076),
.QN(net9075)
);

OAI222_X2 c8615(
.A1(net9002),
.A2(net9076),
.B1(net9063),
.B2(net8986),
.C1(net9019),
.C2(net8111),
.ZN(net9077)
);

INV_X8 c8616(
.A(net9853),
.ZN(net9078)
);

AOI21_X1 c8617(
.A(net8910),
.B1(net8685),
.B2(net10699),
.ZN(net9079)
);

AOI21_X4 c8618(
.A(net9059),
.B1(net9078),
.B2(net9065),
.ZN(net9080)
);

AND3_X1 c8619(
.A1(net9066),
.A2(net8986),
.A3(net10714),
.ZN(net9081)
);

NAND3_X1 c8620(
.A1(net9021),
.A2(net9072),
.A3(net10414),
.ZN(net9082)
);

NOR3_X4 c8621(
.A1(net9061),
.A2(net8819),
.A3(net11018),
.ZN(net9083)
);

NOR3_X2 c8622(
.A1(net9079),
.A2(net8916),
.A3(net11096),
.ZN(net9084)
);

AND3_X4 c8623(
.A1(net9072),
.A2(net9078),
.A3(net10893),
.ZN(net9085)
);

SDFF_X1 c8624(
.D(net9028),
.SE(net9024),
.SI(net9070),
.CK(clk),
.Q(net9087),
.QN(net9086)
);

NAND3_X2 c8625(
.A1(net9001),
.A2(net9087),
.A3(net11018),
.ZN(net9088)
);

SDFF_X2 c8626(
.D(net9084),
.SE(net9051),
.SI(net9028),
.CK(clk),
.Q(net9090),
.QN(net9089)
);

OR3_X1 c8627(
.A1(net9088),
.A2(net9075),
.A3(net9067),
.ZN(net9091)
);

MUX2_X1 c8628(
.A(net9042),
.B(net8991),
.S(net10794),
.Z(net9092)
);

OAI21_X4 c8629(
.A(net9085),
.B1(net9019),
.B2(net10967),
.ZN(net9093)
);

CLKGATETST_X8 c8630(
.E(net8993),
.SE(net9091),
.CK(clk),
.GCK(net9094)
);

DFFRS_X1 c8631(
.D(net9011),
.RN(net9067),
.SN(net10415),
.CK(clk),
.Q(net9096),
.QN(net9095)
);

MUX2_X2 c8632(
.A(net9032),
.B(net8883),
.S(net8936),
.Z(net9097)
);

NOR2_X4 c8633(
.A1(net8057),
.A2(net8996),
.ZN(net9098)
);

NAND3_X4 c8634(
.A1(net9083),
.A2(net9032),
.A3(net8195),
.ZN(net9099)
);

INV_X16 c8635(
.A(net11110),
.ZN(net9100)
);

INV_X32 c8636(
.A(net11110),
.ZN(net9101)
);

NOR2_X2 c8637(
.A1(net9008),
.A2(net8820),
.ZN(net9102)
);

OR3_X4 c8638(
.A1(net9007),
.A2(net8861),
.A3(net8202),
.ZN(net9103)
);

AND3_X2 c8639(
.A1(net9089),
.A2(net9063),
.A3(net11077),
.ZN(net9104)
);

NOR3_X1 c8640(
.A1(net8097),
.A2(net8912),
.A3(net11110),
.ZN(net9105)
);

XOR2_X2 c8641(
.A(net8979),
.B(net7221),
.Z(net9106)
);

DFFRS_X2 c8642(
.D(net8105),
.RN(net9047),
.SN(net9098),
.CK(clk),
.Q(net9108),
.QN(net9107)
);

XNOR2_X1 c8643(
.A(net9096),
.B(net6768),
.ZN(net9109)
);

INV_X4 c8644(
.A(net10232),
.ZN(net9110)
);

OR2_X4 c8645(
.A1(net8913),
.A2(net9048),
.ZN(net9111)
);

OR2_X1 c8646(
.A1(net9006),
.A2(net9000),
.ZN(net9112)
);

XNOR2_X2 c8647(
.A(net7199),
.B(net9100),
.ZN(net9113)
);

SDFF_X1 c8648(
.D(net7096),
.SE(net8105),
.SI(net9112),
.CK(clk),
.Q(net9115),
.QN(net9114)
);

AND2_X4 c8649(
.A1(net8861),
.A2(net9104),
.ZN(net9116)
);

OR3_X2 c8650(
.A1(net9046),
.A2(net8812),
.A3(net7996),
.ZN(net9117)
);

AND2_X1 c8651(
.A1(net8202),
.A2(net7123),
.ZN(net9118)
);

NAND2_X1 c8652(
.A1(net8181),
.A2(net9103),
.ZN(net9119)
);

NAND2_X2 c8653(
.A1(net8097),
.A2(net7096),
.ZN(net9120)
);

NAND2_X4 c8654(
.A1(net8198),
.A2(net9087),
.ZN(net9121)
);

AND2_X2 c8655(
.A1(net8153),
.A2(net8213),
.ZN(net9122)
);

SDFFR_X2 c8656(
.D(net8195),
.RN(net9064),
.SE(net9107),
.SI(net8912),
.CK(clk),
.Q(net9124),
.QN(net9123)
);

XOR2_X1 c8657(
.A(net8160),
.B(net9123),
.Z(net9125)
);

OAI21_X2 c8658(
.A(net8980),
.B1(net9018),
.B2(net9125),
.ZN(net9126)
);

NOR2_X1 c8659(
.A1(net9124),
.A2(net9017),
.ZN(net9127)
);

OAI21_X1 c8660(
.A(net9065),
.B1(net9115),
.B2(net9095),
.ZN(net9128)
);

AOI21_X2 c8661(
.A(net8998),
.B1(net7996),
.B2(net10473),
.ZN(net9129)
);

AOI21_X1 c8662(
.A(net9120),
.B1(net7965),
.B2(net11098),
.ZN(net9130)
);

OR2_X2 c8663(
.A1(net9005),
.A2(net10918),
.ZN(net9131)
);

AOI21_X4 c8664(
.A(net8741),
.B1(net7965),
.B2(net9067),
.ZN(net9132)
);

AND3_X1 c8665(
.A1(net9118),
.A2(net8186),
.A3(net8153),
.ZN(net9133)
);

NAND3_X1 c8666(
.A1(net9117),
.A2(net9090),
.A3(net9035),
.ZN(net9134)
);

NOR3_X4 c8667(
.A1(net9102),
.A2(net9132),
.A3(net9098),
.ZN(net9135)
);

NOR3_X2 c8668(
.A1(net9128),
.A2(net9131),
.A3(net8096),
.ZN(net9136)
);

NOR2_X4 c8669(
.A1(net8003),
.A2(net8116),
.ZN(net9137)
);

AND3_X4 c8670(
.A1(net8751),
.A2(net8913),
.A3(net8918),
.ZN(net9138)
);

NAND3_X2 c8671(
.A1(net9125),
.A2(net9034),
.A3(net5315),
.ZN(net9139)
);

SDFF_X2 c8672(
.D(net9056),
.SE(net9132),
.SI(net7965),
.CK(clk),
.Q(net9141),
.QN(net9140)
);

OR3_X1 c8673(
.A1(net8939),
.A2(net9120),
.A3(net8152),
.ZN(net9142)
);

MUX2_X1 c8674(
.A(net7996),
.B(net8760),
.S(net9114),
.Z(net9143)
);

OAI21_X4 c8675(
.A(net9017),
.B1(net9105),
.B2(net9120),
.ZN(net9144)
);

MUX2_X2 c8676(
.A(net9137),
.B(net8105),
.S(net6273),
.Z(net9145)
);

NAND3_X4 c8677(
.A1(net8812),
.A2(net9121),
.A3(net8741),
.ZN(net9146)
);

AOI222_X1 c8678(
.A1(net9106),
.A2(net7965),
.B1(net8198),
.B2(net9120),
.C1(net9098),
.C2(net9086),
.ZN(net9147)
);

OR3_X4 c8679(
.A1(net9130),
.A2(net9142),
.A3(net8195),
.ZN(net9148)
);

NOR2_X2 c8680(
.A1(net8037),
.A2(net8181),
.ZN(net9149)
);

AND3_X2 c8681(
.A1(net7221),
.A2(net9144),
.A3(net9055),
.ZN(net9150)
);

NOR3_X1 c8682(
.A1(net9044),
.A2(net9146),
.A3(net9098),
.ZN(net9151)
);

DFFRS_X1 c8683(
.D(net9039),
.RN(net5315),
.SN(net9140),
.CK(clk),
.Q(net9153),
.QN(net9152)
);

XOR2_X2 c8684(
.A(net8912),
.B(net8884),
.Z(net9154)
);

OR3_X2 c8685(
.A1(net8116),
.A2(net9152),
.A3(net11110),
.ZN(net9155)
);

OAI21_X2 c8686(
.A(net9018),
.B1(net9007),
.B2(net10667),
.ZN(net9156)
);

OAI21_X1 c8687(
.A(net9155),
.B1(net9146),
.B2(net9137),
.ZN(net9157)
);

XNOR2_X1 c8688(
.A(net10867),
.B(net10918),
.ZN(net9158)
);

OR2_X4 c8689(
.A1(net7796),
.A2(net9143),
.ZN(net9159)
);

AOI21_X2 c8690(
.A(net8186),
.B1(net7243),
.B2(net8178),
.ZN(net9160)
);

AOI21_X1 c8691(
.A(net9159),
.B1(net9157),
.B2(net9142),
.ZN(net9161)
);

AOI21_X4 c8692(
.A(net6882),
.B1(net8898),
.B2(net9078),
.ZN(net9162)
);

AND3_X1 c8693(
.A1(net8218),
.A2(net9101),
.A3(net9019),
.ZN(net9163)
);

OR2_X1 c8694(
.A1(net9161),
.A2(net8918),
.ZN(net9164)
);

AOI211_X1 c8695(
.A(net9156),
.B(net9110),
.C1(out13),
.C2(net11077),
.ZN(net9165)
);

NAND3_X1 c8696(
.A1(net9109),
.A2(net9158),
.A3(net9140),
.ZN(net9166)
);

NOR3_X4 c8697(
.A1(net8884),
.A2(net9150),
.A3(net9159),
.ZN(net9167)
);

NOR3_X2 c8698(
.A1(net9138),
.A2(net9166),
.A3(net8186),
.ZN(net9168)
);

AND3_X4 c8699(
.A1(net9166),
.A2(net8860),
.A3(net8218),
.ZN(net9169)
);

NAND3_X2 c8700(
.A1(net8898),
.A2(net9169),
.A3(net9044),
.ZN(net9170)
);

OR3_X1 c8701(
.A1(net9168),
.A2(net9125),
.A3(net10842),
.ZN(net9171)
);

XNOR2_X2 c8702(
.A(net9156),
.B(net9143),
.ZN(net9172)
);

NAND4_X2 c8703(
.A1(net7243),
.A2(net9172),
.A3(net9166),
.A4(net9019),
.ZN(net9173)
);

MUX2_X1 c8704(
.A(net8991),
.B(net9157),
.S(net9112),
.Z(net9174)
);

OAI21_X4 c8705(
.A(net9146),
.B1(net9166),
.B2(net10667),
.ZN(net9175)
);

MUX2_X2 c8706(
.A(net9048),
.B(net8860),
.S(net8116),
.Z(net9176)
);

SDFFRS_X2 c8707(
.D(net9127),
.RN(net9167),
.SE(net9160),
.SI(net8998),
.SN(net8182),
.CK(clk),
.Q(net9178),
.QN(net9177)
);

NAND3_X4 c8708(
.A1(net8155),
.A2(net9158),
.A3(net9153),
.ZN(net9179)
);

OR4_X4 c8709(
.A1(net9154),
.A2(net9169),
.A3(net9177),
.A4(net10917),
.ZN(net9180)
);

OR3_X4 c8710(
.A1(net9022),
.A2(net9142),
.A3(net9172),
.ZN(net9181)
);

AND3_X2 c8711(
.A1(net9180),
.A2(net9176),
.A3(net10755),
.ZN(net9182)
);

OAI22_X2 c8712(
.A1(net9182),
.A2(net9172),
.B1(net9000),
.B2(net10842),
.ZN(net9183)
);

NOR3_X1 c8713(
.A1(net9150),
.A2(net9153),
.A3(net7996),
.ZN(net9184)
);

AOI222_X4 c8714(
.A1(net9165),
.A2(net9184),
.B1(net9183),
.B2(net9112),
.C1(net9086),
.C2(net9098),
.ZN(net9185)
);

AND2_X4 c8715(
.A1(net9122),
.A2(net10709),
.ZN(net9186)
);

OAI211_X4 c8716(
.A(net8240),
.B(net9035),
.C1(net8883),
.C2(net9120),
.ZN(net9187)
);

AND2_X1 c8717(
.A1(net8178),
.A2(net9186),
.ZN(net9188)
);

DFFRS_X2 c8718(
.D(net8987),
.RN(net9019),
.SN(net8731),
.CK(clk),
.Q(net9190),
.QN(net9189)
);

INV_X1 c8719(
.A(net11036),
.ZN(net9191)
);

OR3_X2 c8720(
.A1(net8946),
.A2(net7724),
.A3(net9019),
.ZN(net9192)
);

SDFF_X1 c8721(
.D(net8306),
.SE(net9183),
.SI(net8998),
.CK(clk),
.Q(net9194),
.QN(net9193)
);

NAND2_X1 c8722(
.A1(net8292),
.A2(net8820),
.ZN(net9195)
);

OAI21_X2 c8723(
.A(net9000),
.B1(net9094),
.B2(net10881),
.ZN(net9196)
);

INV_X2 c8724(
.A(net10160),
.ZN(net9197)
);

SDFF_X2 c8725(
.D(net8241),
.SE(net7199),
.SI(net9181),
.CK(clk),
.Q(net9199),
.QN(net9198)
);

NAND2_X2 c8726(
.A1(net9113),
.A2(net9110),
.ZN(net9200)
);

OAI21_X1 c8727(
.A(net9110),
.B1(net7822),
.B2(net10406),
.ZN(net9201)
);

NAND2_X4 c8728(
.A1(net8260),
.A2(net8312),
.ZN(net9202)
);

INV_X8 c8729(
.A(net9753),
.ZN(net9203)
);

AOI21_X2 c8730(
.A(net8230),
.B1(net8187),
.B2(net9203),
.ZN(net9204)
);

INV_X16 c8731(
.A(net9821),
.ZN(net9205)
);

AND2_X2 c8732(
.A1(net9186),
.A2(net8936),
.ZN(net9206)
);

XOR2_X1 c8733(
.A(net9134),
.B(net8260),
.Z(net9207)
);

AOI21_X1 c8734(
.A(net6282),
.B1(net9094),
.B2(net8771),
.ZN(net9208)
);

INV_X32 c8735(
.A(net9668),
.ZN(net9209)
);

NOR2_X1 c8736(
.A1(net6273),
.A2(net9116),
.ZN(net9210)
);

OAI33_X1 c8737(
.A1(net7317),
.A2(net8176),
.A3(net9172),
.B1(net8705),
.B2(net9120),
.B3(net9098),
.ZN(net9211)
);

AOI21_X4 c8738(
.A(net9191),
.B1(net3403),
.B2(net9186),
.ZN(net9212)
);

AND3_X1 c8739(
.A1(net9169),
.A2(net8240),
.A3(net11229),
.ZN(net9213)
);

NAND3_X1 c8740(
.A1(net9034),
.A2(net9197),
.A3(net9212),
.ZN(net9214)
);

OR2_X2 c8741(
.A1(net9188),
.A2(net9205),
.ZN(net9215)
);

NOR3_X4 c8742(
.A1(net7212),
.A2(net9122),
.A3(net9203),
.ZN(net9216)
);

NOR3_X2 c8743(
.A1(net9201),
.A2(net9035),
.A3(net8178),
.ZN(net9217)
);

AND3_X4 c8744(
.A1(net8121),
.A2(net7212),
.A3(net9160),
.ZN(net9218)
);

NAND3_X2 c8745(
.A1(net6356),
.A2(net9203),
.A3(net8827),
.ZN(net9219)
);

DFFRS_X1 c8746(
.D(net8731),
.RN(net8111),
.SN(net8121),
.CK(clk),
.Q(net9221),
.QN(net9220)
);

NOR2_X4 c8747(
.A1(net9181),
.A2(net8273),
.ZN(net9222)
);

DFFRS_X2 c8748(
.D(net9164),
.RN(net9216),
.SN(net6356),
.CK(clk),
.Q(net9224),
.QN(net9223)
);

OR3_X1 c8749(
.A1(net9160),
.A2(net8998),
.A3(net8312),
.ZN(net9225)
);

SDFF_X1 c8750(
.D(net3403),
.SE(net9209),
.SI(net8998),
.CK(clk),
.Q(net9227),
.QN(net9226)
);

MUX2_X1 c8751(
.A(net7087),
.B(net9087),
.S(net9205),
.Z(net9228)
);

OAI21_X4 c8752(
.A(net9216),
.B1(net9195),
.B2(net10737),
.ZN(net9229)
);

MUX2_X2 c8753(
.A(net9018),
.B(net9198),
.S(net9098),
.Z(net9230)
);

INV_X4 c8754(
.A(net9840),
.ZN(net9231)
);

NOR2_X2 c8755(
.A1(net9111),
.A2(net9207),
.ZN(net9232)
);

NAND3_X4 c8756(
.A1(net9221),
.A2(net9169),
.A3(net9197),
.ZN(net9233)
);

OR3_X4 c8757(
.A1(net8176),
.A2(net9190),
.A3(net9216),
.ZN(net9234)
);

SDFFS_X1 c8758(
.D(net9231),
.SE(net9232),
.SI(net7199),
.SN(net11230),
.CK(clk),
.Q(net9236),
.QN(net9235)
);

AND3_X2 c8759(
.A1(net9222),
.A2(net9085),
.A3(net10819),
.ZN(net9237)
);

INV_X1 c8760(
.A(net9667),
.ZN(net9238)
);

NOR3_X1 c8761(
.A1(net9209),
.A2(net9228),
.A3(net9215),
.ZN(net9239)
);

OAI211_X1 c8762(
.A(net9143),
.B(net9238),
.C1(net9220),
.C2(net7311),
.ZN(net9240)
);

SDFF_X2 c8763(
.D(net8187),
.SE(net8946),
.SI(net9234),
.CK(clk),
.Q(net9242),
.QN(net9241)
);

DFFRS_X1 c8764(
.D(net8911),
.RN(net9116),
.SN(net9019),
.CK(clk),
.Q(net9244),
.QN(net9243)
);

XOR2_X2 c8765(
.A(net9215),
.B(net8987),
.Z(net9245)
);

OR3_X2 c8766(
.A1(net9232),
.A2(net9239),
.A3(net7087),
.ZN(net9246)
);

OAI21_X2 c8767(
.A(net8996),
.B1(net9239),
.B2(net10755),
.ZN(net9247)
);

AOI221_X1 c8768(
.A(net9098),
.B1(net9236),
.B2(net9214),
.C1(net8883),
.C2(net8187),
.ZN(net9248)
);

OAI21_X1 c8769(
.A(net9000),
.B1(net9234),
.B2(net9236),
.ZN(net9249)
);

XNOR2_X1 c8770(
.A(net9241),
.B(net11090),
.ZN(net9250)
);

AOI21_X2 c8771(
.A(net9234),
.B1(net9226),
.B2(net7918),
.ZN(net9251)
);

OR2_X4 c8772(
.A1(net9212),
.A2(net10863),
.ZN(net9252)
);

NOR4_X4 c8773(
.A1(net7807),
.A2(net9227),
.A3(net8178),
.A4(net9235),
.ZN(net9253)
);

NOR4_X2 c8774(
.A1(net9141),
.A2(net9253),
.A3(net9235),
.A4(net10699),
.ZN(net9254)
);

OR2_X1 c8775(
.A1(net9168),
.A2(net8962),
.ZN(net9255)
);

DFFRS_X2 c8776(
.D(net9249),
.RN(net9254),
.SN(net9234),
.CK(clk),
.Q(net9257),
.QN(net9256)
);

XNOR2_X2 c8777(
.A(net9251),
.B(net9252),
.ZN(net9258)
);

AOI211_X4 c8778(
.A(net9250),
.B(net9242),
.C1(net4127),
.C2(net9252),
.ZN(net9259)
);

OAI221_X1 c8779(
.A(net9175),
.B1(net9108),
.B2(net9179),
.C1(net8014),
.C2(net9252),
.ZN(net9260)
);

AND2_X4 c8780(
.A1(net9085),
.A2(net8911),
.ZN(net9261)
);

OAI221_X4 c8781(
.A(net9233),
.B1(net9254),
.B2(net9205),
.C1(net9098),
.C2(net9235),
.ZN(net9262)
);

AOI21_X1 c8782(
.A(net9247),
.B1(net8998),
.B2(net9035),
.ZN(net9263)
);

AOI21_X4 c8783(
.A(net9242),
.B1(net9258),
.B2(net6927),
.ZN(net9264)
);

AND3_X1 c8784(
.A1(net9175),
.A2(net9236),
.A3(net10865),
.ZN(net9265)
);

NAND3_X1 c8785(
.A1(net8293),
.A2(net9259),
.A3(net6356),
.ZN(net9266)
);

NOR4_X1 c8786(
.A1(net9229),
.A2(net9265),
.A3(net9226),
.A4(net9235),
.ZN(net9267)
);

NOR3_X4 c8787(
.A1(net9227),
.A2(net9168),
.A3(net10862),
.ZN(net9268)
);

SDFF_X1 c8788(
.D(net9126),
.SE(net8827),
.SI(net9267),
.CK(clk),
.Q(net9270),
.QN(net9269)
);

AND2_X1 c8789(
.A1(net9213),
.A2(net9260),
.ZN(net9271)
);

SDFFRS_X1 c8790(
.D(net9271),
.RN(net9108),
.SE(net9238),
.SI(net9000),
.SN(net9098),
.CK(clk),
.Q(net9273),
.QN(net9272)
);

SDFF_X2 c8791(
.D(net9268),
.SE(net9254),
.SI(net10876),
.CK(clk),
.Q(net9275),
.QN(net9274)
);

NOR3_X2 c8792(
.A1(net9267),
.A2(net9265),
.A3(net10928),
.ZN(net9276)
);

AND3_X4 c8793(
.A1(net8936),
.A2(net9264),
.A3(net9265),
.ZN(net9277)
);

NAND3_X2 c8794(
.A1(net9258),
.A2(net9270),
.A3(net9252),
.ZN(net9278)
);

OR3_X1 c8795(
.A1(net9278),
.A2(net9269),
.A3(net10626),
.ZN(net9279)
);

DFFRS_X1 c8796(
.D(net9112),
.RN(net9274),
.SN(net10583),
.CK(clk),
.Q(net9281),
.QN(net9280)
);

DFFRS_X2 c8797(
.D(net9275),
.RN(net9268),
.SN(net10775),
.CK(clk),
.Q(net9283),
.QN(net9282)
);

NAND2_X1 c8798(
.A1(net8335),
.A2(net8376),
.ZN(net9284)
);

MUX2_X1 c8799(
.A(net9257),
.B(net9178),
.S(net6799),
.Z(net9285)
);

NAND2_X2 c8800(
.A1(net8996),
.A2(net11231),
.ZN(net9286)
);

NAND2_X4 c8801(
.A1(net4476),
.A2(net9081),
.ZN(net9287)
);

OAI21_X4 c8802(
.A(net9204),
.B1(net9236),
.B2(net10405),
.ZN(net9288)
);

INV_X2 c8803(
.A(net9977),
.ZN(net9289)
);

AND2_X2 c8804(
.A1(net9200),
.A2(net9240),
.ZN(net9290)
);

XOR2_X1 c8805(
.A(net9236),
.B(net11107),
.Z(net9291)
);

INV_X8 c8806(
.A(net9574),
.ZN(net9292)
);

OAI221_X2 c8807(
.A(net9287),
.B1(net8316),
.B2(net8376),
.C1(net9240),
.C2(net9086),
.ZN(net9293)
);

NOR2_X1 c8808(
.A1(net8182),
.A2(net8988),
.ZN(net9294)
);

MUX2_X2 c8809(
.A(net8142),
.B(net8771),
.S(net9256),
.Z(net9295)
);

NAND3_X4 c8810(
.A1(net9284),
.A2(net9081),
.A3(net9193),
.ZN(net9296)
);

OR3_X4 c8811(
.A1(net9288),
.A2(net8988),
.A3(net8278),
.ZN(net9297)
);

OR2_X2 c8812(
.A1(net5166),
.A2(net9285),
.ZN(net9298)
);

DFFR_X1 c8813(
.D(net8975),
.RN(net8370),
.CK(clk),
.Q(net9300),
.QN(net9299)
);

INV_X16 c8814(
.A(net11022),
.ZN(net9301)
);

AOI211_X2 c8815(
.A(net7347),
.B(net7421),
.C1(net8312),
.C2(net9296),
.ZN(net9302)
);

AOI22_X1 c8816(
.A1(net6226),
.A2(net8302),
.B1(net9223),
.B2(net8827),
.ZN(net9303)
);

SDFF_X1 c8817(
.D(net8111),
.SE(net6927),
.SI(net9296),
.CK(clk),
.Q(net9305),
.QN(net9304)
);

AND3_X2 c8818(
.A1(net7818),
.A2(net9178),
.A3(net9296),
.ZN(net9306)
);

NOR3_X1 c8819(
.A1(net8347),
.A2(out13),
.A3(net9252),
.ZN(net9307)
);

OR3_X2 c8820(
.A1(net9176),
.A2(net9094),
.A3(net9288),
.ZN(net9308)
);

OAI21_X2 c8821(
.A(net9307),
.B1(net9141),
.B2(net9218),
.ZN(net9309)
);

OAI21_X1 c8822(
.A(net9208),
.B1(net9272),
.B2(net11090),
.ZN(net9310)
);

AOI21_X2 c8823(
.A(net8370),
.B1(net9288),
.B2(net9214),
.ZN(net9311)
);

NOR2_X4 c8824(
.A1(net9303),
.A2(net9301),
.ZN(net9312)
);

AOI21_X1 c8825(
.A(net9195),
.B1(net7147),
.B2(net11225),
.ZN(net9313)
);

AOI21_X4 c8826(
.A(net9301),
.B1(net9064),
.B2(net9253),
.ZN(net9314)
);

AND3_X1 c8827(
.A1(net9217),
.A2(net9289),
.A3(net7421),
.ZN(net9315)
);

NOR2_X2 c8828(
.A1(net9081),
.A2(net9314),
.ZN(net9316)
);

XOR2_X2 c8829(
.A(net9312),
.B(net9309),
.Z(net9317)
);

XNOR2_X1 c8830(
.A(net9311),
.B(net9176),
.ZN(net9318)
);

SDFFRS_X2 c8831(
.D(net8921),
.RN(net9305),
.SE(net8988),
.SI(net8111),
.SN(net7357),
.CK(clk),
.Q(net9320),
.QN(net9319)
);

DFFR_X2 c8832(
.D(net9255),
.RN(net9294),
.CK(clk),
.Q(net9322),
.QN(net9321)
);

NAND3_X1 c8833(
.A1(net9252),
.A2(net7372),
.A3(net9063),
.ZN(net9323)
);

OR2_X4 c8834(
.A1(net9172),
.A2(net9311),
.ZN(net9324)
);

NOR3_X4 c8835(
.A1(net7421),
.A2(net10583),
.A3(net10752),
.ZN(net9325)
);

INV_X32 c8836(
.A(net9976),
.ZN(net9326)
);

SDFF_X2 c8837(
.D(net7395),
.SE(net9217),
.SI(net8921),
.CK(clk),
.Q(net9328),
.QN(net9327)
);

NOR3_X2 c8838(
.A1(net9322),
.A2(net9288),
.A3(net8369),
.ZN(net9329)
);

DFFS_X1 c8839(
.D(net7421),
.SN(net9318),
.CK(clk),
.Q(net9331),
.QN(net9330)
);

OR2_X1 c8840(
.A1(net8771),
.A2(net9316),
.ZN(net9332)
);

AND3_X4 c8841(
.A1(net8369),
.A2(net8883),
.A3(net8301),
.ZN(net9333)
);

NAND3_X2 c8842(
.A1(net9323),
.A2(net7311),
.A3(net11224),
.ZN(net9334)
);

XNOR2_X2 c8843(
.A(net8332),
.B(net9326),
.ZN(net9335)
);

INV_X4 c8844(
.A(net10044),
.ZN(net9336)
);

OR3_X1 c8845(
.A1(net7311),
.A2(out13),
.A3(net10923),
.ZN(net9337)
);

MUX2_X1 c8846(
.A(net9286),
.B(net9328),
.S(net10965),
.Z(net9338)
);

INV_X1 c8847(
.A(net9704),
.ZN(net9339)
);

OAI21_X4 c8848(
.A(net9199),
.B1(net9308),
.B2(net9319),
.ZN(net9340)
);

MUX2_X2 c8849(
.A(net8365),
.B(net9337),
.S(net9240),
.Z(net9341)
);

NAND3_X4 c8850(
.A1(net9290),
.A2(net7394),
.A3(net10549),
.ZN(net9342)
);

OR3_X4 c8851(
.A1(net8376),
.A2(net9304),
.A3(net9207),
.ZN(net9343)
);

AND3_X2 c8852(
.A1(net9218),
.A2(net9176),
.A3(net9319),
.ZN(net9344)
);

AND2_X4 c8853(
.A1(net9306),
.A2(net8988),
.ZN(net9345)
);

NOR3_X1 c8854(
.A1(net9334),
.A2(net7364),
.A3(net8771),
.ZN(net9346)
);

OR3_X2 c8855(
.A1(net9136),
.A2(net9214),
.A3(net9208),
.ZN(net9347)
);

OAI21_X2 c8856(
.A(net9311),
.B1(net8142),
.B2(net10384),
.ZN(net9348)
);

OAI21_X1 c8857(
.A(net9309),
.B1(net9327),
.B2(net10738),
.ZN(net9349)
);

AND2_X1 c8858(
.A1(net8312),
.A2(net9216),
.ZN(net9350)
);

AOI21_X2 c8859(
.A(net8014),
.B1(net9344),
.B2(net9285),
.ZN(net9351)
);

DFFRS_X1 c8860(
.D(net9339),
.RN(net9324),
.SN(net9308),
.CK(clk),
.Q(net9353),
.QN(net9352)
);

NAND2_X1 c8861(
.A1(net9332),
.A2(net9353),
.ZN(net9354)
);

AOI21_X1 c8862(
.A(net9345),
.B1(net9344),
.B2(net11231),
.ZN(net9355)
);

INV_X2 c8863(
.A(net9573),
.ZN(net9356)
);

AOI21_X4 c8864(
.A(net9338),
.B1(net9354),
.B2(net9299),
.ZN(net9357)
);

AND3_X1 c8865(
.A1(net9357),
.A2(net9354),
.A3(net9321),
.ZN(net9358)
);

NAND3_X1 c8866(
.A1(net9327),
.A2(net10548),
.A3(net10906),
.ZN(net9359)
);

AOI222_X2 c8867(
.A1(net9313),
.A2(net9309),
.B1(net9086),
.B2(net9340),
.C1(net8316),
.C2(net9352),
.ZN(net9360)
);

NOR3_X4 c8868(
.A1(net8322),
.A2(net9358),
.A3(net9356),
.ZN(net9361)
);

NOR3_X2 c8869(
.A1(net9361),
.A2(net9356),
.A3(net10820),
.ZN(net9362)
);

AND3_X4 c8870(
.A1(net9343),
.A2(net9337),
.A3(net8369),
.ZN(net9363)
);

NAND3_X2 c8871(
.A1(net8274),
.A2(net9326),
.A3(net9361),
.ZN(net9364)
);

NAND2_X2 c8872(
.A1(net9356),
.A2(net10953),
.ZN(net9365)
);

OR3_X1 c8873(
.A1(net7326),
.A2(net9291),
.A3(net9203),
.ZN(net9366)
);

NAND2_X4 c8874(
.A1(net9273),
.A2(net9203),
.ZN(net9367)
);

OAI222_X1 c8875(
.A1(net9366),
.A2(net9367),
.B1(net9078),
.B2(net9340),
.C1(net9361),
.C2(net11230),
.ZN(net9368)
);

MUX2_X1 c8876(
.A(net9330),
.B(net10735),
.S(net10885),
.Z(net9369)
);

OAI21_X4 c8877(
.A(net9369),
.B1(net9177),
.B2(net10965),
.ZN(net9370)
);

MUX2_X2 c8878(
.A(net9365),
.B(net10917),
.S(net11232),
.Z(net9371)
);

NAND3_X4 c8879(
.A1(net9370),
.A2(net9371),
.A3(net9120),
.ZN(net9372)
);

AOI221_X4 c8880(
.A(net9341),
.B1(net9334),
.B2(net9372),
.C1(net6391),
.C2(net11233),
.ZN(net9373)
);

AND2_X2 c8881(
.A1(net8705),
.A2(net9331),
.ZN(net9374)
);

OR3_X4 c8882(
.A1(net9356),
.A2(net9183),
.A3(net9336),
.ZN(net9375)
);

AND4_X4 c8883(
.A1(net8399),
.A2(net8231),
.A3(net8495),
.A4(net9020),
.ZN(net9376)
);

AND3_X2 c8884(
.A1(net9348),
.A2(net9208),
.A3(net9020),
.ZN(net9377)
);

AOI221_X2 c8885(
.A(net9194),
.B1(net9324),
.B2(net6391),
.C1(net9296),
.C2(net9356),
.ZN(net9378)
);

NOR3_X1 c8886(
.A1(net7372),
.A2(net7326),
.A3(net7431),
.ZN(net9379)
);

XOR2_X1 c8887(
.A(net9325),
.B(net11068),
.Z(net9380)
);

NOR2_X1 c8888(
.A1(net9342),
.A2(net7473),
.ZN(net9381)
);

DFFRS_X2 c8889(
.D(net9145),
.RN(net10625),
.SN(net10962),
.CK(clk),
.Q(net9383),
.QN(net9382)
);

OR2_X2 c8890(
.A1(net7123),
.A2(net9380),
.ZN(net9384)
);

OR3_X2 c8891(
.A1(net7147),
.A2(net9296),
.A3(net9206),
.ZN(net9385)
);

INV_X8 c8892(
.A(net9576),
.ZN(net9386)
);

SDFF_X1 c8893(
.D(net9245),
.SE(net9361),
.SI(net10871),
.CK(clk),
.Q(net9388),
.QN(net9387)
);

SDFF_X2 c8894(
.D(net8883),
.SE(net9240),
.SI(net11067),
.CK(clk),
.Q(net9390),
.QN(net9389)
);

OAI21_X2 c8895(
.A(net9224),
.B1(net9390),
.B2(net11089),
.ZN(net9391)
);

NOR2_X4 c8896(
.A1(net6388),
.A2(net9356),
.ZN(net9392)
);

OAI21_X1 c8897(
.A(net7357),
.B1(net9283),
.B2(net9177),
.ZN(net9393)
);

NOR2_X2 c8898(
.A1(net9380),
.A2(net11107),
.ZN(net9394)
);

AOI21_X2 c8899(
.A(net5530),
.B1(net9380),
.B2(net9240),
.ZN(net9395)
);

INV_X16 c8900(
.A(net9834),
.ZN(net9396)
);

XOR2_X2 c8901(
.A(net9376),
.B(net9380),
.Z(net9397)
);

AOI21_X1 c8902(
.A(net9208),
.B1(net8255),
.B2(net9396),
.ZN(net9398)
);

XNOR2_X1 c8903(
.A(net9020),
.B(net8319),
.ZN(net9399)
);

OR2_X4 c8904(
.A1(net7364),
.A2(net7372),
.ZN(net9400)
);

AOI21_X4 c8905(
.A(net7456),
.B1(net9386),
.B2(net9356),
.ZN(net9401)
);

INV_X32 c8906(
.A(net9575),
.ZN(net9402)
);

NAND4_X1 c8907(
.A1(net9401),
.A2(net9087),
.A3(net8412),
.A4(net9387),
.ZN(net9403)
);

AND3_X1 c8908(
.A1(net9320),
.A2(net9342),
.A3(net9193),
.ZN(net9404)
);

OR4_X1 c8909(
.A1(net9265),
.A2(net9383),
.A3(net8493),
.A4(net8827),
.ZN(net9405)
);

NAND3_X1 c8910(
.A1(net4534),
.A2(net8139),
.A3(net8412),
.ZN(net9406)
);

NOR3_X4 c8911(
.A1(net9336),
.A2(net9380),
.A3(net9382),
.ZN(net9407)
);

NOR3_X2 c8912(
.A1(net8412),
.A2(net9405),
.A3(net9401),
.ZN(net9408)
);

AND3_X4 c8913(
.A1(net9402),
.A2(net1708),
.A3(net10701),
.ZN(net9409)
);

OAI22_X1 c8914(
.A1(net5513),
.A2(net9300),
.B1(net8705),
.B2(net10878),
.ZN(net9410)
);

NAND3_X2 c8915(
.A1(net9328),
.A2(net9396),
.A3(net9020),
.ZN(net9411)
);

OR3_X1 c8916(
.A1(net9402),
.A2(net9078),
.A3(net9381),
.ZN(net9412)
);

MUX2_X1 c8917(
.A(net9194),
.B(net7357),
.S(net11067),
.Z(net9413)
);

OR2_X1 c8918(
.A1(net9411),
.A2(net10451),
.ZN(net9414)
);

OAI21_X4 c8919(
.A(net9396),
.B1(net7357),
.B2(net11119),
.ZN(net9415)
);

MUX2_X2 c8920(
.A(net9293),
.B(net9399),
.S(net8820),
.Z(net9416)
);

NAND3_X4 c8921(
.A1(net7519),
.A2(net9240),
.A3(net3565),
.ZN(net9417)
);

OR3_X4 c8922(
.A1(net9412),
.A2(net9413),
.A3(net9327),
.ZN(net9418)
);

AND3_X2 c8923(
.A1(net9417),
.A2(net9064),
.A3(net9253),
.ZN(net9419)
);

NOR3_X1 c8924(
.A1(net9331),
.A2(net8490),
.A3(net9388),
.ZN(net9420)
);

OR3_X2 c8925(
.A1(net9381),
.A2(net8420),
.A3(net11229),
.ZN(net9421)
);

OAI21_X2 c8926(
.A(net9078),
.B1(net9418),
.B2(net9243),
.ZN(net9422)
);

OAI21_X1 c8927(
.A(net8255),
.B1(net8412),
.B2(net10760),
.ZN(net9423)
);

AOI21_X2 c8928(
.A(net8439),
.B1(net7918),
.B2(net9410),
.ZN(net9424)
);

AOI21_X1 c8929(
.A(net7470),
.B1(net9372),
.B2(net9293),
.ZN(net9425)
);

SDFFS_X2 c8930(
.D(net9397),
.SE(net9394),
.SI(net9178),
.SN(net9425),
.CK(clk),
.Q(net9427),
.QN(net9426)
);

DFFRS_X1 c8931(
.D(net9404),
.RN(net9403),
.SN(net9410),
.CK(clk),
.Q(net9429),
.QN(net9428)
);

AOI21_X4 c8932(
.A(net9407),
.B1(net9423),
.B2(net9265),
.ZN(net9430)
);

AND3_X1 c8933(
.A1(net9424),
.A2(net9395),
.A3(net9340),
.ZN(net9431)
);

NAND3_X1 c8934(
.A1(net9359),
.A2(net9426),
.A3(net11119),
.ZN(net9432)
);

NOR3_X4 c8935(
.A1(net8319),
.A2(net9328),
.A3(net11026),
.ZN(net9433)
);

NOR3_X2 c8936(
.A1(net9325),
.A2(net9396),
.A3(net9265),
.ZN(net9434)
);

AND3_X4 c8937(
.A1(net7474),
.A2(net9429),
.A3(net9427),
.ZN(net9435)
);

XNOR2_X2 c8938(
.A(net8349),
.B(net9415),
.ZN(net9436)
);

NAND3_X2 c8939(
.A1(net9423),
.A2(net9392),
.A3(net9425),
.ZN(net9437)
);

AND2_X4 c8940(
.A1(net9400),
.A2(net9178),
.ZN(net9438)
);

OR3_X1 c8941(
.A1(net9416),
.A2(net9414),
.A3(net9342),
.ZN(net9439)
);

MUX2_X1 c8942(
.A(net9436),
.B(net9427),
.S(net9425),
.Z(net9440)
);

OAI21_X4 c8943(
.A(net6391),
.B1(net7456),
.B2(net9330),
.ZN(net9441)
);

MUX2_X2 c8944(
.A(net3565),
.B(net5513),
.S(net9418),
.Z(net9442)
);

NAND3_X4 c8945(
.A1(net9438),
.A2(net9420),
.A3(net8410),
.ZN(net9443)
);

OR3_X4 c8946(
.A1(net9419),
.A2(net7475),
.A3(net3575),
.ZN(net9444)
);

INV_X4 c8947(
.A(net9703),
.ZN(net9445)
);

AND3_X2 c8948(
.A1(net9435),
.A2(net9361),
.A3(net11068),
.ZN(net9446)
);

NOR3_X1 c8949(
.A1(net9141),
.A2(net9245),
.A3(net8421),
.ZN(net9447)
);

OR3_X2 c8950(
.A1(net9441),
.A2(net9409),
.A3(net9410),
.ZN(net9448)
);

OAI21_X2 c8951(
.A(net9418),
.B1(net9389),
.B2(net11091),
.ZN(net9449)
);

OAI21_X1 c8952(
.A(net9449),
.B1(net9381),
.B2(net10929),
.ZN(net9450)
);

OAI222_X4 c8953(
.A1(net9393),
.A2(net9442),
.B1(net9418),
.B2(net8420),
.C1(net7357),
.C2(net9292),
.ZN(net9451)
);

AOI21_X2 c8954(
.A(net9300),
.B1(net9422),
.B2(net9418),
.ZN(net9452)
);

AOI221_X1 c8955(
.A(net9421),
.B1(net8421),
.B2(net9425),
.C1(net7357),
.C2(net11235),
.ZN(net9453)
);

AOI21_X1 c8956(
.A(net9444),
.B1(net7357),
.B2(net10943),
.ZN(net9454)
);

AOI21_X4 c8957(
.A(net9432),
.B1(net9448),
.B2(net9320),
.ZN(net9455)
);

AND3_X1 c8958(
.A1(net8316),
.A2(net9447),
.A3(net11234),
.ZN(net9456)
);

NAND3_X1 c8959(
.A1(net9419),
.A2(net10966),
.A3(net11228),
.ZN(net9457)
);

OAI222_X2 c8960(
.A1(net9444),
.A2(net9436),
.B1(net9457),
.B2(net9410),
.C1(net9402),
.C2(net10947),
.ZN(net9458)
);

NOR3_X4 c8961(
.A1(net8435),
.A2(net9455),
.A3(net9428),
.ZN(net9459)
);

NOR3_X2 c8962(
.A1(net9434),
.A2(net9457),
.A3(net10742),
.ZN(net9460)
);

OAI221_X1 c8963(
.A(net9381),
.B1(net9457),
.B2(net9425),
.C1(net10934),
.C2(net11091),
.ZN(net9461)
);

AND3_X4 c8964(
.A1(net9361),
.A2(net7123),
.A3(net9389),
.ZN(net9462)
);

NAND3_X2 c8965(
.A1(net8231),
.A2(net8535),
.A3(net8827),
.ZN(net9463)
);

AND2_X1 c8966(
.A1(net7489),
.A2(net8225),
.ZN(net9464)
);

OR3_X1 c8967(
.A1(net7271),
.A2(net9390),
.A3(net9425),
.ZN(net9465)
);

NAND2_X1 c8968(
.A1(net9298),
.A2(net8501),
.ZN(net9466)
);

INV_X1 c8969(
.A(net9578),
.ZN(net9467)
);

MUX2_X1 c8970(
.A(net9464),
.B(net6477),
.S(net9410),
.Z(net9468)
);

DFFRS_X2 c8971(
.D(net8827),
.RN(net8535),
.SN(net10451),
.CK(clk),
.Q(net9470),
.QN(net9469)
);

OAI21_X4 c8972(
.A(net9280),
.B1(net9391),
.B2(net10761),
.ZN(net9471)
);

NAND2_X2 c8973(
.A1(net2737),
.A2(net10872),
.ZN(net9472)
);

MUX2_X2 c8974(
.A(net9244),
.B(net7431),
.S(net8225),
.Z(net9473)
);

NAND3_X4 c8975(
.A1(net9466),
.A2(net7561),
.A3(net9388),
.ZN(net9474)
);

NAND2_X4 c8976(
.A1(net8495),
.A2(net11225),
.ZN(net9475)
);

AND2_X2 c8977(
.A1(net8547),
.A2(net10878),
.ZN(net9476)
);

OR3_X4 c8978(
.A1(net9340),
.A2(net10866),
.A3(net11211),
.ZN(net9477)
);

AND3_X2 c8979(
.A1(net8419),
.A2(net9325),
.A3(net9340),
.ZN(net9478)
);

INV_X2 c8980(
.A(net9577),
.ZN(net9479)
);

NOR3_X1 c8981(
.A1(net8501),
.A2(net8587),
.A3(net9470),
.ZN(net9480)
);

OR3_X2 c8982(
.A1(net8341),
.A2(net9253),
.A3(net9425),
.ZN(net9481)
);

OAI21_X2 c8983(
.A(net9253),
.B1(net8182),
.B2(net9387),
.ZN(net9482)
);

OAI21_X1 c8984(
.A(net8568),
.B1(net9374),
.B2(net9335),
.ZN(net9483)
);

AOI21_X2 c8985(
.A(net8576),
.B1(net9394),
.B2(net10769),
.ZN(net9484)
);

XOR2_X1 c8986(
.A(net9340),
.B(net9484),
.Z(net9485)
);

AND4_X2 c8987(
.A1(net9203),
.A2(net9361),
.A3(net9374),
.A4(net8528),
.ZN(net9486)
);

NOR2_X1 c8988(
.A1(net8495),
.A2(net10968),
.ZN(net9487)
);

AOI21_X1 c8989(
.A(net7596),
.B1(net8583),
.B2(net10768),
.ZN(net9488)
);

AOI21_X4 c8990(
.A(net8516),
.B1(net9470),
.B2(net9479),
.ZN(net9489)
);

SDFF_X1 c8991(
.D(net3575),
.SE(net8535),
.SI(net9479),
.CK(clk),
.Q(net9491),
.QN(net9490)
);

AND3_X1 c8992(
.A1(net6414),
.A2(net9374),
.A3(net10935),
.ZN(net9492)
);

NAND3_X1 c8993(
.A1(net6554),
.A2(net9488),
.A3(net9490),
.ZN(net9493)
);

NOR3_X4 c8994(
.A1(net8820),
.A2(net9482),
.A3(net8529),
.ZN(net9494)
);

NOR3_X2 c8995(
.A1(net9474),
.A2(net9469),
.A3(net10990),
.ZN(net9495)
);

AND3_X4 c8996(
.A1(net9206),
.A2(net9340),
.A3(net11061),
.ZN(net9496)
);

AND4_X1 c8997(
.A1(net9425),
.A2(net8582),
.A3(net9469),
.A4(net7431),
.ZN(net9497)
);

NAND3_X2 c8998(
.A1(net8410),
.A2(net9475),
.A3(net8529),
.ZN(net9498)
);

OR3_X1 c8999(
.A1(net9372),
.A2(net8341),
.A3(net10523),
.ZN(net9499)
);

MUX2_X1 c9000(
.A(net9494),
.B(net9388),
.S(net9335),
.Z(net9500)
);

OAI21_X4 c9001(
.A(net9171),
.B1(net9476),
.B2(net9253),
.ZN(net9501)
);

MUX2_X2 c9002(
.A(net8494),
.B(net9394),
.S(out15),
.Z(net9502)
);

NAND3_X4 c9003(
.A1(net9296),
.A2(net9492),
.A3(net6477),
.ZN(net9503)
);

INV_X8 c9004(
.A(net9762),
.ZN(net9504)
);

INV_X16 c9005(
.A(net9763),
.ZN(net9505)
);

OR2_X2 c9006(
.A1(net9487),
.A2(net10668),
.ZN(net9506)
);

OR3_X4 c9007(
.A1(net9498),
.A2(net9471),
.A3(net8341),
.ZN(net9507)
);

AND3_X2 c9008(
.A1(net9491),
.A2(net9479),
.A3(net11089),
.ZN(net9508)
);

NOR3_X1 c9009(
.A1(net8331),
.A2(net9505),
.A3(net9507),
.ZN(net9509)
);

OR3_X2 c9010(
.A1(net9480),
.A2(net9509),
.A3(net9506),
.ZN(net9510)
);

OAI21_X2 c9011(
.A(net9374),
.B1(net9504),
.B2(net11008),
.ZN(net9511)
);

OAI21_X1 c9012(
.A(net9500),
.B1(net9511),
.B2(net10879),
.ZN(net9512)
);

AOI21_X2 c9013(
.A(net6593),
.B1(net8583),
.B2(net9388),
.ZN(net9513)
);

AOI21_X1 c9014(
.A(net8421),
.B1(net9281),
.B2(net9491),
.ZN(net9514)
);

AOI21_X4 c9015(
.A(net9491),
.B1(net10452),
.B2(net10990),
.ZN(net9515)
);

AOI222_X1 c9016(
.A1(net9489),
.A2(net9506),
.B1(net9504),
.B2(net9514),
.C1(net9490),
.C2(net9387),
.ZN(net9516)
);

AND3_X1 c9017(
.A1(net9467),
.A2(net9472),
.A3(net8410),
.ZN(net9517)
);

NAND3_X1 c9018(
.A1(net9477),
.A2(net9512),
.A3(net9502),
.ZN(net9518)
);

NOR3_X4 c9019(
.A1(net9308),
.A2(net9511),
.A3(net9498),
.ZN(net9519)
);

NOR3_X2 c9020(
.A1(net9514),
.A2(net9483),
.A3(net9506),
.ZN(net9520)
);

AOI222_X4 c9021(
.A1(net5551),
.A2(net9519),
.B1(net9506),
.B2(net9514),
.C1(net8182),
.C2(net9490),
.ZN(net9521)
);

AND3_X4 c9022(
.A1(net8513),
.A2(net9292),
.A3(net9502),
.ZN(net9522)
);

NAND3_X2 c9023(
.A1(net7584),
.A2(net9335),
.A3(net9514),
.ZN(net9523)
);

AOI22_X4 c9024(
.A1(net9516),
.A2(net9410),
.B1(net9512),
.B2(net9514),
.ZN(net9524)
);

OR3_X1 c9025(
.A1(net9315),
.A2(net9508),
.A3(net9514),
.ZN(net9525)
);

MUX2_X1 c9026(
.A(net7561),
.B(net9517),
.S(net9521),
.Z(net9526)
);

OAI21_X4 c9027(
.A(net9479),
.B1(net9518),
.B2(net9502),
.ZN(net9527)
);

MUX2_X2 c9028(
.A(net9523),
.B(net9493),
.S(net9499),
.Z(net9528)
);

NAND3_X4 c9029(
.A1(net9485),
.A2(net9527),
.A3(net9525),
.ZN(net9529)
);

OR3_X4 c9030(
.A1(net9510),
.A2(net9491),
.A3(net10546),
.ZN(net9530)
);

AND3_X2 c9031(
.A1(net9515),
.A2(net9525),
.A3(net11014),
.ZN(net9531)
);

OAI33_X1 c9032(
.A1(net9520),
.A2(net9445),
.A3(net9525),
.B1(net9387),
.B2(net8528),
.B3(net9514),
.ZN(net9532)
);

NOR3_X1 c9033(
.A1(net9391),
.A2(net9532),
.A3(net11014),
.ZN(net9533)
);

OR3_X2 c9034(
.A1(net9457),
.A2(net9525),
.A3(net9522),
.ZN(net9534)
);

OAI21_X2 c9035(
.A(net9524),
.B1(net9390),
.B2(net9533),
.ZN(net9535)
);

OAI21_X1 c9036(
.A(net9394),
.B1(net10523),
.B2(net11007),
.ZN(net9536)
);

AOI21_X2 c9037(
.A(net9526),
.B1(net9514),
.B2(net10844),
.ZN(net9537)
);

AOI21_X1 c9038(
.A(net9533),
.B1(net9537),
.B2(net9536),
.ZN(net9538)
);

OAI22_X4 c9039(
.A1(net8225),
.A2(net9531),
.B1(net10452),
.B2(net11016)
);

SDFFR_X1 merge9040(
.D(net5089),
.RN(net6120),
.SE(net6122),
.SI(net5953),
.CK(clk),
.Q(net9540),
.QN(net9539)
);

INV_X32 merge9041(
.A(net9950),
.ZN(net9541)
);

SDFF_X2 merge9042(
.D(net1783),
.SE(net1661),
.SI(net1759),
.CK(clk),
.Q(net9543),
.QN(net9542)
);

DFFRS_X1 merge9043(
.D(net4843),
.RN(net3850),
.SN(net3880),
.CK(clk),
.Q(net9545),
.QN(net9544)
);

DFFS_X2 merge9044(
.D(net876),
.SN(net852),
.CK(clk),
.Q(net9547),
.QN(net9546)
);

CLKGATETST_X1 merge9045(
.E(net414),
.SE(net147),
.CK(clk),
.GCK(net9548)
);

CLKGATETST_X2 merge9046(
.E(net6855),
.SE(net7778),
.CK(clk),
.GCK(net9549)
);

NOR2_X4 merge9047(
.A1(net1515),
.A2(net1522),
.ZN(net9550)
);

SDFFR_X2 merge9048(
.D(net2833),
.RN(net3369),
.SE(net3780),
.SI(net3769),
.CK(clk),
.Q(net9552),
.QN(net9551)
);

SDFFS_X1 merge9049(
.D(net7359),
.SE(net5315),
.SI(net7514),
.SN(net11210),
.CK(clk),
.Q(net9554),
.QN(net9553)
);

DFFRS_X2 merge9050(
.D(net2879),
.RN(net2885),
.SN(net1942),
.CK(clk),
.Q(net9556),
.QN(net9555)
);

CLKGATETST_X4 merge9051(
.E(net3198),
.SE(net3124),
.CK(clk),
.GCK(net9557)
);

INV_X4 merge9052(
.A(net9891),
.ZN(net9558)
);

AOI22_X2 merge9053(
.A1(net6534),
.A2(net8279),
.B1(net8443),
.B2(net8462),
.ZN(net9559)
);

CLKGATETST_X8 merge9054(
.E(net87),
.SE(net519),
.CK(clk),
.GCK(net9560)
);

SDFFS_X2 merge9055(
.D(net5315),
.SE(net6467),
.SI(net5604),
.SN(net5622),
.CK(clk),
.Q(net9562),
.QN(net9561)
);

NAND4_X4 merge9056(
.A1(net5454),
.A2(net5496),
.A3(net5539),
.A4(net5565),
.ZN(net9563)
);

INV_X1 merge9057(
.A(net9792),
.ZN(net9564)
);

INV_X2 merge9058(
.A(net10253),
.ZN(net9565)
);

INV_X8 merge9059(
.A(net10903),
.ZN(net9566)
);

DFFR_X1 merge9060(
.D(net1078),
.RN(net1051),
.CK(clk),
.Q(net9568),
.QN(net9567)
);

SDFFR_X1 merge9061(
.D(net8055),
.RN(net8060),
.SE(net8076),
.SI(net8119),
.CK(clk),
.Q(net9570),
.QN(net9569)
);

DFFR_X2 merge9062(
.D(net1920),
.RN(net2960),
.CK(clk),
.Q(net9572),
.QN(net9571)
);

SDFFR_X2 merge9063(
.D(net9207),
.RN(net9119),
.SE(net9344),
.SI(net10663),
.CK(clk),
.Q(net9574),
.QN(net9573)
);

SDFFS_X1 merge9064(
.D(net7509),
.SE(net9381),
.SI(net9282),
.SN(net9384),
.CK(clk),
.Q(net9576),
.QN(net9575)
);

SDFFS_X2 merge9065(
.D(net8528),
.SE(net9425),
.SI(net9478),
.SN(net9145),
.CK(clk),
.Q(net9578),
.QN(net9577)
);

NOR2_X2 merge9066(
.A1(net8317),
.A2(net7724),
.ZN(net9579)
);

SDFFR_X1 merge9067(
.D(net8216),
.RN(net8164),
.SE(net8242),
.SI(net8306),
.CK(clk),
.Q(net9581),
.QN(net9580)
);

INV_X16 merge9068(
.A(net10008),
.ZN(net9582)
);

DFFS_X1 merge9069(
.D(net6807),
.SN(net4961),
.CK(clk),
.Q(net9584),
.QN(net9583)
);

SDFFR_X2 merge9070(
.D(net8807),
.RN(net8855),
.SE(net8875),
.SI(net8789),
.CK(clk),
.Q(net9586),
.QN(net9585)
);

AOI21_X4 merge9071(
.A(net3141),
.B1(net2943),
.B2(net3119),
.ZN(net9587)
);

INV_X32 merge9072(
.A(net10161),
.ZN(net9588)
);

AND3_X1 merge9073(
.A1(net552),
.A2(net1525),
.A3(net2209),
.ZN(net9589)
);

NAND3_X1 merge9074(
.A1(net4443),
.A2(net4437),
.A3(net10567),
.ZN(net9590)
);

INV_X4 merge9075(
.A(net9982),
.ZN(net9591)
);

DFFS_X2 merge9076(
.D(net208),
.SN(net186),
.CK(clk),
.Q(net9593),
.QN(net9592)
);

INV_X1 merge9077(
.A(net9908),
.ZN(net9594)
);

XOR2_X2 merge9078(
.A(net3454),
.B(net3562),
.Z(net9595)
);

NOR3_X4 merge9079(
.A1(net3303),
.A2(net4150),
.A3(net10680),
.ZN(net9596)
);

CLKGATETST_X1 merge9080(
.E(net843),
.SE(net760),
.CK(clk),
.GCK(net9597)
);

OAI211_X2 merge9081(
.A(net8931),
.B(net8921),
.C1(net7922),
.C2(net9049),
.ZN(net9598)
);

SDFFRS_X1 merge9082(
.D(net6683),
.RN(net6700),
.SE(net7181),
.SI(net7654),
.SN(net6452),
.CK(clk),
.Q(net9600),
.QN(net9599)
);

SDFFS_X1 merge9083(
.D(net3784),
.SE(net2808),
.SI(net3764),
.SN(net1844),
.CK(clk),
.Q(net9602),
.QN(net9601)
);

OR4_X2 merge9084(
.A1(net8886),
.A2(net8891),
.A3(net8825),
.A4(net8730),
.ZN(net9603)
);

INV_X2 merge9085(
.A(net9862),
.ZN(net9604)
);

INV_X8 merge9086(
.A(net10998),
.ZN(net9605)
);

SDFF_X1 merge9087(
.D(net6726),
.SE(net4341),
.SI(net6283),
.CK(clk),
.Q(net9607),
.QN(net9606)
);

CLKGATETST_X2 merge9088(
.E(net1011),
.SE(net1103),
.CK(clk),
.GCK(net9608)
);

INV_X16 merge9089(
.A(net9885),
.ZN(net9609)
);

XNOR2_X1 merge9090(
.A(net213),
.B(net1124),
.ZN(net9610)
);

CLKGATETST_X4 merge9091(
.E(net3322),
.SE(net4299),
.CK(clk),
.GCK(net9611)
);

INV_X32 merge9092(
.A(net11123),
.ZN(net9612)
);

OR2_X4 merge9093(
.A1(net1288),
.A2(net1435),
.ZN(net9613)
);

AOI222_X2 merge9094(
.A1(net8573),
.A2(net8523),
.B1(net8633),
.B2(net7553),
.C1(net8619),
.C2(net6650),
.ZN(net9614)
);

SDFFS_X2 merge9095(
.D(net8502),
.SE(net5474),
.SI(net8526),
.SN(net11062),
.CK(clk),
.Q(net9616),
.QN(net9615)
);

AOI211_X1 merge9096(
.A(net4457),
.B(net4672),
.C1(net4673),
.C2(net11099),
.ZN(net9617)
);

CLKGATETST_X8 merge9097(
.E(net3918),
.SE(net3930),
.CK(clk),
.GCK(net9618)
);

INV_X4 merge9098(
.A(net9693),
.ZN(net9619)
);

DFFR_X1 merge9099(
.D(net1374),
.RN(net458),
.CK(clk),
.Q(net9621),
.QN(net9620)
);

INV_X1 merge9100(
.A(net10226),
.ZN(net9622)
);

OR2_X1 merge9101(
.A1(net506),
.A2(net668),
.ZN(net9623)
);

DFFR_X2 merge9102(
.D(net5824),
.RN(net5838),
.CK(clk),
.Q(net9625),
.QN(net9624)
);

DFFS_X1 merge9103(
.D(net7707),
.SN(net7726),
.CK(clk),
.Q(net9627),
.QN(net9626)
);

INV_X2 merge9104(
.A(net10850),
.ZN(net9628)
);

INV_X8 merge9105(
.A(net10049),
.ZN(net9629)
);

INV_X16 merge9106(
.A(net10072),
.ZN(net9630)
);

SDFF_X2 merge9107(
.D(net8119),
.SE(net6027),
.SI(net8206),
.CK(clk),
.Q(net9632),
.QN(net9631)
);

INV_X32 merge9108(
.A(net9989),
.ZN(net9633)
);

NAND4_X2 merge9109(
.A1(net5512),
.A2(net4691),
.A3(net5666),
.A4(net5664),
.ZN(net9634)
);

INV_X4 merge9110(
.A(net10268),
.ZN(net9635)
);

XNOR2_X2 merge9111(
.A(net213),
.B(net347),
.ZN(net9636)
);

DFFRS_X1 merge9112(
.D(net6284),
.RN(net6197),
.SN(net6395),
.CK(clk),
.Q(net9638),
.QN(net9637)
);

DFFRS_X2 merge9113(
.D(net3377),
.RN(net3364),
.SN(net11048),
.CK(clk),
.Q(net9640),
.QN(net9639)
);

OR4_X4 merge9114(
.A1(net7015),
.A2(net7708),
.A3(net8027),
.A4(net8039),
.ZN(net9641)
);

INV_X1 merge9115(
.A(net10065),
.ZN(net9642)
);

SDFFR_X1 merge9116(
.D(net1745),
.RN(net1856),
.SE(net1880),
.SI(net2825),
.CK(clk),
.Q(net9644),
.QN(net9643)
);

DFFS_X2 merge9117(
.D(net5764),
.SN(net5864),
.CK(clk),
.Q(net9646),
.QN(net9645)
);

SDFFR_X2 merge9118(
.D(net3794),
.RN(net5672),
.SE(net5717),
.SI(net5586),
.CK(clk),
.Q(net9648),
.QN(net9647)
);

CLKGATETST_X1 merge9119(
.E(net2946),
.SE(net1920),
.CK(clk),
.GCK(net9649)
);

SDFFS_X1 merge9120(
.D(net4007),
.SE(net5103),
.SI(net5101),
.SN(net5059),
.CK(clk),
.Q(net9651),
.QN(net9650)
);

OAI22_X2 merge9121(
.A1(net1638),
.A2(net1505),
.B1(net1643),
.B2(net1647),
.ZN(net9652)
);

SDFF_X1 merge9122(
.D(net6558),
.SE(net5580),
.SI(net3723),
.CK(clk),
.Q(net9654),
.QN(net9653)
);

AND2_X4 merge9123(
.A1(net1934),
.A2(net1023),
.ZN(net9655)
);

INV_X2 merge9124(
.A(net10190),
.ZN(net9656)
);

INV_X8 merge9125(
.A(net9931),
.ZN(net9657)
);

INV_X16 merge9126(
.A(net9695),
.ZN(net9658)
);

CLKGATETST_X2 merge9127(
.E(net483),
.SE(net484),
.CK(clk),
.GCK(net9659)
);

CLKGATETST_X4 merge9128(
.E(net7716),
.SE(net6786),
.CK(clk),
.GCK(net9660)
);

INV_X32 merge9129(
.A(net10252),
.ZN(net9661)
);

OAI211_X4 merge9130(
.A(net8147),
.B(net9085),
.C1(net8992),
.C2(net7918),
.ZN(net9662)
);

INV_X4 merge9131(
.A(net10111),
.ZN(net9663)
);

INV_X1 merge9132(
.A(net10064),
.ZN(net9664)
);

SDFFS_X2 merge9133(
.D(net7251),
.SE(net7257),
.SI(net6372),
.SN(net7047),
.CK(clk),
.Q(net9666),
.QN(net9665)
);

SDFFR_X1 merge9134(
.D(net8278),
.RN(net9160),
.SE(net9210),
.SI(net8292),
.CK(clk),
.Q(net9668),
.QN(net9667)
);

NOR3_X2 merge9135(
.A1(net4070),
.A2(net4167),
.A3(net4005),
.ZN(net9669)
);

INV_X2 merge9136(
.A(net9696),
.ZN(net9670)
);

OAI211_X1 merge9137(
.A(net482),
.B(net4305),
.C1(net4410),
.C2(net3469),
.ZN(net9671)
);

AND3_X4 merge9138(
.A1(net5899),
.A2(net6038),
.A3(net6991),
.ZN(net9672)
);

CLKGATETST_X8 merge9139(
.E(net5763),
.SE(net5781),
.CK(clk),
.GCK(net9673)
);

INV_X8 merge9140(
.A(net10057),
.ZN(net9674)
);

DFFR_X1 merge9141(
.D(net5976),
.RN(net6026),
.CK(clk),
.Q(net9676),
.QN(net9675)
);

SDFF_X2 merge9142(
.D(net5808),
.SE(net8732),
.SI(net8735),
.CK(clk),
.Q(net9678),
.QN(net9677)
);

DFFR_X2 merge9143(
.D(net6149),
.RN(net5296),
.CK(clk),
.Q(net9680),
.QN(net9679)
);

INV_X16 merge9144(
.A(net9802),
.ZN(net9681)
);

DFFS_X1 merge9145(
.D(net1010),
.SN(net1007),
.CK(clk),
.Q(net9683),
.QN(net9682)
);

INV_X32 merge9146(
.A(net10835),
.ZN(net9684)
);

SDFFR_X2 merge9147(
.D(net3758),
.RN(net3825),
.SE(net5748),
.SI(net5692),
.CK(clk),
.Q(net9686),
.QN(net9685)
);

INV_X4 merge9148(
.A(net10188),
.ZN(net9687)
);

SDFFS_X1 merge9149(
.D(net5264),
.SE(net4691),
.SI(net1615),
.SN(net3685),
.CK(clk),
.Q(net9689),
.QN(net9688)
);

INV_X1 merge9150(
.A(net10114),
.ZN(net9690)
);

SDFFS_X2 merge9151(
.D(net8423),
.SE(net8111),
.SI(net6563),
.SN(net4600),
.CK(clk),
.Q(net9692),
.QN(net9691)
);

INV_X2 merge9152(
.A(net10528),
.ZN(net9693)
);

NOR4_X4 merge9153(
.A1(net6526),
.A2(net6550),
.A3(net2809),
.A4(net5704),
.ZN(net9694)
);

DFFRS_X1 merge9154(
.D(net41),
.RN(net37),
.SN(net106),
.CK(clk),
.Q(net9696),
.QN(net9695)
);

DFFS_X2 merge9155(
.D(net228),
.SN(net1092),
.CK(clk),
.Q(net9698),
.QN(net9697)
);

INV_X8 merge9156(
.A(net10031),
.ZN(net9699)
);

INV_X16 merge9157(
.A(net10235),
.ZN(net9700)
);

CLKGATETST_X1 merge9158(
.E(net5775),
.SE(net5781),
.CK(clk),
.GCK(net9701)
);

INV_X32 merge9159(
.A(net11116),
.ZN(net9702)
);

SDFFR_X1 merge9160(
.D(net4449),
.RN(net8975),
.SE(net9442),
.SI(net9433),
.CK(clk),
.Q(net9704),
.QN(net9703)
);

NOR4_X2 merge9161(
.A1(net8334),
.A2(net4524),
.A3(net7601),
.A4(net7586),
.ZN(net9705)
);

CLKGATETST_X2 merge9162(
.E(net6767),
.SE(net6904),
.CK(clk),
.GCK(net9706)
);

CLKGATETST_X4 merge9163(
.E(net4303),
.SE(net5261),
.CK(clk),
.GCK(net9707)
);

AND2_X1 merge9164(
.A1(net1174),
.A2(net335),
.ZN(net9708)
);

INV_X4 merge9165(
.A(net9901),
.ZN(net9709)
);

CLKGATETST_X8 merge9166(
.E(net6738),
.SE(net6783),
.CK(clk),
.GCK(net9710)
);

INV_X1 merge9167(
.A(net9991),
.ZN(net9711)
);

INV_X2 merge9168(
.A(net10176),
.ZN(net9712)
);

SDFFR_X2 merge9169(
.D(net2732),
.RN(net5307),
.SE(net6543),
.SI(net6547),
.CK(clk),
.Q(net9714),
.QN(net9713)
);

SDFFS_X1 merge9170(
.D(net6575),
.SE(net7407),
.SI(net8496),
.SN(net8519),
.CK(clk),
.Q(net9716),
.QN(net9715)
);

DFFR_X1 merge9171(
.D(net7710),
.RN(net5019),
.CK(clk),
.Q(net9718),
.QN(net9717)
);

DFFR_X2 merge9172(
.D(net8649),
.RN(net5766),
.CK(clk),
.Q(net9720),
.QN(net9719)
);

DFFS_X1 merge9173(
.D(net3969),
.SN(net4103),
.CK(clk),
.Q(net9722),
.QN(net9721)
);

INV_X8 merge9174(
.A(net10019),
.ZN(net9723)
);

NAND2_X1 merge9175(
.A1(net186),
.A2(net277),
.ZN(net9724)
);

INV_X16 merge9176(
.A(net11125),
.ZN(net9725)
);

SDFFS_X2 merge9177(
.D(net8200),
.SE(net7224),
.SI(net9062),
.SN(net8853),
.CK(clk),
.Q(net9727),
.QN(net9726)
);

INV_X32 merge9178(
.A(net11120),
.ZN(net9728)
);

INV_X4 merge9179(
.A(net11101),
.ZN(net9729)
);

INV_X1 merge9180(
.A(net10286),
.ZN(net9730)
);

DFFS_X2 merge9181(
.D(net6750),
.SN(net6765),
.CK(clk),
.Q(net9732),
.QN(net9731)
);

INV_X2 merge9182(
.A(net10073),
.ZN(net9733)
);

CLKGATETST_X1 merge9183(
.E(net519),
.SE(net632),
.CK(clk),
.GCK(net9734)
);

INV_X8 merge9184(
.A(net10121),
.ZN(net9735)
);

CLKGATETST_X2 merge9185(
.E(net3396),
.SE(net4437),
.CK(clk),
.GCK(net9736)
);

INV_X16 merge9186(
.A(net10265),
.ZN(net9737)
);

CLKGATETST_X4 merge9187(
.E(net1944),
.SE(net160),
.CK(clk),
.GCK(net9738)
);

CLKGATETST_X8 merge9188(
.E(net5871),
.SE(net5807),
.CK(clk),
.GCK(net9739)
);

NAND2_X2 merge9189(
.A1(net252),
.A2(net211),
.ZN(net9740)
);

INV_X32 merge9190(
.A(net9916),
.ZN(net9741)
);

NAND2_X4 merge9191(
.A1(net5857),
.A2(net6858),
.ZN(net9742)
);

SDFFR_X1 merge9192(
.D(net7463),
.RN(net7271),
.SE(net5283),
.SI(net11093),
.CK(clk),
.Q(net9744),
.QN(net9743)
);

INV_X4 merge9193(
.A(net10221),
.ZN(net9745)
);

INV_X1 merge9194(
.A(net10527),
.ZN(net9746)
);

NAND3_X2 merge9195(
.A1(net4495),
.A2(net6397),
.A3(net5485),
.ZN(net9747)
);

DFFRS_X2 merge9196(
.D(net6228),
.RN(net7079),
.SN(net7167),
.CK(clk),
.Q(net9749),
.QN(net9748)
);

DFFR_X1 merge9197(
.D(net4975),
.RN(net5009),
.CK(clk),
.Q(net9751),
.QN(net9750)
);

SDFFR_X2 merge9198(
.D(net9196),
.RN(net7807),
.SE(net8246),
.SI(net8233),
.CK(clk),
.Q(net9753),
.QN(net9752)
);

DFFR_X2 merge9199(
.D(net1007),
.RN(net1016),
.CK(clk),
.Q(net9755),
.QN(net9754)
);

SDFFS_X1 merge9200(
.D(net6133),
.SE(net5524),
.SI(net4618),
.SN(net4524),
.CK(clk),
.Q(net9757),
.QN(net9756)
);

INV_X2 merge9201(
.A(net10304),
.ZN(net9758)
);

DFFS_X1 merge9202(
.D(net5811),
.SN(net5862),
.CK(clk),
.Q(net9760),
.QN(net9759)
);

INV_X8 merge9203(
.A(net10916),
.ZN(net9761)
);

SDFFS_X2 merge9204(
.D(net7546),
.SE(net8567),
.SI(net7431),
.SN(net9502),
.CK(clk),
.Q(net9763),
.QN(net9762)
);

INV_X16 merge9205(
.A(net10115),
.ZN(net9764)
);

INV_X32 merge9206(
.A(net10193),
.ZN(net9765)
);

INV_X4 merge9207(
.A(net10068),
.ZN(net9766)
);

INV_X1 merge9208(
.A(net10001),
.ZN(net9767)
);

OR3_X1 merge9209(
.A1(net6898),
.A2(net8842),
.A3(net7021),
.ZN(net9768)
);

AOI211_X4 merge9210(
.A(net3560),
.B(net1783),
.C1(net4620),
.C2(net3728),
.ZN(net9769)
);

SDFFR_X1 merge9211(
.D(net7098),
.RN(net5114),
.SE(net8090),
.SI(net8070),
.CK(clk),
.Q(net9771),
.QN(net9770)
);

INV_X2 merge9212(
.A(net10833),
.ZN(net9772)
);

DFFS_X2 merge9213(
.D(net2939),
.SN(net3845),
.CK(clk),
.Q(net9774),
.QN(net9773)
);

SDFFR_X2 merge9214(
.D(net8004),
.RN(net7994),
.SE(net8054),
.SI(net8118),
.CK(clk),
.Q(net9776),
.QN(net9775)
);

NOR4_X1 merge9215(
.A1(net5592),
.A2(net5612),
.A3(net5562),
.A4(net5597),
.ZN(net9777)
);

INV_X8 merge9216(
.A(net9981),
.ZN(net9778)
);

AOI211_X2 merge9217(
.A(net1363),
.B(net3969),
.C1(net4152),
.C2(net3081),
.ZN(net9779)
);

SDFFS_X1 merge9218(
.D(net4374),
.SE(net4368),
.SI(net3463),
.SN(net2593),
.CK(clk),
.Q(net9781),
.QN(net9780)
);

INV_X16 merge9219(
.A(net10085),
.ZN(net9782)
);

INV_X32 merge9220(
.A(net10960),
.ZN(net9783)
);

SDFFS_X2 merge9221(
.D(net8345),
.SE(net6460),
.SI(net4627),
.SN(net6381),
.CK(clk),
.Q(net9785),
.QN(net9784)
);

INV_X4 merge9222(
.A(net10939),
.ZN(net9786)
);

MUX2_X1 merge9223(
.A(net2564),
.B(net3639),
.S(net4524),
.Z(net9787)
);

INV_X1 merge9224(
.A(net10026),
.ZN(net9788)
);

INV_X2 merge9225(
.A(net9894),
.ZN(net9789)
);

CLKGATETST_X1 merge9226(
.E(net403),
.SE(net632),
.CK(clk),
.GCK(net9790)
);

SDFFR_X1 merge9227(
.D(net5144),
.RN(net2261),
.SE(net5148),
.SI(net4260),
.CK(clk),
.Q(net9792),
.QN(net9791)
);

INV_X8 merge9228(
.A(net10018),
.ZN(net9793)
);

SDFFR_X2 merge9229(
.D(net4611),
.RN(net4662),
.SE(net2587),
.SI(net2822),
.CK(clk),
.Q(net9795),
.QN(net9794)
);

SDFF_X1 merge9230(
.D(net5975),
.SE(net4994),
.SI(net5951),
.CK(clk),
.Q(net9797),
.QN(net9796)
);

SDFFS_X1 merge9231(
.D(net8169),
.SE(net8132),
.SI(net7200),
.SN(net8119),
.CK(clk),
.Q(net9799),
.QN(net9798)
);

SDFFS_X2 merge9232(
.D(net7282),
.SE(net7268),
.SI(net6353),
.SN(net6356),
.CK(clk),
.Q(net9801),
.QN(net9800)
);

SDFFR_X1 merge9233(
.D(net3600),
.RN(net3480),
.SE(net1700),
.SI(net2465),
.CK(clk),
.Q(net9803),
.QN(net9802)
);

CLKGATETST_X2 merge9234(
.E(net2942),
.SE(net1958),
.CK(clk),
.GCK(net9804)
);

SDFF_X2 merge9235(
.D(net8372),
.SE(net8139),
.SI(net8291),
.CK(clk),
.Q(net9806),
.QN(net9805)
);

CLKGATETST_X4 merge9236(
.E(net1434),
.SE(net1464),
.CK(clk),
.GCK(net9807)
);

CLKGATETST_X8 merge9237(
.E(net6739),
.SE(net5824),
.CK(clk),
.GCK(net9808)
);

AND2_X2 merge9238(
.A1(net450),
.A2(net1454),
.ZN(net9809)
);

SDFFR_X2 merge9239(
.D(net7371),
.RN(net5320),
.SE(net7207),
.SI(net6441),
.CK(clk),
.Q(net9811),
.QN(net9810)
);

DFFRS_X1 merge9240(
.D(net1416),
.RN(net2582),
.SN(net2581),
.CK(clk),
.Q(net9813),
.QN(net9812)
);

DFFR_X1 merge9241(
.D(net2923),
.RN(net3845),
.CK(clk),
.Q(net9815),
.QN(net9814)
);

SDFFS_X1 merge9242(
.D(net7876),
.SE(net6908),
.SI(net7139),
.SN(net7136),
.CK(clk),
.Q(net9817),
.QN(net9816)
);

DFFR_X2 merge9243(
.D(net7733),
.RN(net6739),
.CK(clk),
.Q(net9819),
.QN(net9818)
);

AOI22_X1 merge9244(
.A1(net2238),
.A2(net5067),
.B1(net4122),
.B2(net4070),
.ZN(net9820)
);

SDFFS_X2 merge9245(
.D(net7263),
.SE(net7260),
.SI(net9189),
.SN(net8946),
.CK(clk),
.Q(net9822),
.QN(net9821)
);

INV_X16 merge9246(
.A(net10005),
.ZN(net9823)
);

SDFFR_X1 merge9247(
.D(net6573),
.RN(net7554),
.SE(net5654),
.SI(net5590),
.CK(clk),
.Q(net9825),
.QN(net9824)
);

OAI21_X4 merge9248(
.A(net942),
.B1(net216),
.B2(net1274),
.ZN(net9826)
);

SDFFR_X2 merge9249(
.D(net8132),
.RN(net7199),
.SE(net6179),
.SI(net7204),
.CK(clk),
.Q(net9828),
.QN(net9827)
);

SDFFS_X1 merge9250(
.D(net1653),
.SE(net1660),
.SI(net3404),
.SN(net3479),
.CK(clk),
.Q(net9830),
.QN(net9829)
);

AND4_X4 merge9251(
.A1(net5528),
.A2(net6410),
.A3(net5557),
.A4(net5525),
.ZN(net9831)
);

XOR2_X1 merge9252(
.A(net6764),
.B(net5790),
.Z(net9832)
);

NAND4_X1 merge9253(
.A1(net2427),
.A2(net2324),
.A3(net2209),
.A4(net3125),
.ZN(net9833)
);

SDFFS_X2 merge9254(
.D(net7333),
.SE(net6534),
.SI(net9261),
.SN(net9149),
.CK(clk),
.Q(net9835),
.QN(net9834)
);

SDFFR_X1 merge9255(
.D(net5543),
.RN(net3448),
.SE(net6441),
.SI(net6391),
.CK(clk),
.Q(net9837),
.QN(net9836)
);

SDFFR_X2 merge9256(
.D(net1659),
.RN(net1672),
.SE(net732),
.SI(net85),
.CK(clk),
.Q(net9839),
.QN(net9838)
);

SDFFS_X1 merge9257(
.D(net8229),
.SE(net6158),
.SI(net8231),
.SN(net11208),
.CK(clk),
.Q(net9841),
.QN(net9840)
);

SDFFS_X2 merge9258(
.D(net2614),
.SE(net1670),
.SI(net1690),
.SN(net10882),
.CK(clk),
.Q(net9843),
.QN(net9842)
);

SDFFR_X1 merge9259(
.D(net5110),
.RN(net6054),
.SE(net3134),
.SI(net6951),
.CK(clk),
.Q(net9845),
.QN(net9844)
);

SDFFR_X2 merge9260(
.D(net7231),
.RN(net7810),
.SE(net6084),
.SI(net5345),
.CK(clk),
.Q(net9847),
.QN(net9846)
);

SDFFS_X1 merge9261(
.D(net8353),
.SE(net8370),
.SI(net4547),
.SN(net4556),
.CK(clk),
.Q(net9849),
.QN(net9848)
);

SDFFS_X2 merge9262(
.D(net7448),
.SE(net7539),
.SI(net7348),
.SN(net6337),
.CK(clk),
.Q(net9851),
.QN(net9850)
);

SDFFR_X1 merge9263(
.D(net8117),
.RN(net1270),
.SE(net4113),
.SI(net11130),
.CK(clk),
.Q(net9853),
.QN(net9852)
);

SDFFR_X2 merge9264(
.D(net6786),
.RN(net7288),
.SE(net7189),
.SI(net8283),
.CK(clk),
.Q(net9855),
.QN(net9854)
);

DFFS_X1 merge9265(
.D(net5771),
.SN(net2942),
.CK(clk),
.Q(net9857),
.QN(net9856)
);

OR4_X1 merge9266(
.A1(net3583),
.A2(net3562),
.A3(net3612),
.A4(net3305),
.ZN(net9858)
);

OAI22_X1 merge9267(
.A1(net6425),
.A2(net4471),
.B1(net8223),
.B2(net7908),
.ZN(net9859)
);

AND4_X2 merge9268(
.A1(net6093),
.A2(net6282),
.A3(net6212),
.A4(net6283),
.ZN(net9860)
);

SDFFS_X1 merge9269(
.D(net2501),
.SE(net2516),
.SI(net665),
.SN(net1604),
.CK(clk),
.Q(net9862),
.QN(net9861)
);

DFFRS_X2 merge9270(
.D(net2020),
.RN(net1114),
.SN(net3124),
.CK(clk),
.Q(net9864),
.QN(net9863)
);

DFFS_X2 merge9271(
.D(net1892),
.SN(net1923),
.CK(clk),
.Q(net9866),
.QN(net9865)
);

AND4_X1 merge9272(
.A1(net6491),
.A2(net6489),
.A3(net8013),
.A4(net8193),
.ZN(net9867)
);

AOI22_X4 merge9273(
.A1(net4287),
.A2(net2553),
.B1(net3344),
.B2(net4556),
.ZN(net9868)
);

OAI22_X4 merge9274(
.A1(net1701),
.A2(net1726),
.B1(net2625),
.B2(net1768),
.ZN(net9869)
);

SDFFS_X2 merge9275(
.D(net6428),
.SE(net6457),
.SI(net3571),
.SN(net3565),
.CK(clk),
.Q(net9871),
.QN(net9870)
);

AOI22_X2 merge9276(
.A1(net3625),
.A2(net3561),
.B1(net3626),
.B2(net4531),
.ZN(net9872)
);

SDFFR_X1 merge9277(
.D(net4076),
.RN(net4064),
.SE(net5053),
.SI(net10418),
.CK(clk),
.Q(net9874),
.QN(net9873)
);

NAND4_X4 merge9278(
.A1(net8402),
.A2(net4648),
.A3(net5580),
.A4(net10855),
.ZN(net9875)
);

OAI211_X2 merge9279(
.A(net309),
.B(net308),
.C1(net3048),
.C2(net3036),
.ZN(net9876)
);

SDFF_X1 merge9280(
.D(net7756),
.SE(net7893),
.SI(net5877),
.CK(clk),
.Q(net9878),
.QN(net9877)
);

OR4_X2 merge9281(
.A1(net552),
.A2(net515),
.A3(net456),
.A4(net10804),
.ZN(net9879)
);

AOI211_X1 merge9282(
.A(net63),
.B(net147),
.C1(net3051),
.C2(net1022),
.ZN(net9880)
);

SDFFR_X2 merge9283(
.D(net2642),
.RN(net3609),
.SE(net4549),
.SI(net4432),
.CK(clk),
.Q(net9882),
.QN(net9881)
);

NAND4_X2 merge9284(
.A1(net4005),
.A2(net3992),
.A3(net4152),
.A4(net10690),
.ZN(net9883)
);

OR4_X4 merge9285(
.A1(net748),
.A2(net1718),
.A3(net4563),
.A4(net3637),
.ZN(net9884)
);

SDFFS_X1 merge9286(
.D(net3319),
.SE(net2410),
.SI(net3367),
.SN(net2281),
.CK(clk),
.Q(net9886),
.QN(net9885)
);

OAI22_X2 merge9287(
.A1(net2095),
.A2(net1433),
.B1(net408),
.B2(net343),
.ZN(net9887)
);

SDFFS_X2 merge9288(
.D(net3101),
.SE(net4368),
.SI(net1407),
.SN(net1382),
.CK(clk),
.Q(net9889),
.QN(net9888)
);

OAI211_X4 merge9289(
.A(net128),
.B(net226),
.C1(net3927),
.C2(net3979),
.ZN(net9890)
);

SDFFR_X1 merge9290(
.D(net7095),
.RN(net6726),
.SE(net7010),
.SI(net4179),
.CK(clk),
.Q(net9892),
.QN(net9891)
);

SDFFR_X2 merge9291(
.D(net1754),
.RN(net732),
.SE(net816),
.SI(net821),
.CK(clk),
.Q(net9894),
.QN(net9893)
);

OAI211_X1 merge9292(
.A(net1193),
.B(net2188),
.C1(net1234),
.C2(net1023),
.ZN(net9895)
);

SDFFS_X1 merge9293(
.D(net3260),
.SE(net2549),
.SI(net515),
.SN(net512),
.CK(clk),
.Q(net9897),
.QN(net9896)
);

SDFFS_X2 merge9294(
.D(net5577),
.SE(net3758),
.SI(net7405),
.SN(net5480),
.CK(clk),
.Q(net9899),
.QN(net9898)
);

SDFFR_X1 merge9295(
.D(net3342),
.RN(net2285),
.SE(net4331),
.SI(net3969),
.CK(clk),
.Q(net9901),
.QN(net9900)
);

SDFFR_X2 merge9296(
.D(net6444),
.RN(net6253),
.SE(net8378),
.SI(net6391),
.CK(clk),
.Q(net9903),
.QN(net9902)
);

SDFFS_X1 merge9297(
.D(net6556),
.SE(net5574),
.SI(net6253),
.SN(net11026),
.CK(clk),
.Q(net9905),
.QN(net9904)
);

NOR4_X4 merge9298(
.A1(net8834),
.A2(net8822),
.A3(net8824),
.A4(net10744),
.ZN(net9906)
);

NOR4_X2 merge9299(
.A1(net6930),
.A2(net6904),
.A3(net6909),
.A4(net6911),
.ZN(net9907)
);

SDFFS_X2 merge9300(
.D(net7399),
.SE(net7288),
.SI(net7236),
.SN(net4145),
.CK(clk),
.Q(net9909),
.QN(net9908)
);

SDFFR_X1 merge9301(
.D(net4154),
.RN(net5070),
.SE(net5095),
.SI(net10800),
.CK(clk),
.Q(net9911),
.QN(net9910)
);

SDFFR_X2 merge9302(
.D(net4990),
.RN(net5053),
.SE(net6850),
.SI(net6898),
.CK(clk),
.Q(net9913),
.QN(net9912)
);

SDFFS_X1 merge9303(
.D(net7138),
.SE(net7127),
.SI(net6908),
.SN(net8101),
.CK(clk),
.Q(net9915),
.QN(net9914)
);

SDFFS_X2 merge9304(
.D(net5949),
.SE(net5951),
.SI(net3850),
.SN(net6988),
.CK(clk),
.Q(net9917),
.QN(net9916)
);

SDFFR_X1 merge9305(
.D(net5533),
.RN(net5580),
.SE(net8361),
.SI(net6534),
.CK(clk),
.Q(net9919),
.QN(net9918)
);

AOI211_X4 merge9306(
.A(net3595),
.B(net4556),
.C1(net1551),
.C2(net476),
.ZN(net9920)
);

SDFFR_X2 merge9307(
.D(net5999),
.RN(net6005),
.SE(net6942),
.SI(net6904),
.CK(clk),
.Q(net9922),
.QN(net9921)
);

NOR4_X1 merge9308(
.A1(net1506),
.A2(net1398),
.A3(net2500),
.A4(net2495),
.ZN(net9923)
);

AOI211_X2 merge9309(
.A(net5875),
.B(net5899),
.C1(net5783),
.C2(net2993),
.ZN(net9924)
);

SDFFS_X1 merge9310(
.D(net8749),
.SE(net8759),
.SI(net6855),
.SN(net6884),
.CK(clk),
.Q(net9926),
.QN(net9925)
);

SDFFS_X2 merge9311(
.D(net5852),
.SE(net3933),
.SI(net4950),
.SN(net4868),
.CK(clk),
.Q(net9928),
.QN(net9927)
);

SDFFR_X1 merge9312(
.D(net106),
.RN(net961),
.SE(net1042),
.SI(net1075),
.CK(clk),
.Q(net9930),
.QN(net9929)
);

SDFFR_X2 merge9313(
.D(net1840),
.RN(net1856),
.SE(net760),
.SI(net765),
.CK(clk),
.Q(net9932),
.QN(net9931)
);

SDFFS_X1 merge9314(
.D(net5177),
.SE(net3925),
.SI(net1383),
.SN(net1416),
.CK(clk),
.Q(net9934),
.QN(net9933)
);

AOI22_X1 merge9315(
.A1(net6222),
.A2(net7185),
.B1(net8021),
.B2(net11081),
.ZN(net9935)
);

AND4_X4 merge9316(
.A1(net2635),
.A2(net2648),
.A3(net3569),
.A4(net3447),
.ZN(net9936)
);

NAND4_X1 merge9317(
.A1(net6410),
.A2(net6116),
.A3(net5518),
.A4(net4432),
.ZN(net9937)
);

SDFFS_X2 merge9318(
.D(net4141),
.SE(net6970),
.SI(net8000),
.SN(net7708),
.CK(clk),
.Q(net9939),
.QN(net9938)
);

SDFFR_X1 merge9319(
.D(net454),
.RN(net458),
.SE(net2266),
.SI(net2209),
.CK(clk),
.Q(net9941),
.QN(net9940)
);

OR4_X1 merge9320(
.A1(net5260),
.A2(net5292),
.A3(net5289),
.A4(net6093),
.ZN(net9942)
);

OAI22_X1 merge9321(
.A1(net5190),
.A2(net6306),
.B1(net6996),
.B2(net6133),
.ZN(net9943)
);

AND4_X2 merge9322(
.A1(net8368),
.A2(net8239),
.A3(net7417),
.A4(net7420),
.ZN(net9944)
);

SDFFR_X2 merge9323(
.D(net6888),
.RN(net4961),
.SE(net5874),
.SI(net5805),
.CK(clk),
.Q(net9946),
.QN(net9945)
);

SDFFS_X1 merge9324(
.D(net6284),
.SE(net1526),
.SI(net551),
.SN(net10647),
.CK(clk),
.Q(net9948),
.QN(net9947)
);

AND4_X1 merge9325(
.A1(net6447),
.A2(net8268),
.A3(net9237),
.A4(net9293),
.ZN(net9949)
);

SDFFS_X2 merge9326(
.D(net2549),
.SE(net3397),
.SI(net1433),
.SN(net3543),
.CK(clk),
.Q(net9951),
.QN(net9950)
);

AOI22_X4 merge9327(
.A1(net3689),
.A2(net3653),
.B1(net2721),
.B2(net2733),
.ZN(net9952)
);

OAI22_X4 merge9328(
.A1(net7250),
.A2(net6474),
.B1(net6452),
.B2(net10780),
.ZN(net9953)
);

AOI22_X2 merge9329(
.A1(net4009),
.A2(net2103),
.B1(net4995),
.B2(net5027),
.ZN(net9954)
);

SDFFR_X1 merge9330(
.D(net268),
.RN(net25),
.SE(net1965),
.SI(net2103),
.CK(clk),
.Q(net9956),
.QN(net9955)
);

NAND4_X4 merge9331(
.A1(net6159),
.A2(net6158),
.A3(net1372),
.A4(net3209),
.ZN(net9957)
);

SDFFR_X2 merge9332(
.D(net7262),
.RN(net5389),
.SE(net2354),
.SI(net3178),
.CK(clk),
.Q(net9959),
.QN(net9958)
);

SDFFS_X1 merge9333(
.D(net6395),
.SE(net8319),
.SI(net7161),
.SN(net8035),
.CK(clk),
.Q(net9961),
.QN(net9960)
);

SDFFS_X2 merge9334(
.D(net5006),
.SE(net5022),
.SI(net5801),
.SN(net5050),
.CK(clk),
.Q(net9963),
.QN(net9962)
);

OAI211_X2 merge9335(
.A(net4650),
.B(net4531),
.C1(net5402),
.C2(net5403),
.ZN(net9964)
);

SDFFR_X1 merge9336(
.D(net5516),
.RN(net5531),
.SE(net3789),
.SI(net5691),
.CK(clk),
.Q(net9966),
.QN(net9965)
);

SDFFR_X2 merge9337(
.D(net6385),
.RN(net6596),
.SE(net5485),
.SI(net5482),
.CK(clk),
.Q(net9968),
.QN(net9967)
);

SDFFS_X1 merge9338(
.D(net3458),
.SE(net3414),
.SI(net584),
.SN(net546),
.CK(clk),
.Q(net9970),
.QN(net9969)
);

SDFFS_X2 merge9339(
.D(net3015),
.SE(net3013),
.SI(net3091),
.SN(net3085),
.CK(clk),
.Q(net9972),
.QN(net9971)
);

OR4_X2 merge9340(
.A1(net950),
.A2(net2046),
.A3(net147),
.A4(net2943),
.ZN(net9973)
);

SDFFR_X1 merge9341(
.D(net7278),
.RN(net7101),
.SE(net6451),
.SI(net6452),
.CK(clk),
.Q(net9975),
.QN(net9974)
);

SDFFR_X2 merge9342(
.D(net9120),
.RN(net8139),
.SE(net9179),
.SI(net9295),
.CK(clk),
.Q(net9977),
.QN(net9976)
);

AOI211_X1 merge9343(
.A(net1055),
.B(net1092),
.C1(net1994),
.C2(net2046),
.ZN(net9978)
);

SDFFS_X1 merge9344(
.D(net1177),
.SE(net4174),
.SI(net4213),
.SN(net4108),
.CK(clk),
.Q(net9980),
.QN(net9979)
);

SDFFS_X2 merge9345(
.D(net987),
.SE(net1292),
.SI(net1094),
.SN(net1280),
.CK(clk),
.Q(net9982),
.QN(net9981)
);

SDFFR_X1 merge9346(
.D(net1022),
.RN(net318),
.SE(net269),
.SI(net1116),
.CK(clk),
.Q(net9984),
.QN(net9983)
);

NAND4_X2 merge9347(
.A1(net5849),
.A2(net6182),
.A3(net8091),
.A4(net7005),
.ZN(net9985)
);

SDFFR_X2 merge9348(
.D(net4601),
.RN(net5474),
.SE(net4457),
.SI(net4638),
.CK(clk),
.Q(net9987),
.QN(net9986)
);

OR4_X4 merge9349(
.A1(net403),
.A2(net1398),
.A3(net6117),
.A4(net6119),
.ZN(net9988)
);

SDFFS_X1 merge9350(
.D(net4275),
.SE(net4531),
.SI(net2691),
.SN(net2656),
.CK(clk),
.Q(net9990),
.QN(net9989)
);

SDFFS_X2 merge9351(
.D(net1239),
.SE(net1233),
.SI(net1064),
.SN(net2148),
.CK(clk),
.Q(net9992),
.QN(net9991)
);

OAI22_X2 merge9352(
.A1(net3190),
.A2(net3198),
.B1(net1251),
.B2(net4100),
.ZN(net9993)
);

SDFFR_X1 merge9353(
.D(net6783),
.RN(net5025),
.SE(net6908),
.SI(net10909),
.CK(clk),
.Q(net9995),
.QN(net9994)
);

SDFFR_X2 merge9354(
.D(net6463),
.RN(net6303),
.SE(net2590),
.SI(net3459),
.CK(clk),
.Q(net9997),
.QN(net9996)
);

SDFFS_X1 merge9355(
.D(net7910),
.SE(net8760),
.SI(net8855),
.SN(net8824),
.CK(clk),
.Q(net9999),
.QN(net9998)
);

SDFFS_X2 merge9356(
.D(net7726),
.SE(net3979),
.SI(net6981),
.SN(net6979),
.CK(clk),
.Q(net10001),
.QN(net10000)
);

SDFFR_X1 merge9357(
.D(net2475),
.RN(net2455),
.SE(net3417),
.SI(net3260),
.CK(clk),
.Q(net10003),
.QN(net10002)
);

OAI211_X4 merge9358(
.A(net3584),
.B(net2687),
.C1(net2707),
.C2(net10972),
.ZN(net10004)
);

SDFFR_X2 merge9359(
.D(net2013),
.RN(net1920),
.SE(net2068),
.SI(net1124),
.CK(clk),
.Q(net10006),
.QN(net10005)
);

OAI211_X1 merge9360(
.A(net3527),
.B(net3515),
.C1(net4372),
.C2(net4494),
.ZN(net10007)
);

SDFFS_X1 merge9361(
.D(net6868),
.SE(net6896),
.SI(net5856),
.SN(net5871),
.CK(clk),
.Q(net10009),
.QN(net10008)
);

NOR4_X4 merge9362(
.A1(net5227),
.A2(net6120),
.A3(net2382),
.A4(net2381),
.ZN(net10010)
);

NOR4_X2 merge9363(
.A1(net1718),
.A2(net1714),
.A3(net3598),
.A4(net3582),
.ZN(net10011)
);

SDFFS_X2 merge9364(
.D(net4966),
.SE(net4057),
.SI(net5955),
.SN(net5951),
.CK(clk),
.Q(net10013),
.QN(net10012)
);

AOI211_X4 merge9365(
.A(net1789),
.B(net2696),
.C1(net891),
.C2(net913),
.ZN(net10014)
);

SDFFR_X1 merge9366(
.D(net5156),
.RN(net8089),
.SE(net9027),
.SI(net10864),
.CK(clk),
.Q(net10016),
.QN(net10015)
);

SDFFR_X2 merge9367(
.D(net476),
.RN(net663),
.SE(net3495),
.SI(net2423),
.CK(clk),
.Q(net10018),
.QN(net10017)
);

SDFFS_X1 merge9368(
.D(net6137),
.SE(net6179),
.SI(net5231),
.SN(net5103),
.CK(clk),
.Q(net10020),
.QN(net10019)
);

SDFFS_X2 merge9369(
.D(net6417),
.SE(net6412),
.SI(net7417),
.SN(net11050),
.CK(clk),
.Q(net10022),
.QN(net10021)
);

NOR4_X1 merge9370(
.A1(net414),
.A2(net863),
.A3(net3522),
.A4(net3396),
.ZN(net10023)
);

SDFFR_X1 merge9371(
.D(net4430),
.RN(net5429),
.SE(net5459),
.SI(net6337),
.CK(clk),
.Q(net10025),
.QN(net10024)
);

SDFFR_X2 merge9372(
.D(net3208),
.RN(net1322),
.SE(net410),
.SI(net454),
.CK(clk),
.Q(net10027),
.QN(net10026)
);

SDFFS_X1 merge9373(
.D(net5366),
.SE(net4382),
.SI(net2455),
.SN(net2317),
.CK(clk),
.Q(net10029),
.QN(net10028)
);

SDFFS_X2 merge9374(
.D(net4886),
.SE(net5031),
.SI(net5856),
.SN(net11196),
.CK(clk),
.Q(net10031),
.QN(net10030)
);

SDFFR_X1 merge9375(
.D(net7461),
.RN(net7448),
.SE(net7379),
.SI(net7430),
.CK(clk),
.Q(net10033),
.QN(net10032)
);

AOI211_X2 merge9376(
.A(net2368),
.B(net2382),
.C1(net4481),
.C2(net4425),
.ZN(net10034)
);

SDFFR_X2 merge9377(
.D(net4368),
.RN(net6337),
.SE(net8262),
.SI(net8248),
.CK(clk),
.Q(net10036),
.QN(net10035)
);

AOI22_X1 merge9378(
.A1(net5469),
.A2(net6434),
.B1(net7035),
.B2(net6158),
.ZN(net10037)
);

SDFFS_X1 merge9379(
.D(net6931),
.SE(net6973),
.SI(net6749),
.SN(net6872),
.CK(clk),
.Q(net10039),
.QN(net10038)
);

SDFFS_X2 merge9380(
.D(net6172),
.SE(net6286),
.SI(net8171),
.SN(net6086),
.CK(clk),
.Q(net10041),
.QN(net10040)
);

AND4_X4 merge9381(
.A1(net1436),
.A2(net1396),
.A3(net1584),
.A4(net2613),
.ZN(net10042)
);

SDFFR_X1 merge9382(
.D(net9295),
.RN(net5476),
.SE(net5555),
.SI(net10383),
.CK(clk),
.Q(net10044),
.QN(net10043)
);

SDFFR_X2 merge9383(
.D(net6147),
.RN(net6116),
.SE(net7411),
.SI(net7399),
.CK(clk),
.Q(net10046),
.QN(net10045)
);

SDFFS_X1 merge9384(
.D(net2153),
.SE(net1174),
.SI(net1023),
.SN(net10665),
.CK(clk),
.Q(net10048),
.QN(net10047)
);

SDFFS_X2 merge9385(
.D(net2606),
.SE(net2613),
.SI(net2333),
.SN(net2332),
.CK(clk),
.Q(net10050),
.QN(net10049)
);

SDFFR_X1 merge9386(
.D(net8165),
.RN(net8197),
.SE(net6401),
.SI(net6116),
.CK(clk),
.Q(net10052),
.QN(net10051)
);

NAND4_X1 merge9387(
.A1(net267),
.A2(net287),
.A3(net3044),
.A4(net3024),
.ZN(net10053)
);

OR4_X1 merge9388(
.A1(net5464),
.A2(net5480),
.A3(net4425),
.A4(net5315),
.ZN(net10054)
);

SDFFR_X2 merge9389(
.D(net3469),
.RN(net5326),
.SE(net5605),
.SI(net2732),
.CK(clk),
.Q(net10056),
.QN(net10055)
);

SDFFS_X1 merge9390(
.D(net2278),
.SE(net2288),
.SI(net211),
.SN(net1092),
.CK(clk),
.Q(net10058),
.QN(net10057)
);

SDFFS_X2 merge9391(
.D(net7905),
.SE(net7704),
.SI(net5983),
.SN(net6959),
.CK(clk),
.Q(net10060),
.QN(net10059)
);

OAI22_X1 merge9392(
.A1(net2978),
.A2(net3092),
.B1(net3116),
.B2(net3032),
.ZN(net10061)
);

AND4_X2 merge9393(
.A1(net2385),
.A2(net3291),
.A3(net3374),
.A4(net3380),
.ZN(net10062)
);

SDFFR_X1 merge9394(
.D(net7924),
.RN(net7864),
.SE(net8872),
.SI(net8708),
.CK(clk),
.Q(net10064),
.QN(net10063)
);

SDFFR_X2 merge9395(
.D(net6048),
.RN(net6038),
.SE(net4147),
.SI(net5139),
.CK(clk),
.Q(net10066),
.QN(net10065)
);

SDFFS_X1 merge9396(
.D(net3291),
.SE(net3313),
.SI(net3513),
.SN(net4495),
.CK(clk),
.Q(net10068),
.QN(net10067)
);

AND4_X1 merge9397(
.A1(net3593),
.A2(net2475),
.A3(net3603),
.A4(net2678),
.ZN(net10069)
);

AOI22_X4 merge9398(
.A1(net2597),
.A2(net3571),
.B1(net4624),
.B2(net1579),
.ZN(net10070)
);

OAI22_X4 merge9399(
.A1(net4989),
.A2(net5053),
.B1(net1449),
.B2(net3375),
.ZN(net10071)
);

SDFFS_X2 merge9400(
.D(net6189),
.SE(net5185),
.SI(net5238),
.SN(net5206),
.CK(clk),
.Q(net10073),
.QN(net10072)
);

AOI22_X2 merge9401(
.A1(net4039),
.A2(net4009),
.B1(net4008),
.B2(net3884),
.ZN(net10074)
);

SDFFR_X1 merge9402(
.D(net4064),
.RN(net5898),
.SE(net7915),
.SI(net7922),
.CK(clk),
.Q(net10076),
.QN(net10075)
);

NAND4_X4 merge9403(
.A1(net447),
.A2(net442),
.A3(net5208),
.A4(net6120),
.ZN(net10077)
);

SDFFR_X2 merge9404(
.D(net7029),
.RN(net7161),
.SE(net6965),
.SI(net6964),
.CK(clk),
.Q(net10079),
.QN(net10078)
);

SDFFS_X1 merge9405(
.D(net5217),
.SE(net6130),
.SI(net5229),
.SN(net5262),
.CK(clk),
.Q(net10081),
.QN(net10080)
);

OAI211_X2 merge9406(
.A(net7351),
.B(net6460),
.C1(net8896),
.C2(net8912),
.ZN(net10082)
);

OR4_X2 merge9407(
.A1(net546),
.A2(net551),
.A3(net553),
.A4(net1408),
.ZN(net10083)
);

SDFFS_X2 merge9408(
.D(net1482),
.SE(net626),
.SI(net1585),
.SN(net1556),
.CK(clk),
.Q(net10085),
.QN(net10084)
);

SDFFR_X1 merge9409(
.D(net4492),
.RN(net6425),
.SE(net6484),
.SI(net5474),
.CK(clk),
.Q(net10087),
.QN(net10086)
);

SDFFR_X2 merge9410(
.D(net4766),
.RN(net5412),
.SE(net3467),
.SI(net3532),
.CK(clk),
.Q(net10089),
.QN(net10088)
);

AOI211_X1 merge9411(
.A(net4015),
.B(net4009),
.C1(net4052),
.C2(net4034),
.ZN(net10090)
);

NAND4_X2 merge9412(
.A1(net752),
.A2(net754),
.A3(net1711),
.A4(net1615),
.ZN(net10091)
);

OR4_X4 merge9413(
.A1(net3189),
.A2(net4485),
.A3(net4494),
.A4(net11160),
.ZN(net10092)
);

OAI22_X2 merge9414(
.A1(net3084),
.A2(net4086),
.B1(net5084),
.B2(net5058),
.ZN(net10093)
);

OAI211_X4 merge9415(
.A(net4106),
.B(net3151),
.C1(net4159),
.C2(net5095),
.ZN(net10094)
);

MUX2_X2 merge9416(
.A(net1212),
.B(net3133),
.S(net4099),
.Z(net10095)
);

OAI211_X1 merge9417(
.A(net5775),
.B(net5780),
.C1(net5924),
.C2(net5922),
.ZN(net10096)
);

SDFFS_X1 merge9418(
.D(net1710),
.SE(net2624),
.SI(net2477),
.SN(net2613),
.CK(clk),
.Q(net10098),
.QN(net10097)
);

SDFFS_X2 merge9419(
.D(net1543),
.SE(net4451),
.SI(net3396),
.SN(net11164),
.CK(clk),
.Q(net10100),
.QN(net10099)
);

SDFFR_X1 merge9420(
.D(net6118),
.RN(net3247),
.SE(net7862),
.SI(net8021),
.CK(clk),
.Q(net10102),
.QN(net10101)
);

NOR4_X4 merge9421(
.A1(net1103),
.A2(net3037),
.A3(net3120),
.A4(net4107),
.ZN(net10103)
);

SDFF_X2 merge9422(
.D(net4580),
.SE(net1683),
.SI(net3571),
.CK(clk),
.Q(net10105),
.QN(net10104)
);

NOR4_X2 merge9423(
.A1(net2360),
.A2(net2451),
.A3(net503),
.A4(net1268),
.ZN(net10106)
);

DFFRS_X1 merge9424(
.D(net3178),
.RN(net421),
.SN(net3310),
.CK(clk),
.Q(net10108),
.QN(net10107)
);

AOI211_X4 merge9425(
.A(net4041),
.B(net3056),
.C1(net4100),
.C2(net4213),
.ZN(net10109)
);

NOR4_X1 merge9426(
.A1(net1936),
.A2(net3069),
.A3(net3989),
.A4(net2990),
.ZN(net10110)
);

SDFFR_X2 merge9427(
.D(net3892),
.RN(net4884),
.SE(net3988),
.SI(net4893),
.CK(clk),
.Q(net10112),
.QN(net10111)
);

AOI211_X2 merge9428(
.A(net6964),
.B(net6987),
.C1(net6251),
.C2(net6295),
.ZN(net10113)
);

SDFFS_X1 merge9429(
.D(net1758),
.SE(net1752),
.SI(net3623),
.SN(net4546),
.CK(clk),
.Q(net10115),
.QN(net10114)
);

SDFFS_X2 merge9430(
.D(net6085),
.SE(net6103),
.SI(net7030),
.Q(net6989),
.CK(clk),
.QN(net10116)
);

SDFFR_X1 merge9431(
.D(net7061),
.RN(net7081),
.SE(net5143),
.SI(net5190),
.CK(clk),
.Q(net10119),
.QN(net10118)
);

SDFFR_X2 merge9432(
.D(net5309),
.RN(net2484),
.SE(net670),
.SI(net711),
.CK(clk),
.Q(net10121),
.QN(net10120)
);

SDFFS_X1 merge9433(
.D(net5283),
.SE(net8156),
.SI(net8242),
.SN(net11099),
.CK(clk),
.Q(net10123),
.QN(net10122)
);

AOI22_X1 merge9434(
.A1(net360),
.A2(net396),
.B1(net1292),
.B2(net1343),
.ZN(net10124)
);

SDFFS_X2 merge9435(
.D(net4285),
.SE(net4462),
.SI(net4502),
.SN(net4495),
.CK(clk),
.Q(net10126),
.QN(net10125)
);

AND4_X4 merge9436(
.A1(net3386),
.A2(net551),
.A3(net1660),
.A4(net1652),
.ZN(net10127)
);

SDFFR_X1 merge9437(
.D(net2148),
.RN(net2021),
.SE(net2146),
.SI(net2046),
.CK(clk),
.Q(net10129),
.QN(net10128)
);

SDFFR_X2 merge9438(
.D(net584),
.RN(net488),
.SE(net908),
.SI(net878),
.CK(clk),
.Q(net10131),
.QN(net10130)
);

SDFFS_X1 merge9439(
.D(net4204),
.SE(net4221),
.SI(net481),
.SN(net458),
.CK(clk),
.Q(net10133),
.QN(net10132)
);

NAND4_X1 merge9440(
.A1(net3262),
.A2(net3260),
.A3(net4201),
.A4(net4100),
.ZN(net10134)
);

OR4_X1 merge9441(
.A1(net3069),
.A2(net2863),
.A3(net4045),
.A4(net2090),
.ZN(net10135)
);

SDFFS_X2 merge9442(
.D(net3110),
.SE(net3060),
.SI(net4915),
.SN(net4885),
.CK(clk),
.Q(net10137),
.QN(net10136)
);

SDFFR_X1 merge9443(
.D(net2806),
.RN(net2828),
.SE(net3685),
.SI(net10509),
.CK(clk),
.Q(net10139),
.QN(net10138)
);

OAI22_X1 merge9444(
.A1(net2525),
.A2(net1627),
.B1(net4484),
.B2(net4500),
.ZN(net10140)
);

SDFFR_X2 merge9445(
.D(net4691),
.RN(net5639),
.SE(net5335),
.SI(net5199),
.CK(clk),
.Q(net10142),
.QN(net10141)
);

SDFFS_X1 merge9446(
.D(net2409),
.SE(net1593),
.SI(net6623),
.SN(net10478),
.CK(clk),
.Q(net10144),
.QN(net10143)
);

AND4_X2 merge9447(
.A1(net4397),
.A2(net4462),
.A3(net3552),
.A4(net5454),
.ZN(net10145)
);

SDFFS_X2 merge9448(
.D(net7869),
.SE(net8838),
.SI(net5877),
.SN(net7768),
.CK(clk),
.Q(net10147),
.QN(net10146)
);

SDFFR_X1 merge9449(
.D(net6097),
.RN(net6077),
.SE(net7859),
.SI(net7825),
.CK(clk),
.Q(net10149),
.QN(net10148)
);

SDFFR_X2 merge9450(
.D(net7266),
.RN(net7283),
.SE(net2530),
.SI(net643),
.CK(clk),
.Q(net10151),
.QN(net10150)
);

SDFFS_X1 merge9451(
.D(net4189),
.SE(net5233),
.SI(net5290),
.SN(net5185),
.CK(clk),
.Q(net10153),
.QN(net10152)
);

SDFFS_X2 merge9452(
.D(net476),
.SE(net1626),
.SI(net1590),
.SN(net665),
.CK(clk),
.Q(net10155),
.QN(net10154)
);

AND4_X1 merge9453(
.A1(net269),
.A2(net267),
.A3(net2364),
.A4(net3144),
.ZN(net10156)
);

SDFFR_X1 merge9454(
.D(net8100),
.RN(net5167),
.SE(net3425),
.SI(net1380),
.CK(clk),
.Q(net10158),
.QN(net10157)
);

SDFFR_X2 merge9455(
.D(net8204),
.RN(net8241),
.SE(net7929),
.SI(net8833),
.CK(clk),
.Q(net10160),
.QN(net10159)
);

SDFFS_X1 merge9456(
.D(net7346),
.SE(net6284),
.SI(net6196),
.SN(net6310),
.CK(clk),
.Q(net10162),
.QN(net10161)
);

AOI22_X4 merge9457(
.A1(net1264),
.A2(net1288),
.B1(net3421),
.B2(net3448),
.ZN(net10163)
);

OAI22_X4 merge9458(
.A1(net7019),
.A2(net6936),
.B1(net6073),
.B2(net6056),
.ZN(net10164)
);

SDFFS_X2 merge9459(
.D(net5033),
.SE(net4716),
.SI(net8280),
.SN(net5411),
.CK(clk),
.Q(net10166),
.QN(net10165)
);

AOI22_X2 merge9460(
.A1(net7765),
.A2(net7864),
.B1(net7949),
.B2(net5053),
.ZN(net10167)
);

NAND4_X4 merge9461(
.A1(net1657),
.A2(net1660),
.A3(net3479),
.A4(net3581),
.ZN(net10168)
);

SDFFR_X1 merge9462(
.D(net3742),
.RN(net3570),
.SE(net3392),
.SI(net10858),
.CK(clk),
.Q(net10170),
.QN(net10169)
);

SDFFR_X2 merge9463(
.D(net160),
.RN(net1117),
.SE(net3941),
.SI(net3896),
.CK(clk),
.Q(net10172),
.QN(net10171)
);

SDFFS_X1 merge9464(
.D(net2113),
.SE(net2126),
.SI(net3865),
.SN(net3884),
.CK(clk),
.Q(net10174),
.QN(net10173)
);

SDFFS_X2 merge9465(
.D(net1064),
.SE(net1011),
.SI(net996),
.SN(net1016),
.CK(clk),
.Q(net10176),
.QN(net10175)
);

OAI211_X2 merge9466(
.A(net1305),
.B(net1311),
.C1(net4353),
.C2(net4360),
.ZN(net10177)
);

SDFFR_X1 merge9467(
.D(net6136),
.RN(net4011),
.SE(net1401),
.SI(net1410),
.CK(clk),
.Q(net10179),
.QN(net10178)
);

SDFFR_X2 merge9468(
.D(net7558),
.RN(net6593),
.SE(net5172),
.SI(net5645),
.CK(clk),
.Q(net10181),
.QN(net10180)
);

SDFFS_X1 merge9469(
.D(net6765),
.SE(net6861),
.SI(net8002),
.SN(net7970),
.CK(clk),
.Q(net10183),
.QN(net10182)
);

OR4_X2 merge9470(
.A1(net4868),
.A2(net4894),
.A3(net4837),
.A4(net4893),
.ZN(net10184)
);

SDFFS_X2 merge9471(
.D(net3544),
.SE(net3536),
.SI(net6256),
.SN(net5459),
.CK(clk),
.Q(net10186),
.QN(net10185)
);

SDFFR_X1 merge9472(
.D(net6758),
.RN(net7151),
.SE(net7758),
.SI(net6979),
.CK(clk),
.Q(net10188),
.QN(net10187)
);

AOI211_X1 merge9473(
.A(net1719),
.B(net1730),
.C1(net5461),
.C2(net5495),
.ZN(net10189)
);

SDFFR_X2 merge9474(
.D(net4320),
.RN(net3292),
.SE(net3069),
.SI(net4997),
.CK(clk),
.Q(net10191),
.QN(net10190)
);

SDFFS_X1 merge9475(
.D(net1395),
.SE(net609),
.SI(net3442),
.SN(net3421),
.CK(clk),
.Q(net10193),
.QN(net10192)
);

NAND4_X2 merge9476(
.A1(net2690),
.A2(net2569),
.A3(net805),
.A4(net766),
.ZN(net10194)
);

OR4_X4 merge9477(
.A1(net3229),
.A2(net3306),
.A3(net4981),
.A4(net4994),
.ZN(net10195)
);

SDFFS_X2 merge9478(
.D(net6309),
.SE(net6235),
.SI(net631),
.SN(net578),
.CK(clk),
.Q(net10197),
.QN(net10196)
);

SDFFR_X1 merge9479(
.D(net286),
.RN(net291),
.SE(net6954),
.SI(net6968),
.CK(clk),
.Q(net10199),
.QN(net10198)
);

OAI22_X2 merge9480(
.A1(net142),
.A2(net1916),
.B1(net277),
.B2(net1300),
.ZN(net10200)
);

SDFFR_X2 merge9481(
.D(net3145),
.RN(net3107),
.SE(net1767),
.SI(net1793),
.CK(clk),
.Q(net10202),
.QN(net10201)
);

SDFFS_X1 merge9482(
.D(net6763),
.SE(net6988),
.SI(net7952),
.SN(net6020),
.CK(clk),
.Q(net10204),
.QN(net10203)
);

SDFFS_X2 merge9483(
.D(net1507),
.SE(net4368),
.SI(net3112),
.SN(net2112),
.CK(clk),
.Q(net10206),
.QN(net10205)
);

OAI211_X4 merge9484(
.A(net3161),
.B(net3133),
.C1(net5325),
.C2(net7309),
.ZN(net10207)
);

OAI211_X1 merge9485(
.A(net5082),
.B(net8081),
.C1(net11015),
.C2(net11095),
.ZN(net10208)
);

SDFFR_X1 merge9486(
.D(net3710),
.RN(net3704),
.SE(net873),
.SI(net858),
.CK(clk),
.Q(net10210),
.QN(net10209)
);

NOR4_X4 merge9487(
.A1(net261),
.A2(net302),
.A3(net3475),
.A4(net2570),
.ZN(net10211)
);

SDFFR_X2 merge9488(
.D(net2317),
.RN(net2337),
.SE(net3394),
.SI(net1381),
.CK(clk),
.Q(net10213),
.QN(net10212)
);

NOR4_X2 merge9489(
.A1(net3222),
.A2(net4295),
.A3(net418),
.A4(net1372),
.ZN(net10214)
);

AOI211_X4 merge9490(
.A(net4334),
.B(net4245),
.C1(net8021),
.C2(net11206),
.ZN(net10215)
);

SDFFS_X1 merge9491(
.D(net7902),
.SE(net7704),
.SI(net8805),
.SN(net7922),
.CK(clk),
.Q(net10217),
.QN(net10216)
);

SDFFS_X2 merge9492(
.D(net909),
.SE(net878),
.SI(net6371),
.SN(net6185),
.CK(clk),
.Q(net10219),
.QN(net10218)
);

NOR4_X1 merge9493(
.A1(net114),
.A2(net3091),
.A3(net3330),
.A4(net3296),
.ZN(net10220)
);

SDFFR_X1 merge9494(
.D(net3441),
.RN(net3413),
.SE(net289),
.SI(net2977),
.CK(clk),
.Q(net10222),
.QN(net10221)
);

AOI211_X2 merge9495(
.A(net3637),
.B(net4576),
.C1(net4478),
.C2(net4526),
.ZN(net10223)
);

AOI22_X1 merge9496(
.A1(net2192),
.A2(net1219),
.B1(net3144),
.B2(net10979),
.ZN(net10224)
);

AND4_X4 merge9497(
.A1(net793),
.A2(net788),
.A3(net7109),
.A4(net6425),
.ZN(net10225)
);

SDFFR_X2 merge9498(
.D(net4494),
.RN(net5385),
.SE(net551),
.SI(net3554),
.CK(clk),
.Q(net10227),
.QN(net10226)
);

NAND4_X1 merge9499(
.A1(net3374),
.A2(net2478),
.A3(net5074),
.A4(net5082),
.ZN(net10228)
);

OR4_X1 merge9500(
.A1(net5322),
.A2(net5220),
.A3(net1093),
.A4(net2491),
.ZN(net10229)
);

SDFFS_X1 merge9501(
.D(net5036),
.SE(net3364),
.SI(net4330),
.SN(net4333),
.CK(clk),
.Q(net10231),
.QN(net10230)
);

SDFFS_X2 merge9502(
.D(net4455),
.SE(net4457),
.SI(net9005),
.SN(net8975),
.CK(clk),
.Q(net10233),
.QN(net10232)
);

SDFFR_X1 merge9503(
.D(net3070),
.RN(net228),
.SE(net2352),
.SI(net1445),
.CK(clk),
.Q(net10235),
.QN(net10234)
);

OAI22_X1 merge9504(
.A1(net5447),
.A2(net5430),
.B1(net7328),
.B2(net5411),
.ZN(net10236)
);

SDFFR_X2 merge9505(
.D(net3558),
.RN(net2597),
.SE(net4150),
.SI(net5045),
.CK(clk),
.Q(net10238),
.QN(net10237)
);

AND4_X2 merge9506(
.A1(net5002),
.A2(net4016),
.A3(net4154),
.A4(net4097),
.ZN(net10239)
);

SDFFS_X1 merge9507(
.D(net8948),
.SE(net8926),
.SI(net8764),
.SN(net8017),
.CK(clk),
.Q(net10241),
.QN(net10240)
);

SDFFS_X2 merge9508(
.D(net2505),
.SE(net2448),
.SI(net156),
.SN(net277),
.CK(clk),
.Q(net10243),
.QN(net10242)
);

SDFFR_X1 merge9509(
.D(net7102),
.RN(net6283),
.SE(net6599),
.SI(net6558),
.CK(clk),
.Q(net10245),
.QN(net10244)
);

SDFFR_X2 merge9510(
.D(net2835),
.RN(net3742),
.SE(net6333),
.SI(net5283),
.CK(clk),
.Q(net10247),
.QN(net10246)
);

AND4_X1 merge9511(
.A1(net2504),
.A2(net2110),
.A3(net270),
.A4(net267),
.ZN(net10248)
);

SDFFS_X1 merge9512(
.D(net6403),
.SE(net6197),
.SI(net1533),
.SN(net1678),
.CK(clk),
.Q(net10250),
.QN(net10249)
);

AOI22_X4 merge9513(
.A1(net1315),
.A2(net3208),
.B1(net3184),
.B2(net3187),
.ZN(net10251)
);

SDFFS_X2 merge9514(
.D(net1190),
.SE(net2140),
.SI(net3038),
.SN(net1040),
.CK(clk),
.Q(net10253),
.QN(net10252)
);

SDFFR_X1 merge9515(
.D(net5873),
.RN(net5877),
.SE(net2254),
.SI(net2261),
.CK(clk),
.Q(net10255),
.QN(net10254)
);

SDFFR_X2 merge9516(
.D(net913),
.RN(net762),
.SE(net4478),
.SI(net10595),
.CK(clk),
.Q(net10257),
.QN(net10256)
);

SDFFS_X1 merge9517(
.D(net4068),
.SE(net4048),
.SI(net5171),
.SN(net5239),
.CK(clk),
.Q(net10259),
.QN(net10258)
);

SDFFS_X2 merge9518(
.D(net4030),
.SE(net5158),
.SI(net5917),
.SN(net5857),
.CK(clk),
.Q(net10261),
.QN(net10260)
);

SDFFR_X1 merge9519(
.D(net6071),
.RN(net6133),
.SE(net4202),
.SI(net6786),
.CK(clk),
.Q(net10263),
.QN(net10262)
);

SDFFR_X2 merge9520(
.D(net4525),
.RN(net4503),
.SE(net4798),
.SI(net5209),
.CK(clk),
.Q(net10265),
.QN(net10264)
);

SDFFS_X1 merge9521(
.D(net7987),
.SE(net8091),
.SI(net4454),
.SN(net5471),
.CK(clk),
.Q(net10267),
.QN(net10266)
);

SDFFS_X2 merge9522(
.D(net8065),
.SE(net8059),
.SI(net6303),
.SN(net4578),
.CK(clk),
.Q(net10269),
.QN(net10268)
);

SDFFR_X1 merge9523(
.D(net751),
.RN(net2584),
.SE(net2433),
.SI(net3477),
.CK(clk),
.Q(net10271),
.QN(net10270)
);

SDFFR_X2 merge9524(
.D(net5391),
.RN(net5328),
.SE(net2738),
.SI(net920),
.CK(clk),
.Q(net10273),
.QN(net10272)
);

OAI22_X4 merge9525(
.A1(net4436),
.A2(net5249),
.B1(net3169),
.B2(net7214),
.ZN(net10274)
);

AOI22_X2 merge9526(
.A1(net6830),
.A2(net6904),
.B1(net1438),
.B2(net1464),
.ZN(net10275)
);

SDFFS_X1 merge9527(
.D(net6283),
.SE(net7309),
.SI(net5235),
.SN(net2473),
.CK(clk),
.Q(net10277),
.QN(net10276)
);

SDFFS_X2 merge9528(
.D(net1871),
.SE(net2774),
.SI(net5449),
.SN(net5444),
.CK(clk),
.Q(net10279),
.QN(net10278)
);

NAND4_X4 merge9529(
.A1(net1385),
.A2(net458),
.A3(net4118),
.A4(net4295),
.ZN(net10280)
);

SDFFR_X1 merge9530(
.D(net8960),
.RN(net8956),
.SE(net4174),
.SI(net1200),
.CK(clk),
.Q(net10282),
.QN(net10281)
);

SDFFR_X2 merge9531(
.D(net6378),
.RN(net5431),
.SE(net679),
.SI(net506),
.CK(clk),
.Q(net10284),
.QN(net10283)
);

OAI211_X2 merge9532(
.A(net7332),
.B(net7227),
.C1(net5463),
.C2(net5454),
.ZN(net10285)
);

SDFFS_X1 merge9533(
.D(net2663),
.SE(net2653),
.SI(net3199),
.SN(net2188),
.CK(clk),
.Q(net10287),
.QN(net10286)
);

SDFFS_X2 merge9534(
.D(net335),
.SE(net326),
.SI(net3953),
.SN(net3964),
.CK(clk),
.Q(net10289),
.QN(net10288)
);

SDFFR_X1 merge9535(
.D(net5206),
.RN(net8069),
.SE(net8054),
.SI(net11035),
.CK(clk),
.Q(net10291),
.QN(net10290)
);

OR4_X2 merge9536(
.A1(net5525),
.A2(net5583),
.A3(net482),
.A4(net863),
.ZN(net10292)
);

SDFFR_X2 merge9537(
.D(net6221),
.RN(net6247),
.SE(net5269),
.SI(net4341),
.CK(clk),
.Q(net10294),
.QN(net10293)
);

SDFFS_X1 merge9538(
.D(net3126),
.SE(net3144),
.SI(net2685),
.SN(net1768),
.CK(clk),
.Q(net10296),
.QN(net10295)
);

AOI211_X1 merge9539(
.A(net5328),
.B(net5190),
.C1(net4413),
.C2(net3532),
.ZN(net10297)
);

SDFFS_X2 merge9540(
.D(net2434),
.SE(net2536),
.SI(net6456),
.SN(net6461),
.CK(clk),
.Q(net10299),
.QN(net10298)
);

SDFFR_X1 merge9541(
.D(net867),
.RN(net4716),
.SE(net5375),
.SI(net5399),
.CK(clk),
.Q(net10301),
.QN(net10300)
);

SDFFR_X2 merge9542(
.D(net3364),
.RN(net4205),
.SE(net7176),
.SI(net6179),
.CK(clk),
.Q(net10303),
.QN(net10302)
);

SDFFS_X1 merge9543(
.D(net3306),
.SE(net4395),
.SI(net1687),
.SN(net1691),
.CK(clk),
.Q(net10305),
.QN(net10304)
);

NAND4_X2 merge9544(
.A1(net1660),
.A2(net1647),
.A3(net7236),
.A4(net10483),
.ZN(net10306)
);

SDFFS_X2 merge9545(
.D(net7799),
.SE(net7816),
.SI(net225),
.SN(net214),
.CK(clk),
.Q(net10308),
.QN(net10307)
);

OR4_X4 merge9546(
.A1(net7202),
.A2(net7204),
.A3(net8150),
.A4(net6212),
.ZN(net10309)
);

SDFFR_X1 merge9547(
.D(net6116),
.RN(net8268),
.SE(net6288),
.SI(net6098),
.CK(clk),
.Q(net10311),
.QN(net10310)
);

SDFFR_X2 merge9548(
.D(net8110),
.RN(net9016),
.SE(net3373),
.SI(net4237),
.CK(clk),
.Q(net10313),
.QN(net10312)
);

OAI22_X2 merge9549(
.A1(net2598),
.A2(net2689),
.B1(net574),
.B2(net568),
.ZN(net10314)
);

SDFFS_X1 merge9550(
.D(net5849),
.SE(net1988),
.SI(net4100),
.SN(net11052),
.CK(clk),
.Q(net10316),
.QN(net10315)
);

SDFFS_X2 merge9551(
.D(net3610),
.SE(net2553),
.SI(net4105),
.SN(net4103),
.CK(clk),
.Q(net10318),
.QN(net10317)
);

SDFFR_X1 merge9552(
.D(net6134),
.RN(net6071),
.SE(net7094),
.SI(net7081),
.CK(clk),
.Q(net10320),
.QN(net10319)
);

OAI211_X4 merge9553(
.A(net4120),
.B(net4042),
.C1(net3934),
.C2(net3925),
.ZN(net10321)
);

OAI211_X1 merge9554(
.A(net202),
.B(net182),
.C1(net3249),
.C2(net4100),
.ZN(net10322)
);

SDFFR_X2 merge9555(
.D(net6051),
.RN(net5068),
.SE(net3616),
.SI(net3658),
.CK(clk),
.Q(net10324),
.QN(net10323)
);

NOR4_X4 merge9556(
.A1(net6003),
.A2(net5966),
.A3(net7720),
.A4(net7758),
.ZN(net10325)
);

NOR4_X2 merge9557(
.A1(net4048),
.A2(net4052),
.A3(net224),
.A4(net208),
.ZN(net10326)
);

SDFFS_X1 merge9558(
.D(net5903),
.SE(net6828),
.SI(net6070),
.SN(net6103),
.CK(clk),
.Q(net10328),
.QN(net10327)
);

SDFFS_X2 merge9559(
.D(net1787),
.SE(net2685),
.SI(net7469),
.SN(net7437),
.CK(clk),
.Q(net10330),
.QN(net10329)
);

AOI211_X4 merge9560(
.A(net5233),
.B(net5182),
.C1(net5238),
.C2(net10753),
.ZN(net10331)
);

NOR4_X1 merge9561(
.A1(net1719),
.A2(net1794),
.A3(net3636),
.A4(net2569),
.ZN(net10332)
);

SDFFR_X1 merge9562(
.D(net7715),
.RN(net7817),
.SE(net8762),
.SI(net7724),
.CK(clk),
.Q(net10334),
.QN(net10333)
);

SDFFR_X2 merge9563(
.D(net3391),
.RN(net3348),
.SE(net5012),
.SI(net5027),
.CK(clk),
.Q(net10336),
.QN(net10335)
);

SDFFS_X1 merge9564(
.D(net2589),
.SE(net2673),
.SI(net5082),
.SN(net10607),
.CK(clk),
.Q(net10338),
.QN(net10337)
);

AOI211_X2 merge9565(
.A(net1274),
.B(net2224),
.C1(net2993),
.C2(net6860),
.ZN(net10339)
);

SDFFS_X2 merge9566(
.D(net3121),
.SE(net4150),
.SI(net3960),
.SN(net2993),
.CK(clk),
.Q(net10341),
.QN(net10340)
);

SDFFR_X1 merge9567(
.D(net482),
.RN(net1467),
.SE(net3422),
.SI(net10827),
.CK(clk),
.Q(net10343),
.QN(net10342)
);

SDFFR_X2 merge9568(
.D(net509),
.RN(net482),
.SE(net5014),
.SI(net5008),
.CK(clk),
.Q(net10345),
.QN(net10344)
);

SDFFS_X1 merge9569(
.D(net6193),
.SE(net7136),
.SI(net2152),
.SN(net2144),
.CK(clk),
.Q(net10347),
.QN(net10346)
);

SDFFS_X2 merge9570(
.D(net6987),
.SE(net7260),
.SI(net5321),
.SN(net6428),
.CK(clk),
.Q(net10349),
.QN(net10348)
);

AOI22_X1 merge9571(
.A1(net3597),
.A2(net2696),
.B1(net3712),
.B2(net3705),
.ZN(net10350)
);

AND4_X4 merge9572(
.A1(net4330),
.A2(net3334),
.A3(net2093),
.A4(net2914),
.ZN(net10351)
);

SDFFR_X1 merge9573(
.D(net3921),
.RN(net4034),
.SE(net3117),
.SI(net4075),
.CK(clk),
.Q(net10353),
.QN(net10352)
);

NAND4_X1 merge9574(
.A1(net226),
.A2(net1116),
.A3(net2222),
.A4(net3199),
.ZN(net10354)
);

SDFFR_X2 merge9575(
.D(net3659),
.RN(net2664),
.SE(net2382),
.SI(net10874),
.CK(clk),
.Q(net10356),
.QN(net10355)
);

OR4_X1 merge9576(
.A1(net4562),
.A2(net2732),
.A3(net8048),
.A4(net7847),
.ZN(net10357)
);

OAI22_X1 merge9577(
.A1(net2051),
.A2(net2094),
.B1(net5959),
.B2(net5951),
.ZN(net10358)
);

SDFFS_X1 merge9578(
.D(net3136),
.SE(net2943),
.SI(net2959),
.SN(net5086),
.CK(clk),
.Q(net10360),
.QN(net10359)
);

SDFFS_X2 merge9579(
.D(net1320),
.SE(net1378),
.SI(net6337),
.SN(net7445),
.CK(clk),
.Q(net10362),
.QN(net10361)
);

SDFFR_X1 merge9580(
.D(net8328),
.RN(net8249),
.SE(net2733),
.SI(net5515),
.CK(clk),
.Q(net10364),
.QN(net10363)
);

AND4_X2 merge9581(
.A1(net6386),
.A2(net6381),
.A3(net9067),
.A4(net8111),
.ZN(net10365)
);

SDFFR_X2 merge9582(
.D(net1691),
.RN(net2547),
.SE(net2549),
.SI(net10995),
.CK(clk),
.Q(net10367),
.QN(net10366)
);

AND4_X1 merge9583(
.A1(net1159),
.A2(net1146),
.A3(net2461),
.A4(net1521),
.ZN(net10368)
);

SDFFS_X1 merge9584(
.D(net6547),
.SE(net6546),
.SI(net5158),
.SN(net33),
.CK(clk),
.Q(net10370),
.QN(net10369)
);

SDFFS_X2 merge9585(
.D(net7082),
.SE(net7081),
.SI(net9009),
.SN(net8760),
.CK(clk),
.Q(net10372),
.QN(net10371)
);

SDFFR_X1 merge9586(
.D(net5858),
.RN(net2993),
.SE(net3969),
.SI(net3922),
.CK(clk),
.Q(net10374),
.QN(net10373)
);

SDFFR_X2 merge9587(
.D(net4903),
.RN(net5877),
.SE(net3946),
.SI(net6783),
.CK(clk),
.Q(net10376),
.QN(net10375)
);

NOR2_X1 merge9588(
.A1(net3318),
.A2(net3336),
.ZN(net10377)
);

CLKGATETST_X1 merge9589(
.E(net3519),
.SE(net3533),
.CK(clk),
.GCK(net10378)
);

OR2_X2 merge9590(
.A1(net1379),
.A2(net1412),
.ZN(net10379)
);

CLKGATETST_X2 merge9591(
.E(net419),
.SE(net445),
.CK(clk),
.GCK(net10380)
);

CLKGATETST_X4 merge9592(
.E(net7648),
.SE(net7684),
.CK(clk),
.GCK(net10381)
);

CLKGATETST_X8 merge9593(
.E(net8594),
.SE(net8641),
.CK(clk),
.GCK(net10382)
);

DFFR_X1 merge9594(
.D(net9277),
.RN(net9266),
.CK(clk),
.Q(net10384),
.QN(net10383)
);

DFFR_X2 merge9595(
.D(net8087),
.RN(net8120),
.CK(clk),
.Q(net10386),
.QN(net10385)
);

DFFS_X1 merge9596(
.D(net5607),
.SN(net5653),
.CK(clk),
.Q(net10388),
.QN(net10387)
);

DFFS_X2 merge9597(
.D(net7820),
.SN(net7824),
.CK(clk),
.Q(net10390),
.QN(net10389)
);

NOR2_X4 merge9598(
.A1(net1680),
.A2(net1692),
.ZN(net10391)
);

CLKGATETST_X1 merge9599(
.E(net2537),
.SE(net2552),
.CK(clk),
.GCK(net10392)
);

NOR2_X2 merge9600(
.A1(net4289),
.A2(net4290),
.ZN(net10393)
);

XOR2_X2 merge9601(
.A(net8244),
.B(net8308),
.Z(net10394)
);

CLKGATETST_X2 merge9602(
.E(net3660),
.SE(net3719),
.CK(clk),
.GCK(net10395)
);

CLKGATETST_X4 merge9603(
.E(net312),
.GCK(net319),
.CK(clk)
);

CLKGATETST_X8 merge9604(
.E(net1905),
.SE(net1919),
.CK(clk),
.GCK(net10397)
);

DFFR_X1 merge9605(
.D(net60),
.RN(net91),
.CK(clk),
.Q(net10399),
.QN(net10398)
);

DFFR_X2 merge9606(
.D(net2795),
.RN(net2854),
.CK(clk),
.Q(net10401),
.QN(net10400)
);

DFFS_X1 merge9607(
.D(net1209),
.SN(net1216),
.CK(clk),
.Q(net10403),
.QN(net10402)
);

XNOR2_X1 merge9608(
.A(net726),
.B(net753),
.ZN(net10404)
);

DFFS_X2 merge9609(
.D(net9099),
.SN(net9185),
.CK(clk),
.Q(net10406),
.QN(net10405)
);

OR2_X4 merge9610(
.A1(net8522),
.A2(net8558),
.ZN(net10407)
);

CLKGATETST_X1 merge9611(
.E(net5443),
.SE(net5455),
.CK(clk),
.GCK(net10408)
);

CLKGATETST_X2 merge9612(
.E(net838),
.SE(net795),
.CK(clk),
.GCK(net10409)
);

CLKGATETST_X4 merge9613(
.E(net7719),
.SE(net7711),
.CK(clk),
.GCK(net10410)
);

CLKGATETST_X8 merge9614(
.E(net8721),
.GCK(net8725),
.CK(clk)
);

DFFR_X1 merge9615(
.D(net6798),
.RN(net9832),
.CK(clk),
.Q(net10413),
.QN(net10412)
);

DFFR_X2 merge9616(
.D(net9093),
.RN(net9074),
.CK(clk),
.Q(net10415),
.QN(net10414)
);

DFFS_X1 merge9617(
.D(net8405),
.SN(net8479),
.CK(clk),
.Q(net10417),
.QN(net10416)
);

DFFS_X2 merge9618(
.D(net5013),
.SN(net5020),
.CK(clk),
.Q(net10419),
.QN(net10418)
);

OR2_X1 merge9619(
.A1(net4364),
.A2(net4433),
.ZN(net10420)
);

CLKGATETST_X1 merge9620(
.E(net5821),
.SE(net5830),
.CK(clk),
.GCK(net10421)
);

CLKGATETST_X2 merge9621(
.E(net855),
.SE(net896),
.CK(clk),
.GCK(net10422)
);

CLKGATETST_X4 merge9622(
.E(net7906),
.SE(net7912),
.CK(clk),
.GCK(net10423)
);

XNOR2_X2 merge9623(
.A(net1882),
.B(net1808),
.ZN(net10424)
);

AND2_X4 merge9624(
.A1(net641),
.A2(net664),
.ZN(net10425)
);

CLKGATETST_X8 merge9625(
.E(net5176),
.SE(net5179),
.CK(clk),
.GCK(net10426)
);

DFFR_X1 merge9626(
.D(net7436),
.RN(net7466),
.CK(clk),
.Q(net10428),
.QN(net10427)
);

DFFR_X2 merge9627(
.D(net5367),
.RN(net5387),
.CK(clk),
.Q(net10430),
.QN(net10429)
);

AND2_X1 merge9628(
.A1(net9364),
.A2(net9362),
.ZN(net10431)
);

NAND2_X1 merge9629(
.A1(net2081),
.A2(net2084),
.ZN(net10432)
);

DFFS_X1 merge9630(
.D(net6917),
.SN(net6946),
.CK(clk),
.Q(net10434),
.QN(net10433)
);

NAND2_X2 merge9631(
.A1(net7002),
.A2(net7074),
.ZN(net10435)
);

DFFS_X2 merge9632(
.D(net5860),
.SN(net5936),
.CK(clk),
.Q(net10437),
.QN(net10436)
);

CLKGATETST_X1 merge9633(
.E(net6311),
.SE(net6374),
.CK(clk),
.GCK(net10438)
);

CLKGATETST_X2 merge9634(
.E(net2605),
.SE(net2608),
.CK(clk),
.GCK(net10439)
);

NAND2_X4 merge9635(
.A1(net3430),
.A2(net3433),
.ZN(net10440)
);

CLKGATETST_X4 merge9636(
.E(net388),
.SE(net389),
.CK(clk),
.GCK(net10441)
);

CLKGATETST_X8 merge9637(
.E(net9589),
.SE(net9833),
.CK(clk),
.GCK(net10442)
);

DFFR_X1 merge9638(
.D(net1796),
.RN(net1748),
.CK(clk),
.Q(net10444),
.QN(net10443)
);

DFFR_X2 merge9639(
.D(net4967),
.RN(net4935),
.CK(clk),
.Q(net10446),
.QN(net10445)
);

DFFS_X1 merge9640(
.D(net4737),
.SN(net4772),
.CK(clk),
.Q(net10448),
.QN(net10447)
);

DFFS_X2 merge9641(
.D(net8358),
.SN(net8354),
.CK(clk),
.Q(net10450),
.QN(net10449)
);

CLKGATETST_X1 merge9642(
.E(net9377),
.SE(net9461),
.CK(clk),
.GCK(net10451)
);

CLKGATETST_X2 merge9643(
.E(net9463),
.SE(net9538),
.CK(clk),
.GCK(net10452)
);

CLKGATETST_X4 merge9644(
.E(net8201),
.SE(net8222),
.CK(clk),
.GCK(net10453)
);

CLKGATETST_X8 merge9645(
.E(net6208),
.SE(net6244),
.CK(clk),
.GCK(net10454)
);

AND2_X2 merge9646(
.A1(net3613),
.A2(net3634),
.ZN(net10455)
);

XOR2_X1 merge9647(
.A(net1461),
.B(net1519),
.Z(net10456)
);

DFFR_X1 merge9648(
.D(net3040),
.RN(net3086),
.CK(clk),
.Q(net10458),
.QN(net10457)
);

NOR2_X1 merge9649(
.A1(net6153),
.A2(net6175),
.ZN(net10459)
);

OR2_X2 merge9650(
.A1(net4114),
.A2(net4119),
.ZN(net10460)
);

DFFR_X2 merge9651(
.D(net4530),
.RN(net4605),
.CK(clk),
.Q(net10462),
.QN(net10461)
);

DFFS_X1 merge9652(
.D(net4660),
.SN(net4661),
.CK(clk),
.Q(net10464),
.QN(net10463)
);

DFFS_X2 merge9653(
.D(net6832),
.SN(net6845),
.CK(clk),
.Q(net10466),
.QN(net10465)
);

NOR2_X4 merge9654(
.A1(net6497),
.A2(net6521),
.ZN(net10467)
);

NOR2_X2 merge9655(
.A1(net8023),
.A2(net8029),
.ZN(net10468)
);

XOR2_X2 merge9656(
.A(net2723),
.B(net2739),
.Z(net10469)
);

CLKGATETST_X1 merge9657(
.E(net2040),
.SE(net2067),
.CK(clk),
.GCK(net10470)
);

XNOR2_X1 merge9658(
.A(net5088),
.B(net5094),
.ZN(net10471)
);

CLKGATETST_X2 merge9659(
.E(net1001),
.SE(net1002),
.CK(clk),
.GCK(net10472)
);

CLKGATETST_X4 merge9660(
.E(net8930),
.SE(net8997),
.CK(clk),
.GCK(net10473)
);

CLKGATETST_X8 merge9661(
.E(net8829),
.SE(net8895),
.CK(clk),
.GCK(net10474)
);

DFFR_X1 merge9662(
.D(net5678),
.RN(net5690),
.CK(clk),
.Q(net10476),
.QN(net10475)
);

DFFR_X2 merge9663(
.D(net6579),
.RN(net6591),
.CK(clk),
.Q(net10478),
.QN(net10477)
);

DFFS_X1 merge9664(
.D(net4188),
.SN(net4195),
.CK(clk),
.Q(net10480),
.QN(net10479)
);

DFFS_X2 merge9665(
.D(net5499),
.SN(net5520),
.CK(clk),
.Q(net10482),
.QN(net10481)
);

CLKGATETST_X1 merge9666(
.E(net7190),
.SE(net7217),
.CK(clk),
.GCK(net10483)
);

CLKGATETST_X2 merge9667(
.E(net210),
.SE(net215),
.CK(clk),
.GCK(net10484)
);

CLKGATETST_X4 merge9668(
.E(net3833),
.SE(net3837),
.CK(clk),
.GCK(net10485)
);

OR2_X4 merge9669(
.A1(net6076),
.A2(net6095),
.ZN(net10486)
);

OR2_X1 merge9670(
.A1(net7281),
.A2(net7280),
.ZN(net10487)
);

XNOR2_X2 merge9671(
.A(net1588),
.B(net1594),
.ZN(net10488)
);

CLKGATETST_X8 merge9672(
.E(net2950),
.SE(net2905),
.CK(clk),
.GCK(net10489)
);

AND2_X4 merge9673(
.A1(net7341),
.A2(net7349),
.ZN(net10490)
);

DFFR_X1 merge9674(
.D(net6007),
.RN(net6012),
.CK(clk),
.Q(net10492),
.QN(net10491)
);

DFFR_X2 merge9675(
.D(net7555),
.RN(net7557),
.CK(clk),
.Q(net10494),
.QN(net10493)
);

AND2_X1 merge9676(
.A1(net3225),
.A2(net3302),
.ZN(net10495)
);

DFFS_X1 merge9677(
.D(net6398),
.SN(net6446),
.CK(clk),
.Q(net10497),
.QN(net10496)
);

NAND2_X1 merge9678(
.A1(net2161),
.A2(net2196),
.ZN(net10498)
);

NAND2_X2 merge9679(
.A1(net4060),
.A2(net4017),
.ZN(net10499)
);

DFFS_X2 merge9680(
.D(net2973),
.SN(net2988),
.CK(clk),
.Q(net10501),
.QN(net10500)
);

CLKGATETST_X1 merge9681(
.E(net2350),
.SE(net2338),
.CK(clk),
.GCK(net10502)
);

CLKGATETST_X2 merge9682(
.E(net4857),
.SE(net4863),
.CK(clk),
.GCK(net10503)
);

NAND2_X4 merge9683(
.A1(net1180),
.A2(net1182),
.ZN(net10504)
);

CLKGATETST_X4 merge9684(
.E(net3928),
.SE(net3948),
.CK(clk),
.GCK(net10505)
);

AND2_X2 merge9685(
.A1(net1019),
.A2(net1098),
.ZN(net10506)
);

CLKGATETST_X8 merge9686(
.E(net7091),
.SE(net7135),
.CK(clk),
.GCK(net10507)
);

XOR2_X1 merge9687(
.A(net3149),
.B(net3138),
.Z(net10508)
);

DFFR_X1 merge9688(
.D(net3738),
.RN(net3734),
.CK(clk),
.Q(net10510),
.QN(net10509)
);

NOR2_X1 merge9689(
.A1(net5256),
.A2(net5317),
.ZN(net10511)
);

DFFR_X2 merge9690(
.D(net4439),
.RN(net4464),
.CK(clk),
.Q(net10513),
.QN(net10512)
);

DFFS_X1 merge9691(
.D(net6686),
.SN(net6713),
.CK(clk),
.Q(net10515),
.QN(net10514)
);

DFFS_X2 merge9692(
.D(net8756),
.SN(net8816),
.CK(clk),
.Q(net10517),
.QN(net10516)
);

CLKGATETST_X1 merge9693(
.E(net536),
.SE(net539),
.CK(clk),
.GCK(net10518)
);

OR2_X2 merge9694(
.A1(net1318),
.A2(net1328),
.ZN(net10519)
);

NOR2_X4 merge9695(
.A1(net2269),
.A2(net2286),
.ZN(net10520)
);

CLKGATETST_X2 merge9696(
.E(net3980),
.SE(net3104),
.CK(clk),
.GCK(net10521)
);

NOR2_X2 merge9697(
.A1(net4417),
.A2(net3355),
.ZN(net10522)
);

CLKGATETST_X4 merge9698(
.E(net9486),
.SE(net9530),
.CK(clk),
.GCK(net10523)
);

CLKGATETST_X8 merge9699(
.E(net1982),
.SE(net1082),
.CK(clk),
.GCK(net10524)
);

DFFR_X1 merge9700(
.D(net4165),
.RN(net3994),
.CK(clk),
.Q(net10526),
.QN(net10525)
);

DFFR_X2 merge9701(
.D(net1183),
.RN(net10200),
.CK(clk),
.Q(net10528),
.QN(net10527)
);

DFFS_X1 merge9702(
.D(net1621),
.SN(net1614),
.CK(clk),
.Q(net10530),
.QN(net10529)
);

DFFS_X2 merge9703(
.D(net1947),
.SN(net1976),
.CK(clk),
.Q(net10532),
.QN(net10531)
);

XOR2_X2 merge9704(
.A(net2595),
.B(net1513),
.Z(net10533)
);

XNOR2_X1 merge9705(
.A(net3703),
.B(net2760),
.ZN(net10534)
);

OR2_X4 merge9706(
.A1(net1487),
.A2(net1539),
.ZN(net10535)
);

CLKGATETST_X1 merge9707(
.E(net1013),
.SE(net10506),
.CK(clk),
.GCK(net10536)
);

OR2_X1 merge9708(
.A1(net3212),
.A2(net2230),
.ZN(net10537)
);

CLKGATETST_X2 merge9709(
.E(net4696),
.SE(net4774),
.CK(clk),
.GCK(net10538)
);

XNOR2_X2 merge9710(
.A(net3366),
.B(net3157),
.ZN(net10539)
);

CLKGATETST_X4 merge9711(
.E(net1928),
.SE(net3034),
.CK(clk),
.GCK(net10540)
);

CLKGATETST_X8 merge9712(
.E(net8503),
.SE(net8525),
.CK(clk),
.GCK(net10541)
);

DFFR_X1 merge9713(
.D(net3839),
.RN(net3996),
.CK(clk),
.Q(net10543),
.QN(net10542)
);

DFFR_X2 merge9714(
.D(net8298),
.RN(net8400),
.CK(clk),
.Q(net10545),
.QN(net10544)
);

DFFS_X1 merge9715(
.D(net9501),
.SN(net8614),
.CK(clk),
.Q(net10546),
.QN(out4)
);

DFFS_X2 merge9716(
.D(net7393),
.SN(net7242),
.CK(clk),
.Q(net10548),
.QN(net10547)
);

CLKGATETST_X1 merge9717(
.E(net8377),
.SE(net8459),
.CK(clk),
.GCK(net10549)
);

CLKGATETST_X2 merge9718(
.E(net7634),
.SE(net8499),
.CK(clk),
.GCK(net10550)
);

CLKGATETST_X4 merge9719(
.E(net3470),
.SE(net3360),
.CK(clk),
.GCK(net10551)
);

CLKGATETST_X8 merge9720(
.E(net3398),
.SE(net2416),
.CK(clk),
.GCK(net10552)
);

AND2_X4 merge9721(
.A1(net4156),
.A2(net2207),
.ZN(net10553)
);

DFFR_X1 merge9722(
.D(net5867),
.RN(net6889),
.CK(clk),
.Q(net10555),
.QN(net10554)
);

AND2_X1 merge9723(
.A1(net7013),
.A2(net7075),
.ZN(net10556)
);

NAND2_X1 merge9724(
.A1(net2226),
.A2(net3160),
.ZN(net10557)
);

DFFR_X2 merge9725(
.D(net7070),
.RN(net7032),
.CK(clk),
.Q(net10559),
.QN(net10558)
);

NAND2_X2 merge9726(
.A1(net2331),
.A2(net3465),
.ZN(net10560)
);

NAND2_X4 merge9727(
.A1(net3915),
.A2(net4962),
.ZN(net10561)
);

DFFS_X1 merge9728(
.D(net3816),
.SN(net4714),
.CK(clk),
.Q(net10563),
.QN(net10562)
);

DFFS_X2 merge9729(
.D(net7595),
.SN(net7624),
.CK(clk),
.Q(net10565),
.QN(net10564)
);

CLKGATETST_X1 merge9730(
.E(net8063),
.SE(net8969),
.CK(clk),
.GCK(net10566)
);

CLKGATETST_X2 merge9731(
.E(net5291),
.SE(net4504),
.CK(clk),
.GCK(net10567)
);

CLKGATETST_X4 merge9732(
.E(net5908),
.SE(net7787),
.CK(clk),
.GCK(net10568)
);

CLKGATETST_X8 merge9733(
.E(net5130),
.SE(net4244),
.CK(clk),
.GCK(net10569)
);

DFFR_X1 merge9734(
.D(net8125),
.RN(net7144),
.CK(clk),
.Q(net10571),
.QN(net10570)
);

DFFR_X2 merge9735(
.D(net6720),
.RN(net5656),
.CK(clk),
.Q(net10573),
.QN(net10572)
);

AND2_X2 merge9736(
.A1(net7322),
.A2(net8253),
.ZN(net10574)
);

XOR2_X1 merge9737(
.A(net2118),
.B(net1272),
.Z(net10575)
);

DFFS_X1 merge9738(
.D(net1860),
.SN(net1874),
.CK(clk),
.Q(net10577),
.QN(net10576)
);

DFFS_X2 merge9739(
.D(net463),
.SN(net1452),
.CK(clk),
.Q(net10579),
.QN(net10578)
);

NOR2_X1 merge9740(
.A1(net2384),
.A2(net2251),
.ZN(net10580)
);

CLKGATETST_X1 merge9741(
.E(net8849),
.SE(net7943),
.CK(clk),
.GCK(net10581)
);

CLKGATETST_X2 merge9742(
.E(net3982),
.SE(net3959),
.CK(clk),
.GCK(net10582)
);

CLKGATETST_X4 merge9743(
.E(net9202),
.SE(net9279),
.CK(clk),
.GCK(net10583)
);

CLKGATETST_X8 merge9744(
.E(net5213),
.SE(net3286),
.CK(clk),
.GCK(net10584)
);

DFFR_X1 merge9745(
.D(net8040),
.RN(net8814),
.CK(clk),
.Q(net10586),
.QN(net10585)
);

DFFR_X2 merge9746(
.D(net7396),
.RN(net5561),
.CK(clk),
.Q(net10588),
.QN(net10587)
);

DFFS_X1 merge9747(
.D(net1865),
.SN(net925),
.CK(clk),
.Q(net10590),
.QN(net10589)
);

OR2_X2 merge9748(
.A1(net1852),
.A2(net918),
.ZN(net10591)
);

NOR2_X4 merge9749(
.A1(net2291),
.A2(net2330),
.ZN(net10592)
);

DFFS_X2 merge9750(
.D(net4708),
.SN(net6668),
.CK(clk),
.Q(net10594),
.QN(net10593)
);

CLKGATETST_X1 merge9751(
.E(net4513),
.SE(net4537),
.CK(clk),
.GCK(net10595)
);

NOR2_X2 merge9752(
.A1(net1267),
.A2(net2127),
.ZN(net10596)
);

XOR2_X2 merge9753(
.A(net2637),
.B(net2679),
.Z(net10597)
);

XNOR2_X1 merge9754(
.A(net8389),
.B(net6626),
.ZN(net10598)
);

OR2_X4 merge9755(
.A1(net1491),
.A2(net1439),
.ZN(net10599)
);

CLKGATETST_X2 merge9756(
.E(net8815),
.SE(net6901),
.CK(clk),
.GCK(net10600)
);

CLKGATETST_X4 merge9757(
.E(net2805),
.SE(net2845),
.CK(clk),
.GCK(net10601)
);

CLKGATETST_X8 merge9758(
.E(net6285),
.SE(net6334),
.CK(clk),
.GCK(net10602)
);

OR2_X1 merge9759(
.A1(net2128),
.A2(net1361),
.ZN(net10603)
);

XNOR2_X2 merge9760(
.A(net7513),
.B(net7410),
.ZN(net10604)
);

DFFR_X1 merge9761(
.D(net3752),
.RN(net4584),
.CK(clk),
.Q(net10606),
.QN(net10605)
);

DFFR_X2 merge9762(
.D(net4130),
.RN(net4170),
.CK(clk),
.Q(net10608),
.QN(net10607)
);

DFFS_X1 merge9763(
.D(net4940),
.SN(net4085),
.CK(clk),
.Q(net10610),
.QN(net10609)
);

AND2_X4 merge9764(
.A1(net4470),
.A2(net6296),
.ZN(net10611)
);

AND2_X1 merge9765(
.A1(net5280),
.A2(net5111),
.ZN(net10612)
);

NAND2_X1 merge9766(
.A1(net4590),
.A2(net2630),
.ZN(net10613)
);

DFFS_X2 merge9767(
.D(net6362),
.SN(net5308),
.CK(clk),
.Q(net10615),
.QN(net10614)
);

CLKGATETST_X1 merge9768(
.E(net924),
.SE(net1881),
.CK(clk),
.GCK(net10616)
);

CLKGATETST_X2 merge9769(
.E(net2591),
.SE(net3466),
.CK(clk),
.GCK(net10617)
);

CLKGATETST_X4 merge9770(
.E(net8544),
.SE(net8521),
.CK(clk),
.GCK(net10618)
);

CLKGATETST_X8 merge9771(
.E(net4791),
.SE(net6523),
.CK(clk),
.GCK(net10619)
);

NAND2_X2 merge9772(
.A1(net6246),
.A2(net7028),
.ZN(net10620)
);

DFFR_X1 merge9773(
.D(net8728),
.RN(net8810),
.CK(clk),
.Q(net10622),
.QN(net10621)
);

DFFR_X2 merge9774(
.D(net6851),
.RN(net7879),
.CK(clk),
.Q(net10624),
.QN(net10623)
);

DFFS_X1 merge9775(
.D(net9246),
.SN(net8404),
.CK(clk),
.Q(net10626),
.QN(net10625)
);

NAND2_X4 merge9776(
.A1(net8227),
.A2(net9054),
.ZN(net10627)
);

DFFS_X2 merge9777(
.D(net2136),
.SN(net3023),
.CK(clk),
.Q(net10629),
.QN(net10628)
);

AND2_X2 merge9778(
.A1(net4480),
.A2(net5571),
.ZN(net10630)
);

CLKGATETST_X1 merge9779(
.E(net6610),
.SE(net6379),
.CK(clk),
.GCK(net10631)
);

XOR2_X1 merge9780(
.A(net4558),
.B(net2660),
.Z(net10632)
);

CLKGATETST_X2 merge9781(
.E(net1249),
.SE(net9890),
.CK(clk),
.GCK(net10633)
);

CLKGATETST_X4 merge9782(
.E(net7026),
.SE(net6111),
.CK(clk),
.GCK(net10634)
);

CLKGATETST_X8 merge9783(
.E(net6857),
.SE(net4944),
.CK(clk),
.GCK(net10635)
);

DFFR_X1 merge9784(
.D(net398),
.RN(net9740),
.CK(clk),
.Q(net10637),
.QN(net10636)
);

NOR2_X1 merge9785(
.A1(net3163),
.A2(net3207),
.ZN(net10638)
);

DFFR_X2 merge9786(
.D(net6893),
.RN(net8809),
.CK(clk),
.Q(net10640),
.QN(net10639)
);

DFFS_X1 merge9787(
.D(net6724),
.SN(net7570),
.CK(clk),
.Q(net10642),
.QN(net10641)
);

DFFS_X2 merge9788(
.D(net1421),
.SN(net1347),
.CK(clk),
.Q(net10644),
.QN(net10643)
);

OR2_X2 merge9789(
.A1(net7249),
.A2(net9082),
.ZN(net10645)
);

NOR2_X4 merge9790(
.A1(net8904),
.A2(net9030),
.ZN(net10646)
);

CLKGATETST_X1 merge9791(
.E(net5475),
.SE(net6330),
.CK(clk),
.GCK(net10647)
);

CLKGATETST_X2 merge9792(
.E(net4735),
.SE(net5695),
.CK(clk),
.GCK(net10648)
);

NOR2_X2 merge9793(
.A1(net9068),
.A2(net7219),
.ZN(net10649)
);

XOR2_X2 merge9794(
.A(net1489),
.B(net1517),
.Z(net10650)
);

XNOR2_X1 merge9795(
.A(net5132),
.B(net4166),
.ZN(net10651)
);

OR2_X4 merge9796(
.A1(net6280),
.A2(net5183),
.ZN(net10652)
);

CLKGATETST_X4 merge9797(
.E(net7006),
.SE(net7934),
.CK(clk),
.GCK(net10653)
);

CLKGATETST_X8 merge9798(
.E(net3714),
.SE(net2675),
.CK(clk),
.GCK(net10654)
);

DFFR_X1 merge9799(
.D(net8527),
.RN(net8571),
.CK(clk),
.Q(net10656),
.QN(net10655)
);

DFFR_X2 merge9800(
.D(net2201),
.RN(net2417),
.CK(clk),
.Q(net10658),
.QN(net10657)
);

DFFS_X1 merge9801(
.D(net5032),
.SN(net7041),
.CK(clk),
.Q(net10660),
.QN(net10659)
);

OR2_X1 merge9802(
.A1(net5021),
.A2(net6195),
.ZN(net10661)
);

DFFS_X2 merge9803(
.D(net9350),
.SN(net7591),
.CK(clk),
.Q(net10663),
.QN(net10662)
);

XNOR2_X2 merge9804(
.A(net8138),
.B(net8043),
.ZN(net10664)
);

CLKGATETST_X1 merge9805(
.E(net1964),
.SE(net2004),
.CK(clk),
.GCK(net10665)
);

AND2_X4 merge9806(
.A1(net7959),
.A2(net6972),
.ZN(net10666)
);

CLKGATETST_X2 merge9807(
.E(net9133),
.SE(net9151),
.CK(clk),
.GCK(net10667)
);

CLKGATETST_X4 merge9808(
.E(net9459),
.SE(net6666),
.CK(clk),
.GCK(net10668)
);

AND2_X1 merge9809(
.A1(net5105),
.A2(net4408),
.ZN(net10669)
);

CLKGATETST_X8 merge9810(
.E(net2362),
.SE(net1595),
.CK(clk),
.GCK(net10670)
);

DFFR_X1 merge9811(
.D(net4501),
.RN(net3555),
.CK(clk),
.Q(net10672),
.QN(net10671)
);

DFFR_X2 merge9812(
.D(net1849),
.RN(net3808),
.CK(clk),
.Q(net10674),
.QN(net10673)
);

DFFS_X1 merge9813(
.D(net3901),
.SN(net3900),
.CK(clk),
.Q(net10676),
.QN(net10675)
);

DFFS_X2 merge9814(
.D(net2830),
.SN(net4761),
.CK(clk),
.Q(net10678),
.QN(net10677)
);

CLKGATETST_X1 merge9815(
.E(net5281),
.SE(net7337),
.CK(clk),
.GCK(net10679)
);

CLKGATETST_X2 merge9816(
.E(net4163),
.SE(net3214),
.CK(clk),
.GCK(net10680)
);

NAND2_X1 merge9817(
.A1(net6015),
.A2(net8836),
.ZN(net10681)
);

CLKGATETST_X4 merge9818(
.E(net5881),
.SE(net5926),
.CK(clk),
.GCK(net10682)
);

CLKGATETST_X8 merge9819(
.E(net7335),
.SE(net8989),
.CK(clk),
.GCK(net10683)
);

DFFR_X1 merge9820(
.D(net9978),
.RN(net10322),
.CK(clk),
.Q(net10685),
.QN(net10684)
);

NAND2_X2 merge9821(
.A1(net6971),
.A2(net6983),
.ZN(net10686)
);

NAND2_X4 merge9822(
.A1(net8870),
.A2(net7942),
.ZN(net10687)
);

DFFR_X2 merge9823(
.D(net8052),
.RN(net7057),
.CK(clk),
.Q(net10689),
.QN(net10688)
);

DFFS_X1 merge9824(
.D(net4325),
.SN(net4164),
.CK(clk),
.Q(net10691),
.QN(net10690)
);

DFFS_X2 merge9825(
.D(net4680),
.SN(net4552),
.CK(clk),
.Q(net10693),
.QN(net10692)
);

CLKGATETST_X1 merge9826(
.E(net4901),
.SE(net5055),
.CK(clk),
.GCK(net10694)
);

CLKGATETST_X2 merge9827(
.E(net5709),
.SE(net3744),
.CK(clk),
.GCK(net10695)
);

AND2_X2 merge9828(
.A1(net5049),
.A2(net5225),
.ZN(net10696)
);

XOR2_X1 merge9829(
.A(net6100),
.B(net5125),
.Z(net10697)
);

NOR2_X1 merge9830(
.A1(net3650),
.A2(net3368),
.ZN(net10698)
);

CLKGATETST_X4 merge9831(
.E(net9225),
.SE(net9057),
.CK(clk),
.GCK(net10699)
);

CLKGATETST_X8 merge9832(
.E(net8050),
.SE(net5122),
.CK(clk),
.GCK(net10700)
);

DFFR_X1 merge9833(
.D(net8554),
.RN(net9408),
.CK(clk),
.Q(net10702),
.QN(net10701)
);

OR2_X2 merge9834(
.A1(net2304),
.A2(net2297),
.ZN(net10703)
);

NOR2_X4 merge9835(
.A1(net9437),
.A2(net9460),
.ZN(net10704)
);

NOR2_X2 merge9836(
.A1(net5483),
.A2(net6274),
.ZN(net10705)
);

DFFR_X2 merge9837(
.D(net7016),
.RN(net7022),
.CK(clk),
.Q(net10707),
.QN(net10706)
);

DFFS_X1 merge9838(
.D(net8305),
.SN(net6443),
.CK(clk),
.Q(net10709),
.QN(net10708)
);

XOR2_X2 merge9839(
.A(net8876),
.B(net8804),
.Z(net10710)
);

DFFS_X2 merge9840(
.D(net5928),
.SN(net6254),
.CK(clk),
.Q(net10712),
.QN(net10711)
);

XNOR2_X1 merge9841(
.A(net8854),
.B(net9069),
.ZN(net10713)
);

CLKGATETST_X1 merge9842(
.E(net8955),
.SE(net9037),
.CK(clk),
.GCK(net10714)
);

OR2_X4 merge9843(
.A1(net5203),
.A2(net4422),
.ZN(net10715)
);

CLKGATETST_X2 merge9844(
.E(net1823),
.SE(net1845),
.CK(clk),
.GCK(net10716)
);

CLKGATETST_X4 merge9845(
.E(net2050),
.SE(net9724),
.CK(clk),
.GCK(net10717)
);

OR2_X1 merge9846(
.A1(net4352),
.A2(net4254),
.ZN(net10718)
);

XNOR2_X2 merge9847(
.A(net9351),
.B(net8577),
.ZN(net10719)
);

CLKGATETST_X8 merge9848(
.E(net8588),
.SE(net4785),
.CK(clk),
.GCK(net10720)
);

DFFR_X1 merge9849(
.D(net6688),
.RN(net6702),
.CK(clk),
.Q(net10722),
.QN(net10721)
);

DFFR_X2 merge9850(
.D(net8395),
.RN(net8475),
.CK(clk),
.Q(net10724),
.QN(net10723)
);

DFFS_X1 merge9851(
.D(net5718),
.SN(net8566),
.CK(clk),
.Q(net10726),
.QN(net10725)
);

DFFS_X2 merge9852(
.D(net406),
.SN(net2235),
.CK(clk),
.Q(net10728),
.QN(net10727)
);

CLKGATETST_X1 merge9853(
.E(net2763),
.SE(net6678),
.CK(clk),
.GCK(net10729)
);

CLKGATETST_X2 merge9854(
.E(net2655),
.SE(net2651),
.CK(clk),
.GCK(net10730)
);

CLKGATETST_X4 merge9855(
.E(net3800),
.SE(net4369),
.CK(clk),
.GCK(net10731)
);

CLKGATETST_X8 merge9856(
.E(net4176),
.SE(net4258),
.CK(clk),
.GCK(net10732)
);

DFFR_X1 merge9857(
.D(net6696),
.RN(net5564),
.CK(clk),
.Q(net10734),
.QN(net10733)
);

DFFR_X2 merge9858(
.D(net7468),
.RN(net9349),
.CK(clk),
.Q(net10736),
.QN(net10735)
);

DFFS_X1 merge9859(
.D(net9310),
.SN(net9162),
.CK(clk),
.Q(net10738),
.QN(net10737)
);

DFFS_X2 merge9860(
.D(net10603),
.SN(net2119),
.CK(clk),
.Q(net10740),
.QN(net10739)
);

AND2_X4 merge9861(
.A1(net7149),
.A2(net7235),
.ZN(net10741)
);

CLKGATETST_X1 merge9862(
.E(net8512),
.SE(net9454),
.CK(clk),
.GCK(net10742)
);

CLKGATETST_X2 merge9863(
.E(net3351),
.SE(net9880),
.CK(clk),
.GCK(net10743)
);

CLKGATETST_X4 merge9864(
.E(net8880),
.SE(net7873),
.CK(clk),
.GCK(net10744)
);

CLKGATETST_X8 merge9865(
.E(net5029),
.SE(net5048),
.CK(clk),
.GCK(net10745)
);

DFFR_X1 merge9866(
.D(net4565),
.RN(net5282),
.CK(clk),
.Q(net10747),
.QN(net10746)
);

DFFR_X2 merge9867(
.D(net5742),
.RN(net4557),
.CK(clk),
.Q(net10749),
.QN(net10748)
);

DFFS_X1 merge9868(
.D(net8982),
.SN(net9036),
.CK(clk),
.Q(net10751),
.QN(net10750)
);

DFFS_X2 merge9869(
.D(net5274),
.SN(net9097),
.CK(clk),
.Q(net10753),
.QN(net10752)
);

CLKGATETST_X1 merge9870(
.E(net6360),
.SE(net7508),
.CK(clk),
.GCK(net10754)
);

CLKGATETST_X2 merge9871(
.E(net9174),
.SE(net9135),
.CK(clk),
.GCK(net10755)
);

CLKGATETST_X4 merge9872(
.E(net4685),
.SE(net6279),
.CK(clk),
.GCK(net10756)
);

CLKGATETST_X8 merge9873(
.E(net3453),
.SE(net3446),
.CK(clk),
.GCK(net10757)
);

DFFR_X1 merge9874(
.D(net6440),
.RN(net6345),
.CK(clk),
.Q(net10759),
.QN(net10758)
);

DFFR_X2 merge9875(
.D(net9450),
.RN(net9375),
.CK(clk),
.Q(net10761),
.QN(net10760)
);

DFFS_X1 merge9876(
.D(net2823),
.SN(net1803),
.CK(clk),
.Q(net10763),
.QN(net10762)
);

DFFS_X2 merge9877(
.D(net7613),
.SN(net6723),
.CK(clk),
.Q(net10765),
.QN(net10764)
);

CLKGATETST_X1 merge9878(
.E(net7611),
.SE(net9497),
.CK(clk),
.GCK(out15)
);

CLKGATETST_X2 merge9879(
.E(net1873),
.SE(net3824),
.CK(clk),
.GCK(net10766)
);

AND2_X1 merge9880(
.A1(net6540),
.A2(net5671),
.ZN(net10767)
);

CLKGATETST_X4 merge9881(
.E(net9462),
.SE(net7687),
.CK(clk),
.GCK(net10768)
);

CLKGATETST_X8 merge9882(
.E(net8507),
.SE(net9465),
.CK(clk),
.GCK(net10769)
);

DFFR_X1 merge9883(
.D(net10211),
.RN(net10358),
.CK(clk),
.Q(net10771),
.QN(net10770)
);

DFFR_X2 merge9884(
.D(net10533),
.RN(net10488),
.CK(clk),
.Q(net10773),
.QN(net10772)
);

DFFS_X1 merge9885(
.D(net9276),
.SN(net8252),
.CK(clk),
.Q(net10775),
.QN(net10774)
);

DFFS_X2 merge9886(
.D(net8971),
.SN(net5915),
.CK(clk),
.Q(net10777),
.QN(net10776)
);

CLKGATETST_X1 merge9887(
.E(net5929),
.SE(net10096),
.CK(clk),
.GCK(net10778)
);

NAND2_X1 merge9888(
.A1(net4521),
.A2(net5268),
.ZN(net10779)
);

CLKGATETST_X2 merge9889(
.E(net7055),
.SE(net7234),
.CK(clk),
.GCK(net10780)
);

CLKGATETST_X4 merge9890(
.E(net10280),
.SE(net474),
.CK(clk),
.GCK(net10781)
);

CLKGATETST_X8 merge9891(
.E(net649),
.SE(net10248),
.CK(clk),
.GCK(net10782)
);

DFFR_X1 merge9892(
.D(net10184),
.RN(net10561),
.CK(clk),
.Q(net10784),
.QN(net10783)
);

DFFR_X2 merge9893(
.D(net6318),
.RN(net6199),
.CK(clk),
.Q(net10786),
.QN(net10785)
);

DFFS_X1 merge9894(
.D(net4751),
.SN(net4745),
.CK(clk),
.Q(net10788),
.QN(net10787)
);

DFFS_X2 merge9895(
.D(net8972),
.SN(net8924),
.CK(clk),
.Q(net10790),
.QN(net10789)
);

CLKGATETST_X1 merge9896(
.E(net8134),
.SE(net8269),
.CK(clk),
.GCK(net10791)
);

NAND2_X2 merge9897(
.A1(net9092),
.A2(net9163),
.ZN(net10792)
);

CLKGATETST_X2 merge9898(
.E(net9884),
.SE(net3642),
.CK(clk),
.GCK(net10793)
);

CLKGATETST_X4 merge9899(
.E(net9012),
.SE(net9080),
.CK(clk),
.GCK(net10794)
);

CLKGATETST_X8 merge9900(
.E(net6701),
.SE(net5751),
.CK(clk),
.GCK(net10795)
);

NAND2_X4 merge9901(
.A1(net9347),
.A2(net9439),
.ZN(net10796)
);

DFFR_X1 merge9902(
.D(net4497),
.RN(net4695),
.CK(clk),
.Q(net10798),
.QN(net10797)
);

DFFR_X2 merge9903(
.D(net10651),
.RN(net10519),
.CK(clk),
.Q(net10800),
.QN(net10799)
);

DFFS_X1 merge9904(
.D(net8937),
.SN(net9003),
.CK(clk),
.Q(net10802),
.QN(net10801)
);

DFFS_X2 merge9905(
.D(net564),
.SN(net9988),
.CK(clk),
.Q(net10804),
.QN(net10803)
);

CLKGATETST_X1 merge9906(
.E(net6604),
.SE(net5663),
.CK(clk),
.GCK(net10805)
);

CLKGATETST_X2 merge9907(
.E(net9876),
.SE(net10432),
.CK(clk),
.GCK(net10806)
);

CLKGATETST_X4 merge9908(
.E(net6885),
.SE(net9924),
.CK(clk),
.GCK(net10807)
);

CLKGATETST_X8 merge9909(
.E(net10004),
.SE(net10194),
.CK(clk),
.GCK(net10808)
);

DFFR_X1 merge9910(
.D(net10368),
.RN(net285),
.CK(clk),
.Q(net10810),
.QN(net10809)
);

DFFR_X2 merge9911(
.D(net10321),
.RN(net10124),
.CK(clk),
.Q(net10812),
.QN(net10811)
);

DFFS_X1 merge9912(
.D(net10229),
.SN(net9550),
.CK(clk),
.Q(net10814),
.QN(net10813)
);

DFFS_X2 merge9913(
.D(net10703),
.SN(net1534),
.CK(clk),
.Q(net10816),
.QN(net10815)
);

CLKGATETST_X1 merge9914(
.E(net10011),
.SE(net10591),
.CK(clk),
.GCK(net10817)
);

AND2_X2 merge9915(
.A1(net6535),
.A2(net6435),
.ZN(net10818)
);

CLKGATETST_X2 merge9916(
.E(net8390),
.SE(net9230),
.CK(clk),
.GCK(net10819)
);

CLKGATETST_X4 merge9917(
.E(net6711),
.SE(net9360),
.CK(clk),
.GCK(net10820)
);

CLKGATETST_X8 merge9918(
.E(net10251),
.SE(net10520),
.CK(clk),
.GCK(net10821)
);

DFFR_X1 merge9919(
.D(net4734),
.RN(net4710),
.CK(clk),
.Q(net10823),
.QN(net10822)
);

DFFR_X2 merge9920(
.D(net9826),
.RN(net10339),
.CK(clk),
.Q(net10825),
.QN(net10824)
);

DFFS_X1 merge9921(
.D(net1463),
.SN(net10535),
.CK(clk),
.Q(net10827),
.QN(net10826)
);

DFFS_X2 merge9922(
.D(net8874),
.SN(net9015),
.CK(clk),
.Q(net10829),
.QN(net10828)
);

CLKGATETST_X1 merge9923(
.E(net10195),
.SE(net9879),
.CK(clk),
.GCK(net10830)
);

CLKGATETST_X2 merge9924(
.E(net6411),
.SE(net9779),
.CK(clk),
.GCK(net10831)
);

CLKGATETST_X4 merge9925(
.E(net8600),
.SE(net8538),
.CK(clk),
.GCK(net10832)
);

CLKGATETST_X8 merge9926(
.E(net9610),
.SE(net10110),
.CK(clk),
.GCK(net10833)
);

DFFR_X1 merge9927(
.D(net10274),
.RN(net2556),
.CK(clk),
.Q(net10835),
.QN(net10834)
);

DFFR_X2 merge9928(
.D(net6638),
.RN(net6630),
.CK(clk),
.Q(net10837),
.QN(net10836)
);

DFFS_X1 merge9929(
.D(net7428),
.SN(net7331),
.CK(clk),
.Q(net10839),
.QN(net10838)
);

DFFS_X2 merge9930(
.D(net10498),
.SN(net10207),
.CK(clk),
.Q(net10841),
.QN(net10840)
);

CLKGATETST_X1 merge9931(
.E(net9173),
.SE(net9139),
.CK(clk),
.GCK(net10842)
);

CLKGATETST_X2 merge9932(
.E(net8990),
.SE(net8802),
.CK(clk),
.GCK(net10843)
);

CLKGATETST_X4 merge9933(
.E(net6722),
.SE(net9534),
.CK(clk),
.GCK(net10844)
);

CLKGATETST_X8 merge9934(
.E(net10553),
.SE(net6104),
.CK(clk),
.GCK(net10845)
);

DFFR_X1 merge9935(
.D(net4943),
.RN(net3995),
.CK(clk),
.Q(net10847),
.QN(net10846)
);

DFFR_X2 merge9936(
.D(net8044),
.RN(net8046),
.CK(clk),
.Q(net10849),
.QN(net10848)
);

DFFS_X1 merge9937(
.D(net10061),
.SN(net10074),
.CK(clk),
.Q(net10851),
.QN(net10850)
);

XOR2_X1 merge9938(
.A(net7928),
.B(net8841),
.Z(net10852)
);

DFFS_X2 merge9939(
.D(net2280),
.SN(net10134),
.CK(clk),
.Q(net10854),
.QN(net10853)
);

CLKGATETST_X1 merge9940(
.E(net7647),
.SE(net8425),
.CK(clk),
.GCK(net10855)
);

CLKGATETST_X2 merge9941(
.E(net802),
.SE(net2762),
.CK(clk),
.GCK(net10856)
);

CLKGATETST_X4 merge9942(
.E(net1443),
.SE(net10034),
.CK(clk),
.GCK(net10857)
);

CLKGATETST_X8 merge9943(
.E(net3588),
.SE(net10455),
.CK(clk),
.GCK(net10858)
);

DFFR_X1 merge9944(
.D(net6620),
.RN(net1606),
.CK(clk),
.Q(net10860),
.QN(net10859)
);

DFFR_X2 merge9945(
.D(net9192),
.RN(net7631),
.CK(clk),
.Q(net10862),
.QN(net10861)
);

DFFS_X1 merge9946(
.D(net9053),
.SN(net8282),
.CK(clk),
.Q(net10864),
.QN(net10863)
);

DFFS_X2 merge9947(
.D(net9468),
.SN(net9262),
.CK(clk),
.Q(net10866),
.QN(net10865)
);

CLKGATETST_X1 merge9948(
.E(net9147),
.SE(net8953),
.CK(clk),
.GCK(net10867)
);

CLKGATETST_X2 merge9949(
.E(net10135),
.SE(net10504),
.CK(clk),
.GCK(net10868)
);

CLKGATETST_X4 merge9950(
.E(net10325),
.SE(net1221),
.CK(clk),
.GCK(net10869)
);

CLKGATETST_X8 merge9951(
.E(net9936),
.SE(net9595),
.CK(clk),
.GCK(net10870)
);

DFFR_X1 merge9952(
.D(net9458),
.RN(net9385),
.CK(clk),
.Q(net10872),
.QN(net10871)
);

DFFR_X2 merge9953(
.D(net6677),
.RN(net6708),
.CK(clk),
.Q(net10873),
.QN(out5)
);

DFFS_X1 merge9954(
.D(net10539),
.SN(net10580),
.CK(clk),
.Q(net10875),
.QN(net10874)
);

DFFS_X2 merge9955(
.D(net8584),
.SN(net9263),
.CK(clk),
.Q(net10877),
.QN(net10876)
);

CLKGATETST_X1 merge9956(
.E(net9453),
.SE(net9398),
.CK(clk),
.GCK(net10878)
);

CLKGATETST_X2 merge9957(
.E(net7606),
.SE(net7580),
.CK(clk),
.GCK(net10879)
);

NOR2_X1 merge9958(
.A1(net9302),
.A2(net9219),
.ZN(net10880)
);

CLKGATETST_X4 merge9959(
.E(net9187),
.SE(net8476),
.CK(clk),
.GCK(net10881)
);

CLKGATETST_X8 merge9960(
.E(net3605),
.SE(net2628),
.CK(clk),
.GCK(net10882)
);

DFFR_X1 merge9961(
.D(net9858),
.RN(net10306),
.CK(clk),
.Q(net10884),
.QN(net10883)
);

DFFR_X2 merge9962(
.D(net8460),
.RN(net9355),
.CK(clk),
.Q(net10886),
.QN(net10885)
);

DFFS_X1 merge9963(
.D(net8613),
.SN(net7671),
.CK(clk),
.Q(net10888),
.QN(net10887)
);

DFFS_X2 merge9964(
.D(net1260),
.SN(net9895),
.CK(clk),
.Q(net10890),
.QN(net10889)
);

OR2_X2 merge9965(
.A1(net9040),
.A2(net9073),
.ZN(net10891)
);

CLKGATETST_X1 merge9966(
.E(net8609),
.SE(net7661),
.CK(clk),
.GCK(net10892)
);

CLKGATETST_X2 merge9967(
.E(net9050),
.SE(net8873),
.CK(clk),
.GCK(net10893)
);

CLKGATETST_X4 merge9968(
.E(net7692),
.SE(net7629),
.CK(clk),
.GCK(net10894)
);

CLKGATETST_X8 merge9969(
.E(net7698),
.SE(net8261),
.CK(clk),
.GCK(net10895)
);

DFFR_X1 merge9970(
.D(net438),
.RN(net3246),
.CK(clk),
.Q(net10897),
.QN(net10896)
);

DFFR_X2 merge9971(
.D(net10661),
.RN(net10053),
.CK(clk),
.Q(net10899),
.QN(net10898)
);

DFFS_X1 merge9972(
.D(net8871),
.SN(net9038),
.CK(clk),
.Q(net10901),
.QN(net10900)
);

DFFS_X2 merge9973(
.D(net10189),
.SN(net3602),
.CK(clk),
.Q(net10903),
.QN(net10902)
);

CLKGATETST_X1 merge9974(
.E(net4056),
.SE(net10499),
.CK(clk),
.GCK(net10904)
);

CLKGATETST_X2 merge9975(
.E(net9671),
.SE(net659),
.CK(clk),
.GCK(net10905)
);

CLKGATETST_X4 merge9976(
.E(net8228),
.SE(net9333),
.CK(clk),
.GCK(net10906)
);

CLKGATETST_X8 merge9977(
.E(net4128),
.SE(net9820),
.CK(clk),
.GCK(net10907)
);

DFFR_X1 merge9978(
.D(net6102),
.RN(net10113),
.CK(clk),
.Q(net10909),
.QN(net10908)
);

DFFR_X2 merge9979(
.D(net8426),
.RN(net8455),
.CK(clk),
.Q(net10911),
.QN(net10910)
);

DFFS_X1 merge9980(
.D(net10632),
.SN(net10332),
.CK(clk),
.Q(net10913),
.QN(net10912)
);

DFFS_X2 merge9981(
.D(net10460),
.SN(net6101),
.CK(clk),
.Q(net10915),
.QN(net10914)
);

CLKGATETST_X1 merge9982(
.E(net10106),
.SE(net10228),
.CK(clk),
.GCK(net10916)
);

CLKGATETST_X2 merge9983(
.E(net9346),
.SE(net9170),
.CK(clk),
.GCK(net10917)
);

CLKGATETST_X4 merge9984(
.E(net9148),
.SE(net9129),
.CK(clk),
.GCK(net10918)
);

CLKGATETST_X8 merge9985(
.E(net7697),
.SE(net7660),
.CK(clk),
.GCK(net10919)
);

DFFR_X1 merge9986(
.D(net10666),
.RN(net3181),
.CK(clk),
.Q(net10921),
.QN(net10920)
);

DFFR_X2 merge9987(
.D(net9297),
.RN(net8471),
.CK(clk),
.Q(net10923),
.QN(net10922)
);

DFFS_X1 merge9988(
.D(net7538),
.SN(net7572),
.CK(clk),
.Q(net10925),
.QN(net10924)
);

DFFS_X2 merge9989(
.D(net9655),
.SN(net10156),
.CK(clk),
.Q(net10927),
.QN(net10926)
);

CLKGATETST_X1 merge9990(
.E(net9248),
.SE(net10459),
.CK(clk),
.GCK(net10928)
);

CLKGATETST_X2 merge9991(
.E(net8530),
.SE(net9443),
.CK(clk),
.GCK(net10929)
);

CLKGATETST_X4 merge9992(
.E(net10404),
.SE(net2643),
.CK(clk),
.GCK(net10930)
);

CLKGATETST_X8 merge9993(
.E(net9613),
.SE(net10062),
.CK(clk),
.GCK(net10931)
);

DFFR_X1 merge9994(
.D(net10471),
.RN(net10309),
.CK(clk),
.Q(net10933),
.QN(net10932)
);

DFFR_X2 merge9995(
.D(net9481),
.RN(net9446),
.CK(clk),
.Q(net10935),
.QN(net10934)
);

DFFS_X1 merge9996(
.D(net10177),
.SN(net4182),
.CK(clk),
.Q(net10937),
.QN(net10936)
);

DFFS_X2 merge9997(
.D(net9954),
.SN(net10071),
.CK(clk),
.Q(net10939),
.QN(net10938)
);

NOR2_X4 merge9998(
.A1(net9378),
.A2(net8416),
.ZN(net10940)
);

CLKGATETST_X1 merge9999(
.E(net7575),
.SE(net7669),
.CK(clk),
.GCK(net10941)
);

CLKGATETST_X2 merge10000(
.E(net9964),
.SE(net9777),
.CK(clk),
.GCK(net10942)
);

CLKGATETST_X4 merge10001(
.E(net7685),
.SE(net9440),
.CK(clk),
.GCK(net10943)
);

CLKGATETST_X8 merge10002(
.E(net4589),
.SE(net5556),
.CK(clk),
.GCK(net10944)
);

DFFR_X1 merge10003(
.D(net10379),
.RN(net10092),
.CK(clk),
.Q(net10946),
.QN(net10945)
);

DFFR_X2 merge10004(
.D(net8515),
.RN(net9452),
.CK(clk),
.Q(net10948),
.QN(net10947)
);

DFFS_X1 merge10005(
.D(net2122),
.SN(net231),
.CK(clk),
.Q(net10950),
.QN(net10949)
);

DFFS_X2 merge10006(
.D(net8401),
.SN(net10612),
.CK(clk),
.Q(net10952),
.QN(net10951)
);

CLKGATETST_X1 merge10007(
.E(net10431),
.SE(net7689),
.CK(clk),
.GCK(net10953)
);

CLKGATETST_X2 merge10008(
.E(net8832),
.SE(net7931),
.CK(clk),
.GCK(net10954)
);

CLKGATETST_X4 merge10009(
.E(net3282),
.SE(net1352),
.CK(clk),
.GCK(net10955)
);

CLKGATETST_X8 merge10010(
.E(net6924),
.SE(net7935),
.CK(clk),
.GCK(net10956)
);

DFFR_X1 merge10011(
.D(net9641),
.RN(net9603),
.CK(clk),
.Q(net10958),
.QN(net10957)
);

DFFR_X2 merge10012(
.D(net10292),
.RN(net10698),
.CK(clk),
.Q(net10960),
.QN(net10959)
);

DFFS_X1 merge10013(
.D(net9379),
.SN(net8465),
.CK(clk),
.Q(net10962),
.QN(net10961)
);

DFFS_X2 merge10014(
.D(net9652),
.SN(net10168),
.CK(clk),
.Q(net10964),
.QN(net10963)
);

CLKGATETST_X1 merge10015(
.E(net9317),
.SE(net9363),
.CK(clk),
.GCK(net10965)
);

CLKGATETST_X2 merge10016(
.E(net9456),
.SE(net8585),
.CK(clk),
.GCK(net10966)
);

CLKGATETST_X4 merge10017(
.E(net8148),
.SE(net10627),
.CK(clk),
.GCK(net10967)
);

CLKGATETST_X8 merge10018(
.E(net7679),
.SE(net9473),
.CK(clk),
.GCK(net10968)
);

DFFR_X1 merge10019(
.D(net8534),
.RN(net9747),
.CK(clk),
.Q(net10970),
.QN(net10969)
);

DFFR_X2 merge10020(
.D(net3635),
.RN(net10424),
.CK(clk),
.Q(net10972),
.QN(net10971)
);

DFFS_X1 merge10021(
.D(net10224),
.SN(net10508),
.CK(clk),
.Q(net10974),
.QN(net10973)
);

DFFS_X2 merge10022(
.D(net10220),
.SN(net2117),
.CK(clk),
.Q(net10976),
.QN(net10975)
);

CLKGATETST_X1 merge10023(
.E(net8598),
.SE(net8604),
.CK(clk),
.GCK(out23)
);

CLKGATETST_X2 merge10024(
.E(net1368),
.SE(net3315),
.CK(clk),
.GCK(net10977)
);

CLKGATETST_X4 merge10025(
.E(net9993),
.SE(net10093),
.CK(clk),
.GCK(net10978)
);

CLKGATETST_X8 merge10026(
.E(net10638),
.SE(net10669),
.CK(clk),
.GCK(net10979)
);

NOR2_X2 merge10027(
.A1(net9406),
.A2(net9431),
.ZN(net10980)
);

DFFR_X1 merge10028(
.D(net8632),
.RN(net8606),
.CK(clk),
.Q(net10982),
.QN(net10981)
);

DFFR_X2 merge10029(
.D(net10094),
.RN(net6112),
.CK(clk),
.Q(net10984),
.QN(net10983)
);

DFFS_X1 merge10030(
.D(net9887),
.SN(net10351),
.CK(clk),
.Q(net10986),
.QN(net10985)
);

DFFS_X2 merge10031(
.D(net7683),
.SN(net7686),
.CK(clk),
.Q(net10988),
.QN(net10987)
);

CLKGATETST_X1 merge10032(
.E(net10393),
.SE(net10377),
.CK(clk),
.GCK(net10989)
);

CLKGATETST_X2 merge10033(
.E(net9503),
.SE(net9430),
.CK(clk),
.GCK(net10990)
);

CLKGATETST_X4 merge10034(
.E(net8636),
.SE(net8610),
.CK(clk),
.GCK(net10991)
);

CLKGATETST_X8 merge10035(
.E(net10007),
.SE(net10560),
.CK(clk),
.GCK(net10992)
);

XOR2_X2 merge10036(
.A(net9495),
.B(net8617),
.Z(net10993)
);

DFFR_X1 merge10037(
.D(net10391),
.RN(net10070),
.CK(clk),
.Q(net10995),
.QN(net10994)
);

DFFR_X2 merge10038(
.D(net10239),
.RN(net9883),
.CK(clk),
.Q(net10997),
.QN(net10996)
);

DFFS_X1 merge10039(
.D(net10495),
.SN(net10163),
.CK(clk),
.Q(net10999),
.QN(net10998)
);

DFFS_X2 merge10040(
.D(net8605),
.Q(net11000),
.CK(clk),
.QN(out2)
);

CLKGATETST_X1 merge10041(
.E(net10741),
.SE(net7162),
.CK(clk),
.GCK(net11001)
);

CLKGATETST_X2 merge10042(
.E(net1518),
.SE(net10650),
.CK(clk),
.GCK(net11002)
);

CLKGATETST_X4 merge10043(
.E(net10710),
.SE(net9587),
.CK(clk),
.GCK(net11003)
);

CLKGATETST_X8 merge10044(
.E(net10511),
.SE(net4313),
.CK(clk),
.GCK(net11004)
);

DFFR_X1 merge10045(
.D(net10208),
.RN(net10697),
.CK(clk),
.Q(net11006),
.QN(net11005)
);

DFFR_X2 merge10046(
.D(net9496),
.RN(net9513),
.CK(clk),
.Q(net11008),
.QN(net11007)
);

DFFS_X1 merge10047(
.D(net10014),
.SN(net10350),
.CK(clk),
.Q(net11010),
.QN(net11009)
);

DFFS_X2 merge10048(
.D(net8615),
.SN(net8616),
.CK(clk),
.Q(out10),
.QN(net11011)
);

CLKGATETST_X1 merge10049(
.E(net2189),
.SE(net10326),
.CK(clk),
.GCK(net11012)
);

CLKGATETST_X2 merge10050(
.E(net4232),
.SE(net10592),
.CK(clk),
.GCK(net11013)
);

CLKGATETST_X4 merge10051(
.E(net9528),
.SE(net9529),
.CK(clk),
.GCK(net11014)
);

CLKGATETST_X8 merge10052(
.E(net10095),
.SE(net5091),
.CK(clk),
.GCK(net11015)
);

DFFR_X1 merge10053(
.D(net9535),
.RN(net8618),
.CK(clk),
.Q(net11016),
.QN(out7)
);

DFFR_X2 merge10054(
.D(net10891),
.RN(net9598),
.CK(clk),
.Q(net11018),
.QN(net11017)
);

DFFS_X1 merge10055(
.D(net9907),
.SN(net9768),
.CK(clk),
.Q(net11020),
.QN(net11019)
);

DFFS_X2 merge10056(
.D(net9949),
.SN(net10037),
.CK(clk),
.Q(net11022),
.QN(net11021)
);

CLKGATETST_X1 merge10057(
.E(net9708),
.SE(net10557),
.CK(clk),
.GCK(net11023)
);

CLKGATETST_X2 merge10058(
.E(net10109),
.SE(net2115),
.CK(clk),
.GCK(net11024)
);

CLKGATETST_X4 merge10059(
.E(net9869),
.SE(net3724),
.CK(clk),
.GCK(net11025)
);

CLKGATETST_X8 merge10060(
.E(net10940),
.SE(net6602),
.CK(clk),
.GCK(net11026)
);

DFFR_X1 merge10061(
.D(net10537),
.RN(net10620),
.CK(clk),
.Q(net11028),
.QN(net11027)
);

DFFR_X2 merge10062(
.D(net10127),
.RN(net10630),
.CK(clk),
.Q(net11030),
.QN(net11029)
);

DFFS_X1 merge10063(
.D(net10652),
.SN(net1456),
.CK(clk),
.Q(net11032),
.QN(net11031)
);

DFFS_X2 merge10064(
.D(net9952),
.SN(net2709),
.CK(clk),
.Q(net11034),
.QN(net11033)
);

CLKGATETST_X1 merge10065(
.E(net10715),
.SE(net9985),
.CK(clk),
.GCK(net11035)
);

CLKGATETST_X2 merge10066(
.E(net10365),
.SE(net6408),
.CK(clk),
.GCK(net11036)
);

CLKGATETST_X4 merge10067(
.E(net10534),
.SE(net10469),
.CK(clk),
.GCK(net11037)
);

CLKGATETST_X8 merge10068(
.E(net9596),
.SE(net2321),
.CK(clk),
.GCK(net11038)
);

DFFR_X1 merge10069(
.D(net9920),
.RN(net10597),
.CK(clk),
.Q(net11040),
.QN(net11039)
);

DFFR_X2 merge10070(
.D(net297),
.RN(net10596),
.CK(clk),
.Q(net11042),
.QN(net11041)
);

DFFS_X1 merge10071(
.D(net9769),
.SN(net9634),
.CK(clk),
.Q(net11044),
.QN(net11043)
);

DFFS_X2 merge10072(
.D(net7210),
.SN(net10331),
.CK(clk),
.Q(net11046),
.QN(net11045)
);

CLKGATETST_X1 merge10073(
.E(net467),
.SE(net10042),
.CK(clk),
.GCK(net11047)
);

CLKGATETST_X2 merge10074(
.E(net10440),
.SE(net9923),
.CK(clk),
.GCK(net11048)
);

CLKGATETST_X4 merge10075(
.E(net4269),
.SE(net2130),
.CK(clk),
.GCK(net11049)
);

CLKGATETST_X8 merge10076(
.E(net9705),
.SE(net10604),
.CK(clk),
.GCK(net11050)
);

DFFR_X1 merge10077(
.D(net10713),
.RN(net9906),
.CK(clk),
.Q(net11052),
.QN(net11051)
);

DFFR_X2 merge10078(
.D(net9742),
.RN(net10686),
.CK(clk),
.Q(net11054),
.QN(net11053)
);

DFFS_X1 merge10079(
.D(net10314),
.SN(net10357),
.CK(clk),
.Q(net11056),
.QN(net11055)
);

DFFS_X2 merge10080(
.D(net9831),
.SN(net9859),
.CK(clk),
.Q(net11058),
.QN(net11057)
);

CLKGATETST_X1 merge10081(
.E(net9953),
.SE(net9860),
.CK(clk),
.GCK(net11059)
);

CLKGATETST_X2 merge10082(
.E(net5215),
.SE(net10077),
.CK(clk),
.GCK(net11060)
);

CLKGATETST_X4 merge10083(
.E(net10082),
.SE(net10993),
.CK(clk),
.GCK(net11061)
);

CLKGATETST_X8 merge10084(
.E(net9937),
.SE(net7486),
.CK(clk),
.GCK(net11062)
);

DFFR_X1 merge10085(
.D(net10167),
.RN(net10687),
.CK(clk),
.Q(net11064),
.QN(net11063)
);

DFFR_X2 merge10086(
.D(net10779),
.RN(net10091),
.CK(clk),
.Q(net11066),
.QN(net11065)
);

DFFS_X1 merge10087(
.D(net10796),
.SN(net9329),
.CK(clk),
.Q(net11068),
.QN(net11067)
);

DFFS_X2 merge10088(
.D(net10575),
.SN(net10456),
.CK(clk),
.Q(net11070),
.QN(net11069)
);

CLKGATETST_X1 merge10089(
.E(net6448),
.SE(net6181),
.CK(clk),
.GCK(net11071)
);

CLKGATETST_X2 merge10090(
.E(net10164),
.SE(net9935),
.CK(clk),
.GCK(net11072)
);

CLKGATETST_X4 merge10091(
.E(net9867),
.SE(net9563),
.CK(clk),
.GCK(net11073)
);

CLKGATETST_X8 merge10092(
.E(net9636),
.SE(net4259),
.CK(clk),
.GCK(net11074)
);

DFFR_X1 merge10093(
.D(net9809),
.RN(net1481),
.CK(clk),
.Q(net11076),
.QN(net11075)
);

DFFR_X2 merge10094(
.D(net10214),
.RN(net10792),
.CK(clk),
.Q(net11078),
.QN(net11077)
);

DFFS_X1 merge10095(
.D(net10467),
.SN(net9872),
.CK(clk),
.Q(net11080),
.QN(net11079)
);

DFFS_X2 merge10096(
.D(net10556),
.SN(net10468),
.CK(clk),
.Q(net11082),
.QN(net11081)
);

CLKGATETST_X1 merge10097(
.E(net10285),
.SE(net7340),
.CK(clk),
.GCK(net11083)
);

CLKGATETST_X2 merge10098(
.E(net9973),
.SE(net10090),
.CK(clk),
.GCK(net11084)
);

CLKGATETST_X4 merge10099(
.E(net10140),
.SE(net10145),
.CK(clk),
.GCK(net11085)
);

CLKGATETST_X8 merge10100(
.E(net4065),
.SE(net10696),
.CK(clk),
.GCK(net11086)
);

DFFR_X1 merge10101(
.D(net10083),
.RN(net10599),
.CK(clk),
.Q(net11088),
.QN(net11087)
);

DFFR_X2 merge10102(
.D(net10880),
.RN(net9373),
.CK(clk),
.Q(net11090),
.QN(net11089)
);

DFFS_X1 merge10103(
.D(net9559),
.SN(net10704),
.CK(clk),
.Q(net11092),
.QN(net11091)
);

DFFS_X2 merge10104(
.D(net9944),
.SN(net10490),
.CK(clk),
.Q(net11094),
.QN(net11093)
);

CLKGATETST_X1 merge10105(
.E(net10394),
.SE(net8259),
.CK(clk),
.GCK(net11095)
);

CLKGATETST_X2 merge10106(
.E(net8220),
.SE(net10645),
.CK(clk),
.GCK(net11096)
);

CLKGATETST_X4 merge10107(
.E(net6105),
.SE(net10435),
.CK(clk),
.GCK(net11097)
);

CLKGATETST_X8 merge10108(
.E(net10649),
.SE(net10664),
.CK(clk),
.GCK(net11098)
);

DFFR_X1 merge10109(
.D(net10705),
.RN(net10611),
.CK(clk),
.Q(net11100),
.QN(net11099)
);

DFFR_X2 merge10110(
.D(net10236),
.RN(net10023),
.CK(clk),
.Q(net11102),
.QN(net11101)
);

DFFS_X1 merge10111(
.D(net10487),
.SN(net10407),
.CK(clk),
.Q(net11104),
.QN(net11103)
);

DFFS_X2 merge10112(
.D(net9590),
.SN(net9623),
.CK(clk),
.Q(net11106),
.QN(net11105)
);

CLKGATETST_X1 merge10113(
.E(net10719),
.SE(net10598),
.CK(clk),
.GCK(net11107)
);

CLKGATETST_X2 merge10114(
.E(net10425),
.SE(net9787),
.CK(clk),
.GCK(net11108)
);

CLKGATETST_X4 merge10115(
.E(net10613),
.SE(net10818),
.CK(clk),
.GCK(net11109)
);

CLKGATETST_X8 merge10116(
.E(net8226),
.SE(net9662),
.CK(clk),
.GCK(net11110)
);

DFFR_X1 merge10117(
.D(net9617),
.RN(net9694),
.CK(clk),
.Q(net11112),
.QN(net11111)
);

DFFR_X2 merge10118(
.D(net9943),
.RN(net10420),
.CK(clk),
.Q(net11114),
.QN(net11113)
);

DFFS_X1 merge10119(
.D(net10297),
.SN(net10215),
.CK(clk),
.Q(net11116),
.QN(net11115)
);

DFFS_X2 merge10120(
.D(net9669),
.SN(net7060),
.CK(clk),
.Q(net11118),
.QN(net11117)
);

CLKGATETST_X1 merge10121(
.E(net9875),
.SE(net10980),
.CK(clk),
.GCK(net11119)
);

CLKGATETST_X2 merge10122(
.E(net3702),
.SE(net10069),
.CK(clk),
.GCK(net11120)
);

CLKGATETST_X4 merge10123(
.E(net2232),
.SE(net10718),
.CK(clk),
.GCK(net11121)
);

CLKGATETST_X8 merge10124(
.E(net10767),
.SE(net10225),
.CK(clk),
.GCK(out0)
);

DFFR_X1 merge10125(
.D(net9868),
.RN(net2672),
.CK(clk),
.Q(net11123),
.QN(net11122)
);

DFFR_X2 merge10126(
.D(net10354),
.RN(net10103),
.CK(clk),
.Q(net11125),
.QN(net11124)
);

DFFS_X1 merge10127(
.D(net9672),
.SN(net10486),
.CK(clk),
.Q(net11127),
.QN(net11126)
);

DFFS_X2 merge10128(
.D(net10275),
.SN(net10522),
.CK(clk),
.Q(net11129),
.QN(net11128)
);

CLKGATETST_X1 merge10129(
.E(net9942),
.SE(net10646),
.CK(clk),
.GCK(net11130)
);

CLKGATETST_X2 merge10130(
.E(net10574),
.SE(net7327),
.CK(clk),
.GCK(net11131)
);

CLKGATETST_X4 merge10131(
.E(net5212),
.SE(net10010),
.CK(clk),
.GCK(net11132)
);

CLKGATETST_X8 merge10132(
.E(net4599),
.SE(net10054),
.CK(clk),
.GCK(net11133)
);

DFFR_X1 merge10133(
.D(net9579),
.RN(net9957),
.CK(clk),
.Q(net11135),
.QN(net11134)
);

DFFR_X2 merge10134(
.D(net10681),
.RN(net10852),
.CK(clk),
.Q(net11137),
.QN(net11136)
);

DFFS_X1 merge10135(
.D(net6537),
.SN(net10223),
.CK(clk),
.Q(net11139),
.QN(net11138)
);

DFF_X1 s10136(
.D(net221),
.CK(clk),
.Q(net11141),
.QN(net11140)
);

DFF_X2 s10137(
.D(net561),
.CK(clk),
.Q(net11143),
.QN(net11142)
);

DFF_X1 s10138(
.D(net582),
.CK(clk),
.Q(net11145),
.QN(net11144)
);

DFF_X2 s10139(
.D(net583),
.CK(clk),
.Q(net11147),
.QN(net11146)
);

DFF_X1 s10140(
.D(net1039),
.CK(clk),
.Q(net11149),
.QN(net11148)
);

DFF_X2 s10141(
.D(net1100),
.CK(clk),
.Q(net11151),
.QN(net11150)
);

DFF_X1 s10142(
.D(net1191),
.CK(clk),
.Q(net11153),
.QN(net11152)
);

DFF_X2 s10143(
.D(net1511),
.CK(clk),
.Q(net11155),
.QN(net11154)
);

DFF_X1 s10144(
.D(net1858),
.CK(clk),
.Q(net11157),
.QN(net11156)
);

DFF_X2 s10145(
.D(net1980),
.CK(clk),
.Q(net11159),
.QN(net11158)
);

DFF_X1 s10146(
.D(net2296),
.CK(clk),
.Q(net11161),
.QN(net11160)
);

DFF_X2 s10147(
.D(net2408),
.CK(clk),
.Q(net11163),
.QN(net11162)
);

DFF_X1 s10148(
.D(net2413),
.CK(clk),
.Q(net11165),
.QN(net11164)
);

DFF_X2 s10149(
.D(net2418),
.CK(clk),
.Q(net11167),
.QN(net11166)
);

DFF_X1 s10150(
.D(net2858),
.CK(clk),
.Q(net11169),
.QN(net11168)
);

DFF_X2 s10151(
.D(net3461),
.CK(clk),
.Q(net11171),
.QN(net11170)
);

DFF_X1 s10152(
.D(net3622),
.CK(clk),
.Q(net11173),
.QN(net11172)
);

DFF_X2 s10153(
.D(net3890),
.CK(clk),
.Q(net11175),
.QN(net11174)
);

DFF_X1 s10154(
.D(net4074),
.CK(clk),
.Q(net11177),
.QN(net11176)
);

DFF_X2 s10155(
.D(net4110),
.CK(clk),
.Q(net11179),
.QN(net11178)
);

DFF_X1 s10156(
.D(net4262),
.CK(clk),
.Q(net11181),
.QN(net11180)
);

DFF_X2 s10157(
.D(net4752),
.CK(clk),
.Q(net11183),
.QN(net11182)
);

DFF_X1 s10158(
.D(net4765),
.CK(clk),
.Q(net11185),
.QN(net11184)
);

DFF_X2 s10159(
.D(net4874),
.CK(clk),
.Q(net11187),
.QN(net11186)
);

DFF_X1 s10160(
.D(net4968),
.CK(clk),
.Q(net11189),
.QN(net11188)
);

DFF_X2 s10161(
.D(net5202),
.CK(clk),
.Q(net11191),
.QN(net11190)
);

DFF_X1 s10162(
.D(net5675),
.CK(clk),
.Q(net11193),
.QN(net11192)
);

DFF_X2 s10163(
.D(net5759),
.CK(clk),
.Q(net11195),
.QN(net11194)
);

DFF_X1 s10164(
.D(net5844),
.CK(clk),
.Q(net11197),
.QN(net11196)
);

DFF_X2 s10165(
.D(net5942),
.CK(clk),
.Q(net11199),
.QN(net11198)
);

DFF_X1 s10166(
.D(net6541),
.CK(clk),
.Q(net11201),
.QN(net11200)
);

DFF_X2 s10167(
.D(net6805),
.CK(clk),
.Q(net11203),
.QN(net11202)
);

DFF_X1 s10168(
.D(net6811),
.CK(clk),
.Q(net11205),
.QN(net11204)
);

DFF_X2 s10169(
.D(net7157),
.CK(clk),
.Q(net11207),
.QN(net11206)
);

DFF_X1 s10170(
.D(net7336),
.CK(clk),
.Q(net11209),
.QN(net11208)
);

DFF_X2 s10171(
.D(net7517),
.CK(clk),
.Q(net11211),
.QN(net11210)
);

DFF_X1 s10172(
.D(net7766),
.CK(clk),
.Q(net11213),
.QN(net11212)
);

DFF_X2 s10173(
.D(net7786),
.CK(clk),
.Q(net11215),
.QN(net11214)
);

DFF_X1 s10174(
.D(net8051),
.CK(clk),
.Q(net11217),
.QN(net11216)
);

DFF_X2 s10175(
.D(net8131),
.CK(clk),
.Q(net11219),
.QN(net11218)
);

DFF_X1 s10176(
.D(net8277),
.CK(clk),
.Q(net11221),
.QN(net11220)
);

DFF_X2 s10177(
.D(net8288),
.CK(clk),
.Q(net11223),
.QN(net11222)
);

DFF_X1 s10178(
.D(net8397),
.CK(clk),
.Q(net11225),
.QN(net11224)
);

DFF_X2 s10179(
.D(net8729),
.CK(clk),
.Q(net11227),
.QN(net11226)
);

DFF_X1 s10180(
.D(net9077),
.CK(clk),
.Q(net11229),
.QN(net11228)
);

DFF_X2 s10181(
.D(net9211),
.CK(clk),
.Q(net11231),
.QN(net11230)
);

DFF_X1 s10182(
.D(net9368),
.CK(clk),
.Q(net11233),
.QN(net11232)
);

DFF_X2 s10183(
.D(net9451),
.CK(clk),
.Q(net11235),
.QN(net11234)
);

DFF_X1 s10184(
.D(net9614),
.CK(clk),
.Q(net11237),
.QN(net11236)
);


endmodule
