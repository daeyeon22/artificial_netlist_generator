module test_circuit (
	input in0,
	input in1,
	input in2,
	input in3,
	input in4,
	input in5,
	input in6,
	input in7,
	input in8,
	input in9,
	input in10,
	input in11,
	input in12,
	input in13,
	input in14,
	input in15,
	input in16,
	input in17,
	input in18,
	input in19,
	input in20,
	input in21,
	input in22,
	input in23,
	input in24,
	input in25,
	input clk,
	input rst,
	output out0,
	output out1,
	output out2,
	output out3,
	output out4,
	output out5,
	output out6,
	output out7,
	output out8,
	output out9,
	output out10,
	output out11,
	output out12,
	output out13,
	output out14,
	output out15,
	output out16,
	output out17,
	output out18,
	output out19,
	output out20,
	output out21,
	output out22,
	output out23,
	output out24,
	output out25
);


wire net10576;
wire net10575;
wire net10574;
wire net10572;
wire net10571;
wire net10567;
wire net10565;
wire net10564;
wire net10563;
wire net10561;
wire net10559;
wire net10558;
wire net10553;
wire net10552;
wire net10551;
wire net10549;
wire net10548;
wire net10546;
wire net10545;
wire net10544;
wire net10538;
wire net10535;
wire net10533;
wire net10532;
wire net10526;
wire net10524;
wire net10523;
wire net10522;
wire net10520;
wire net10519;
wire net10518;
wire net10517;
wire net10515;
wire net10511;
wire net10510;
wire net10509;
wire net10503;
wire net10498;
wire net10497;
wire net10494;
wire net10493;
wire net10492;
wire net10490;
wire net10487;
wire net10485;
wire net10482;
wire net10479;
wire net10475;
wire net10474;
wire net10473;
wire net10472;
wire net10505;
wire net10469;
wire net10468;
wire net10461;
wire net10456;
wire net10455;
wire net10453;
wire net10451;
wire net10448;
wire net10446;
wire net10445;
wire net10440;
wire net10439;
wire net10438;
wire net10436;
wire net10435;
wire net10433;
wire net10431;
wire net10430;
wire net10428;
wire net10425;
wire net10424;
wire net10423;
wire net10422;
wire net10419;
wire net10416;
wire net10414;
wire net10413;
wire net10412;
wire net10411;
wire net10409;
wire net10408;
wire net10404;
wire net10403;
wire net10401;
wire net10400;
wire net10398;
wire net10395;
wire net10394;
wire net10385;
wire net10384;
wire net10382;
wire net10381;
wire net10379;
wire net10378;
wire net10377;
wire net10376;
wire net10375;
wire net10368;
wire net10367;
wire net10364;
wire net10363;
wire net10358;
wire net10353;
wire net10348;
wire net10343;
wire net10341;
wire net10340;
wire net10339;
wire net10335;
wire net10334;
wire net10333;
wire net10332;
wire net10330;
wire net10329;
wire net10328;
wire net10326;
wire net10323;
wire net10322;
wire net10321;
wire net10320;
wire net10318;
wire net10317;
wire net10311;
wire net10310;
wire net10307;
wire net10306;
wire net10305;
wire net10303;
wire net10301;
wire net10300;
wire net10299;
wire net10297;
wire net10295;
wire net10293;
wire net10292;
wire net10291;
wire net10290;
wire net10288;
wire net10286;
wire net10285;
wire net10283;
wire net10280;
wire net10277;
wire net10276;
wire net10275;
wire net10274;
wire net10272;
wire net10271;
wire net10269;
wire net10268;
wire net10267;
wire net10266;
wire net10265;
wire net10260;
wire net10259;
wire net10257;
wire net10256;
wire net10255;
wire net10253;
wire net10252;
wire net10249;
wire net10248;
wire net10244;
wire net10242;
wire net10240;
wire net10239;
wire net10287;
wire net10238;
wire net10236;
wire net10235;
wire net10234;
wire net10232;
wire net10231;
wire net10229;
wire net10226;
wire net10225;
wire net10224;
wire net10222;
wire net10221;
wire net10219;
wire net10218;
wire net10216;
wire net10215;
wire net10214;
wire net10211;
wire net10210;
wire net10209;
wire net10204;
wire net10202;
wire net10201;
wire net10193;
wire net10190;
wire net10186;
wire net10185;
wire net10184;
wire net10183;
wire net10182;
wire net10181;
wire net10180;
wire net10179;
wire net10175;
wire net10174;
wire net10173;
wire net10169;
wire net10168;
wire net10167;
wire net10164;
wire out0;
wire net10160;
wire net10155;
wire net10154;
wire net10152;
wire net10151;
wire net10149;
wire net10146;
wire net10145;
wire net10228;
wire net10144;
wire net10141;
wire net10138;
wire net10136;
wire net10135;
wire net10132;
wire net10131;
wire net10129;
wire net10127;
wire net10126;
wire net10125;
wire net10124;
wire net10118;
wire net10117;
wire net10116;
wire net10114;
wire net10109;
wire net10108;
wire net10107;
wire net10105;
wire net10104;
wire net10102;
wire net10099;
wire net10098;
wire net10096;
wire net10095;
wire net10092;
wire out7;
wire net10091;
wire net10089;
wire net10088;
wire out10;
wire net10087;
wire net10086;
wire net10085;
wire net10082;
wire out2;
wire net10080;
wire net10075;
wire net10073;
wire net10324;
wire net10072;
wire net10071;
wire net10070;
wire net10067;
wire net10066;
wire net10064;
wire net10061;
wire net10053;
wire net10051;
wire net10048;
wire net10047;
wire net10046;
wire net10044;
wire net10043;
wire net10042;
wire net10041;
wire net10039;
wire net10033;
wire net10031;
wire net10030;
wire net10028;
wire net10027;
wire net10024;
wire net10022;
wire net10020;
wire net10017;
wire net10016;
wire net10015;
wire net10011;
wire net10009;
wire net10153;
wire net10008;
wire net10005;
wire net10001;
wire net10000;
wire net9997;
wire out5;
wire net9992;
wire net9991;
wire net9988;
wire net9987;
wire net9985;
wire net9983;
wire net9982;
wire net9980;
wire net9979;
wire net9978;
wire net9976;
wire net9975;
wire net9974;
wire net9973;
wire net9970;
wire net9968;
wire net10465;
wire net9966;
wire net9961;
wire net9960;
wire net9959;
wire net9958;
wire net9957;
wire net9953;
wire net10566;
wire net9951;
wire net9948;
wire net9947;
wire net9938;
wire net9937;
wire net9935;
wire net9934;
wire net9931;
wire net9927;
wire net9925;
wire net9924;
wire net9923;
wire net9922;
wire net9918;
wire net9917;
wire net9916;
wire net9912;
wire net9911;
wire net9995;
wire net9909;
wire net9908;
wire net10270;
wire net9907;
wire net9906;
wire net9905;
wire net9901;
wire net9900;
wire net9899;
wire net9898;
wire net9896;
wire net10464;
wire net9894;
wire net9893;
wire net9891;
wire net9887;
wire net9884;
wire net9883;
wire net9881;
wire net9879;
wire net9878;
wire net9877;
wire net9876;
wire net9871;
wire net9870;
wire net10337;
wire net9869;
wire net9868;
wire net9865;
wire net9863;
wire net9862;
wire net10060;
wire net9861;
wire net9860;
wire net9859;
wire net9858;
wire net9857;
wire net10246;
wire net9856;
wire net9855;
wire net9852;
wire net9850;
wire net9847;
wire net9845;
wire net9843;
wire net10189;
wire net9932;
wire net9841;
wire net9839;
wire net9836;
wire net9833;
wire net9831;
wire net10489;
wire net9830;
wire net9826;
wire net9825;
wire net9823;
wire net9822;
wire net9821;
wire net9820;
wire net9816;
wire net9812;
wire net9809;
wire net9807;
wire net9805;
wire net10313;
wire net9803;
wire net9802;
wire net9801;
wire net9798;
wire net9797;
wire net9796;
wire net9795;
wire net9791;
wire net9790;
wire net9789;
wire net10296;
wire net9788;
wire net9786;
wire net9785;
wire net9783;
wire net9781;
wire net9780;
wire net9778;
wire net9774;
wire net9773;
wire net9772;
wire net9769;
wire net9768;
wire net9766;
wire net9765;
wire net9764;
wire net9761;
wire net9760;
wire net9759;
wire net9758;
wire net9757;
wire net9756;
wire net9755;
wire net9751;
wire net9750;
wire net9749;
wire net9748;
wire net9747;
wire net9746;
wire net9743;
wire net9742;
wire net9741;
wire net9739;
wire net9738;
wire net9737;
wire net9735;
wire net9777;
wire net9734;
wire net9732;
wire net9731;
wire net9729;
wire net9727;
wire net9726;
wire net9724;
wire net9723;
wire net9721;
wire net9720;
wire net9715;
wire net9711;
wire net9709;
wire net9708;
wire net9704;
wire net9703;
wire net9700;
wire net9699;
wire net9696;
wire net9695;
wire net9694;
wire net9693;
wire net9692;
wire net9691;
wire net9690;
wire net9689;
wire net9688;
wire net9685;
wire net9683;
wire net9682;
wire net9680;
wire net9678;
wire net9677;
wire net9675;
wire net9673;
wire net9672;
wire net9671;
wire net10369;
wire net9668;
wire net9667;
wire net9665;
wire net10187;
wire net9663;
wire net9661;
wire net9660;
wire net9659;
wire net9657;
wire net9653;
wire net9651;
wire net9679;
wire net9650;
wire net9649;
wire net9648;
wire net9647;
wire net9645;
wire net9641;
wire net9640;
wire net9638;
wire net10282;
wire net9634;
wire net9631;
wire net9629;
wire net9628;
wire net9625;
wire net9623;
wire net9622;
wire net9621;
wire net9753;
wire net9618;
wire net10018;
wire net9617;
wire net9616;
wire net9613;
wire net9612;
wire net9610;
wire net9607;
wire net9606;
wire net9604;
wire net10162;
wire net9603;
wire net9602;
wire net9601;
wire net9600;
wire net9598;
wire net9597;
wire net9596;
wire net9594;
wire net9592;
wire net9591;
wire net9589;
wire net9588;
wire net9587;
wire net9585;
wire net9583;
wire net9581;
wire net10279;
wire net9580;
wire net9579;
wire net9578;
wire net9576;
wire net9575;
wire net9574;
wire net10142;
wire net9573;
wire net9571;
wire net9570;
wire net9568;
wire net9565;
wire net9561;
wire net9555;
wire net9548;
wire net9547;
wire net9545;
wire net9544;
wire net9538;
wire net9537;
wire net9535;
wire net9534;
wire net9533;
wire net9529;
wire net9528;
wire net9525;
wire net9524;
wire net9519;
wire net9518;
wire net9516;
wire net9515;
wire net9514;
wire net9513;
wire net9512;
wire net9511;
wire net9508;
wire net9507;
wire net9506;
wire net9505;
wire net9504;
wire net9503;
wire net9502;
wire net9500;
wire net9499;
wire net9496;
wire net9492;
wire net9484;
wire net10365;
wire net9483;
wire net9479;
wire net9474;
wire net9473;
wire net9470;
wire net9469;
wire net9467;
wire net9464;
wire net9462;
wire net10254;
wire net9459;
wire net9457;
wire net9455;
wire net9454;
wire net9452;
wire net9449;
wire net9448;
wire net9444;
wire net9443;
wire net9439;
wire net9438;
wire net9437;
wire net9436;
wire net9434;
wire net9432;
wire net9431;
wire net9430;
wire net9429;
wire net9427;
wire net9424;
wire net9423;
wire net9422;
wire net9421;
wire net9419;
wire net9418;
wire net9416;
wire net9415;
wire net9412;
wire net9411;
wire net9632;
wire net9407;
wire net9406;
wire net9405;
wire net9404;
wire net9399;
wire net9398;
wire net9394;
wire net9393;
wire net9392;
wire net9390;
wire net9389;
wire net9387;
wire net9386;
wire net9385;
wire net9384;
wire net9383;
wire net9381;
wire net9378;
wire net9377;
wire net9376;
wire net9375;
wire net9373;
wire net9369;
wire net9364;
wire net9363;
wire net9362;
wire net9361;
wire net9360;
wire net9358;
wire net9357;
wire net9356;
wire net9352;
wire net9351;
wire net9350;
wire net10396;
wire net9349;
wire net9347;
wire net9346;
wire net9344;
wire net9343;
wire net9342;
wire net9341;
wire net9338;
wire net9337;
wire net9336;
wire net9333;
wire net9332;
wire net9331;
wire net9330;
wire net9326;
wire net9325;
wire net9324;
wire net9323;
wire net9320;
wire net9316;
wire net10161;
wire net9315;
wire net9314;
wire net9313;
wire net9311;
wire net9310;
wire net9309;
wire net9306;
wire net9305;
wire net9304;
wire net10525;
wire net9303;
wire net10094;
wire net9300;
wire net9299;
wire net9298;
wire net9294;
wire net9293;
wire net9291;
wire net9290;
wire net9295;
wire net9289;
wire net9288;
wire net9283;
wire net9282;
wire net9281;
wire net9280;
wire net9278;
wire net9276;
wire net9275;
wire net9269;
wire net9268;
wire net9266;
wire net9265;
wire net9263;
wire net9261;
wire net9256;
wire net9253;
wire net9252;
wire net9251;
wire net9250;
wire net9248;
wire net9244;
wire net9240;
wire net9239;
wire net9237;
wire net9236;
wire net9234;
wire net9231;
wire net9228;
wire net9227;
wire net9226;
wire net9339;
wire net9224;
wire net9222;
wire net9221;
wire net9220;
wire net9215;
wire net9213;
wire net9212;
wire net9211;
wire net9210;
wire net9209;
wire net9208;
wire net9207;
wire net9205;
wire net10176;
wire net9204;
wire net9200;
wire net9199;
wire net9197;
wire net9195;
wire net9194;
wire net9193;
wire net9190;
wire net9188;
wire net9185;
wire net9183;
wire net10506;
wire net9182;
wire net9536;
wire net9181;
wire net9180;
wire net9178;
wire net9176;
wire net9175;
wire net9171;
wire net9167;
wire net9166;
wire net9165;
wire net9164;
wire net9161;
wire net9160;
wire net9159;
wire net9158;
wire net9258;
wire net9157;
wire net9156;
wire net9154;
wire net9153;
wire net9152;
wire net9151;
wire net9147;
wire net9146;
wire net9145;
wire net9144;
wire net10447;
wire net9142;
wire net9141;
wire net9139;
wire net9136;
wire net9133;
wire net9132;
wire net9131;
wire net9130;
wire net9967;
wire net9126;
wire net9116;
wire net9174;
wire net9114;
wire net9112;
wire net9108;
wire net9107;
wire net9106;
wire net9105;
wire net9103;
wire net9100;
wire net9099;
wire net9095;
wire net9091;
wire net9090;
wire net9089;
wire net9088;
wire net9087;
wire net9674;
wire net9086;
wire net9084;
wire net9083;
wire net9081;
wire net9080;
wire net9076;
wire net9075;
wire net9488;
wire net9074;
wire net9073;
wire net9071;
wire net9069;
wire net9068;
wire net9063;
wire net9061;
wire net9059;
wire net9058;
wire net9057;
wire net9056;
wire net9710;
wire net9054;
wire net9053;
wire net9052;
wire net9051;
wire net9050;
wire net9046;
wire net9989;
wire net9045;
wire net9040;
wire net9039;
wire net9038;
wire net9035;
wire net9032;
wire net9029;
wire net9027;
wire net9026;
wire net9020;
wire net9019;
wire net9018;
wire net9016;
wire net9015;
wire net10504;
wire net9014;
wire net9013;
wire net9011;
wire net9010;
wire net9007;
wire net9005;
wire net9463;
wire net9004;
wire net9003;
wire net9002;
wire net9001;
wire net9000;
wire net8998;
wire net10359;
wire net8997;
wire net8996;
wire net8995;
wire net8993;
wire net8992;
wire net8991;
wire net8989;
wire net8986;
wire net8984;
wire net8983;
wire net8982;
wire net8980;
wire net9475;
wire net8978;
wire net8976;
wire net8975;
wire net8974;
wire net8973;
wire net8972;
wire net10543;
wire net8970;
wire net8969;
wire net8968;
wire net8966;
wire net8965;
wire net8961;
wire net8959;
wire net8958;
wire net8956;
wire net8954;
wire net8953;
wire net8946;
wire net8945;
wire net8941;
wire net8940;
wire net8939;
wire net8937;
wire net10312;
wire net8934;
wire net8927;
wire net9630;
wire net8924;
wire net8921;
wire net9155;
wire net8920;
wire net8919;
wire net8917;
wire net8915;
wire net8913;
wire net8905;
wire net8903;
wire net8902;
wire net8901;
wire net8900;
wire net8899;
wire net8897;
wire net8895;
wire net8893;
wire net8890;
wire net8889;
wire net8887;
wire net8885;
wire net8884;
wire net8882;
wire net9238;
wire net8880;
wire net8877;
wire net8876;
wire net8875;
wire net8873;
wire net8871;
wire net8870;
wire net8869;
wire net8868;
wire net8867;
wire net8865;
wire net8863;
wire net8862;
wire net8861;
wire net8860;
wire net8858;
wire net8857;
wire net8856;
wire net8864;
wire net8855;
wire net8854;
wire net8853;
wire net8852;
wire net8851;
wire net8850;
wire net8849;
wire net8845;
wire net8844;
wire net8838;
wire net8837;
wire net8836;
wire net9055;
wire net8831;
wire net9806;
wire net8827;
wire net8826;
wire net8822;
wire net8821;
wire net8820;
wire net8819;
wire net8816;
wire net10442;
wire net10241;
wire net8814;
wire net8812;
wire net8811;
wire net8810;
wire net8809;
wire net8808;
wire net8806;
wire net8803;
wire net8802;
wire net8799;
wire net8798;
wire net8796;
wire net8795;
wire net10388;
wire net9043;
wire net8791;
wire net8787;
wire net8786;
wire net8785;
wire net8784;
wire net8782;
wire net8780;
wire net8779;
wire net8777;
wire net10081;
wire net8776;
wire net8769;
wire net8768;
wire net8766;
wire net8764;
wire net8763;
wire net9752;
wire net8762;
wire net8761;
wire net8760;
wire net8758;
wire net8753;
wire net8751;
wire net8750;
wire net8749;
wire net8747;
wire net8746;
wire net8745;
wire net8744;
wire net8741;
wire net8740;
wire net8739;
wire net8738;
wire net8737;
wire net8736;
wire net8735;
wire net8733;
wire net8732;
wire net8731;
wire net8728;
wire net10140;
wire net8727;
wire net8726;
wire net10530;
wire net8725;
wire net10178;
wire net8724;
wire net8723;
wire net9828;
wire net8722;
wire net8721;
wire net8720;
wire net8719;
wire net8717;
wire net8715;
wire net8714;
wire net8713;
wire net8712;
wire net8805;
wire net8710;
wire net8708;
wire net8707;
wire net8705;
wire net8704;
wire net8702;
wire net8701;
wire net8699;
wire net8696;
wire net8695;
wire net8693;
wire net8692;
wire net8691;
wire net8689;
wire net8918;
wire net8688;
wire net8686;
wire net8683;
wire net8682;
wire net9490;
wire net8681;
wire net8680;
wire net8678;
wire net8677;
wire net8675;
wire net8673;
wire net8672;
wire net8671;
wire net8669;
wire net8668;
wire net8667;
wire net8666;
wire net8665;
wire net8661;
wire net8660;
wire net10084;
wire net8658;
wire net8653;
wire net8652;
wire net8651;
wire net8648;
wire net8646;
wire net9170;
wire net8644;
wire net8643;
wire net8642;
wire net8641;
wire net8639;
wire net10529;
wire net8638;
wire net8718;
wire net8637;
wire net8636;
wire net8635;
wire net8634;
wire net9192;
wire net8633;
wire net8632;
wire net8631;
wire net8628;
wire net8626;
wire net8625;
wire net8624;
wire net8623;
wire net8621;
wire net8619;
wire net8615;
wire net8874;
wire net8613;
wire net8611;
wire net8981;
wire net8607;
wire net8606;
wire net8605;
wire net8600;
wire net8598;
wire net8597;
wire net8589;
wire net8588;
wire net8587;
wire net10148;
wire net8585;
wire net8584;
wire net8971;
wire net8580;
wire net8579;
wire net8577;
wire net9875;
wire net8576;
wire net8574;
wire net8572;
wire net8571;
wire net8570;
wire net8569;
wire net8568;
wire net8567;
wire net8564;
wire net8560;
wire net8558;
wire net8556;
wire net8555;
wire net8554;
wire net8553;
wire net8552;
wire net9892;
wire net8551;
wire net8911;
wire net8549;
wire net8547;
wire net8546;
wire net8545;
wire net8544;
wire net8929;
wire net8541;
wire net8539;
wire net8538;
wire net8534;
wire net8530;
wire net9371;
wire net8529;
wire net8528;
wire net8527;
wire net10012;
wire net8526;
wire net8525;
wire net8524;
wire net8815;
wire net8521;
wire net10437;
wire net8520;
wire net8519;
wire net8518;
wire net8513;
wire net8512;
wire net10345;
wire net9225;
wire net8510;
wire net8509;
wire net8507;
wire net8498;
wire net8497;
wire net9840;
wire net8495;
wire net8493;
wire net8492;
wire net8489;
wire net8488;
wire net8486;
wire net8480;
wire net8479;
wire net10247;
wire net8478;
wire net8477;
wire net8475;
wire net8474;
wire net8471;
wire net8469;
wire net8468;
wire net8466;
wire net8462;
wire net8460;
wire net8459;
wire net8458;
wire net8456;
wire net8523;
wire net8455;
wire net8454;
wire net8453;
wire net8452;
wire net8450;
wire net8449;
wire net8444;
wire net8442;
wire net8438;
wire net8437;
wire net8434;
wire net8433;
wire net8432;
wire net8429;
wire net8842;
wire net8428;
wire net8427;
wire net8426;
wire net8425;
wire net8423;
wire net8421;
wire net8418;
wire net8417;
wire net8414;
wire net8413;
wire net8412;
wire net8411;
wire net8410;
wire net8409;
wire net8781;
wire net8408;
wire net8407;
wire net8406;
wire net8405;
wire net8404;
wire net8400;
wire net8397;
wire net8396;
wire net8395;
wire net8394;
wire net8391;
wire net8390;
wire net8389;
wire net8388;
wire net8387;
wire net8382;
wire net8381;
wire net8378;
wire net9955;
wire net8377;
wire net8374;
wire net8372;
wire net8371;
wire net8369;
wire net8368;
wire net8367;
wire net8366;
wire net8365;
wire net8363;
wire net8362;
wire net8360;
wire net8358;
wire net8355;
wire net8353;
wire net10237;
wire net8350;
wire net8348;
wire net9522;
wire net8347;
wire net8685;
wire net8345;
wire net9374;
wire net8344;
wire net8343;
wire net8342;
wire net8341;
wire net8339;
wire net9111;
wire net8337;
wire net8335;
wire net8332;
wire net9654;
wire net8331;
wire net8330;
wire net8329;
wire net8328;
wire net8326;
wire net8323;
wire net8322;
wire net8321;
wire net8318;
wire net8317;
wire net8316;
wire net8314;
wire net9030;
wire net8312;
wire net8306;
wire net8304;
wire net8301;
wire net8300;
wire net8297;
wire net8296;
wire net8295;
wire net8292;
wire net8288;
wire net8286;
wire net8284;
wire net8283;
wire net8281;
wire net8280;
wire net8279;
wire net8276;
wire net8273;
wire net8272;
wire net8271;
wire net10230;
wire net8269;
wire net8266;
wire net8265;
wire net8264;
wire net8263;
wire net8261;
wire net9233;
wire net8260;
wire net8357;
wire net8257;
wire net8254;
wire net8253;
wire net8252;
wire out12;
wire net8249;
wire net10036;
wire net8247;
wire out14;
wire net8245;
wire net8244;
wire out22;
wire net8242;
wire net8241;
wire net8240;
wire net8239;
wire net8238;
wire net8236;
wire net8235;
wire net8234;
wire net8232;
wire net8231;
wire net9784;
wire out18;
wire net10177;
wire net8227;
wire net8226;
wire net8225;
wire out11;
wire net8223;
wire net8222;
wire net8220;
wire net8219;
wire net8319;
wire out20;
wire net8218;
wire net8217;
wire net8216;
wire net8213;
wire net8212;
wire net8210;
wire net9279;
wire net8209;
wire out6;
wire net8208;
wire net10386;
wire net8207;
wire net8206;
wire net8205;
wire net8203;
wire net8202;
wire net8201;
wire net8199;
wire net8198;
wire net8754;
wire net8197;
wire net8196;
wire net8195;
wire net8193;
wire net8191;
wire net8190;
wire net8188;
wire net8187;
wire net8186;
wire net8185;
wire net8183;
wire net8179;
wire net8178;
wire net8175;
wire net9187;
wire net8172;
wire net8823;
wire net8168;
wire net8166;
wire net8165;
wire net8164;
wire net8161;
wire net8159;
wire net8158;
wire net9605;
wire net8157;
wire net8156;
wire net8155;
wire net8153;
wire net8516;
wire net8152;
wire net10338;
wire net8150;
wire net8149;
wire net8148;
wire net9713;
wire net8146;
wire net8145;
wire net8144;
wire net8143;
wire net8142;
wire net8140;
wire net8139;
wire net8138;
wire net9493;
wire net8136;
wire net8129;
wire net8128;
wire net8127;
wire net8125;
wire net8124;
wire net8123;
wire net8119;
wire net8118;
wire net8117;
wire net8114;
wire net10194;
wire net8113;
wire net8112;
wire net8448;
wire net8110;
wire net8109;
wire net8106;
wire net8105;
wire net8101;
wire net8100;
wire net8097;
wire net8096;
wire net8095;
wire net8093;
wire net10486;
wire net8092;
wire net9366;
wire net8087;
wire net8084;
wire net9286;
wire net8083;
wire net8082;
wire net9885;
wire net8081;
wire net10200;
wire net8080;
wire net8077;
wire net8076;
wire net9701;
wire net8075;
wire net8074;
wire net8073;
wire net8069;
wire net8068;
wire net8066;
wire net8063;
wire net8062;
wire net8060;
wire net8058;
wire net8057;
wire net8055;
wire net8051;
wire net8050;
wire net8049;
wire net8048;
wire net8047;
wire net8046;
wire net8044;
wire net8043;
wire net8042;
wire net8040;
wire net8039;
wire net8035;
wire net8034;
wire net8032;
wire net10415;
wire net8788;
wire net8030;
wire net8029;
wire net8028;
wire net8027;
wire net8026;
wire net9963;
wire net8025;
wire net8024;
wire net8023;
wire net8021;
wire net8018;
wire net8017;
wire net8016;
wire net8015;
wire net8012;
wire net8011;
wire net8009;
wire net8007;
wire net10355;
wire net8006;
wire net8005;
wire net8004;
wire net8003;
wire net8002;
wire net8001;
wire net7999;
wire net7997;
wire net7996;
wire net10123;
wire net8496;
wire net7994;
wire net7993;
wire net7991;
wire net10387;
wire net7990;
wire net7989;
wire net7988;
wire net7986;
wire net7985;
wire net7983;
wire net7980;
wire net7977;
wire net7974;
wire net7973;
wire net7970;
wire net7960;
wire net7958;
wire net7954;
wire net7953;
wire net7950;
wire net7949;
wire net9322;
wire net7948;
wire net7944;
wire net8305;
wire net7943;
wire net7939;
wire net7937;
wire net7935;
wire net8354;
wire net7934;
wire net7933;
wire net7932;
wire net7930;
wire net7929;
wire net7928;
wire net7926;
wire net7925;
wire net7924;
wire net7923;
wire net7921;
wire net7920;
wire net7919;
wire net7917;
wire net7915;
wire net7914;
wire net7913;
wire net9287;
wire net7912;
wire net7911;
wire net7910;
wire net9666;
wire net7909;
wire net7908;
wire net7906;
wire net7905;
wire net7902;
wire net7892;
wire net7891;
wire net7890;
wire net7889;
wire net7887;
wire net7884;
wire net7881;
wire net7879;
wire net8938;
wire net7878;
wire net7876;
wire net7874;
wire net7873;
wire net7871;
wire net9191;
wire net7870;
wire net7869;
wire out17;
wire net7865;
wire net7864;
wire net7863;
wire net7862;
wire net7861;
wire net8684;
wire net7860;
wire net7857;
wire net8091;
wire net7855;
wire net7852;
wire net7850;
wire net7849;
wire net7848;
wire net7847;
wire net7845;
wire net7843;
wire net7841;
wire net7840;
wire net7836;
wire net7833;
wire net7832;
wire net7824;
wire net7823;
wire net7822;
wire net7816;
wire net7814;
wire net7813;
wire net7812;
wire net7811;
wire net7810;
wire net7809;
wire net7806;
wire net7803;
wire net7802;
wire net7797;
wire net7796;
wire net7795;
wire net7794;
wire net10418;
wire net7791;
wire net7790;
wire net7789;
wire net7787;
wire net7786;
wire net7785;
wire net7781;
wire net7779;
wire net7777;
wire net7776;
wire net7772;
wire net7771;
wire net7770;
wire net7769;
wire net7767;
wire net7765;
wire net9633;
wire net7763;
wire net7762;
wire net7761;
wire net8916;
wire net7760;
wire net7759;
wire net9644;
wire net7758;
wire net7756;
wire net7755;
wire net7754;
wire net7753;
wire net10120;
wire net7752;
wire net7984;
wire net7751;
wire net7749;
wire net7748;
wire net7746;
wire net7745;
wire net7743;
wire net7742;
wire net7740;
wire net7737;
wire net7733;
wire net7732;
wire net7731;
wire net10458;
wire net7730;
wire net7729;
wire net7726;
wire net7725;
wire net7724;
wire net7723;
wire net7721;
wire net7719;
wire net7715;
wire net7714;
wire net7712;
wire net7711;
wire net7710;
wire net7708;
wire net7707;
wire net7706;
wire net7704;
wire net7703;
wire net7699;
wire net9851;
wire net7696;
wire net7694;
wire net7693;
wire net7691;
wire net7688;
wire net7687;
wire net7686;
wire net7679;
wire net7678;
wire net7784;
wire net7675;
wire net7674;
wire net7671;
wire net7670;
wire net7669;
wire net7668;
wire net7666;
wire net7665;
wire net7663;
wire net7662;
wire net7660;
wire net7659;
wire net10470;
wire net7656;
wire net7655;
wire net7654;
wire net7653;
wire net7652;
wire net7651;
wire net8988;
wire net7648;
wire net9260;
wire net7647;
wire net7645;
wire net7644;
wire net7643;
wire net7642;
wire net8550;
wire net7641;
wire net7640;
wire net7636;
wire net7634;
wire net7633;
wire net7632;
wire net7631;
wire net7629;
wire net10480;
wire net7628;
wire net7627;
wire net7626;
wire net7625;
wire net7624;
wire net10143;
wire net7621;
wire net7619;
wire net7617;
wire net7615;
wire net7614;
wire net9025;
wire net7609;
wire net7607;
wire net7605;
wire net8752;
wire net7603;
wire net7601;
wire net7600;
wire net7598;
wire net7595;
wire net7594;
wire net7593;
wire net7592;
wire net7591;
wire net9771;
wire net7590;
wire net8385;
wire net7588;
wire net7587;
wire net7586;
wire net7585;
wire net7584;
wire net7582;
wire net7581;
wire net7579;
wire net9335;
wire net7577;
wire net7572;
wire net9113;
wire net7571;
wire net7570;
wire net7569;
wire net7568;
wire net7566;
wire net7565;
wire net7564;
wire net7562;
wire net7561;
wire net7560;
wire net7559;
wire net8131;
wire net7558;
wire net7556;
wire net9705;
wire net7554;
wire net7553;
wire net7549;
wire net9717;
wire net7547;
wire net7546;
wire net7545;
wire net7543;
wire net7541;
wire net7540;
wire net7539;
wire net9586;
wire net7538;
wire net7537;
wire net7956;
wire net7536;
wire net7535;
wire net7533;
wire net7531;
wire net7530;
wire net7529;
wire net7527;
wire net9611;
wire net7526;
wire net7525;
wire net7523;
wire net7522;
wire net7521;
wire net7520;
wire net7519;
wire net9669;
wire net7518;
wire net7517;
wire net7516;
wire net7514;
wire net7510;
wire net7509;
wire net8102;
wire net7508;
wire net7507;
wire net7505;
wire net7503;
wire net7502;
wire net7501;
wire net7500;
wire net10147;
wire net8979;
wire net7499;
wire net7498;
wire net7657;
wire net7497;
wire net7493;
wire net10488;
wire net7489;
wire net7488;
wire net7486;
wire net7484;
wire net3712;
wire net3650;
wire net5066;
wire net5427;
wire net3699;
wire net4859;
wire net3697;
wire net7427;
wire net3692;
wire net3687;
wire net3684;
wire net4757;
wire net3678;
wire net3673;
wire net2661;
wire net3672;
wire net4673;
wire net8338;
wire net5036;
wire net1050;
wire net3670;
wire net9022;
wire net3669;
wire net6666;
wire net3662;
wire net3657;
wire net10570;
wire net4219;
wire net8888;
wire net5980;
wire net7194;
wire net6390;
wire net3648;
wire net3641;
wire net1859;
wire net3637;
wire net4378;
wire net3635;
wire net8103;
wire net3622;
wire net324;
wire net3615;
wire net3609;
wire net649;
wire net6312;
wire net9079;
wire net3601;
wire net3597;
wire net3596;
wire net3590;
wire net3695;
wire net7859;
wire net4122;
wire net3588;
wire net3390;
wire net2119;
wire net3584;
wire net60;
wire net3582;
wire net3578;
wire net3575;
wire net3574;
wire net3570;
wire net4709;
wire net3567;
wire net3559;
wire net2665;
wire net3557;
wire net3556;
wire net1002;
wire net4495;
wire net3129;
wire net377;
wire net3548;
wire net8832;
wire net3660;
wire net5247;
wire net3546;
wire net2380;
wire net3545;
wire net9569;
wire net8104;
wire net3544;
wire net8593;
wire net6638;
wire net3543;
wire net7268;
wire net9933;
wire net3539;
wire net3538;
wire net3536;
wire net4159;
wire net8346;
wire net3535;
wire net3529;
wire net2047;
wire net3525;
wire net7410;
wire net3523;
wire net3521;
wire net5119;
wire net3517;
wire net7271;
wire net7931;
wire net3512;
wire net3175;
wire net9138;
wire net3511;
wire net3509;
wire net4564;
wire net6676;
wire net3508;
wire net3507;
wire net9740;
wire net3502;
wire net3500;
wire net3494;
wire net919;
wire net7196;
wire net8470;
wire net3493;
wire net5719;
wire net3491;
wire net3489;
wire net10007;
wire net329;
wire net3488;
wire net8908;
wire net7311;
wire net3487;
wire net3532;
wire net3486;
wire net3485;
wire net3484;
wire net3480;
wire net4321;
wire net3478;
wire net3476;
wire net2043;
wire net9033;
wire net3473;
wire net571;
wire net3469;
wire net3466;
wire net3455;
wire net3451;
wire net8303;
wire net3260;
wire net3649;
wire net3449;
wire net5042;
wire net8022;
wire net5709;
wire net3444;
wire net2461;
wire net3442;
wire net3440;
wire net3439;
wire net144;
wire net3519;
wire net872;
wire net5099;
wire net6791;
wire net3426;
wire net8603;
wire net2003;
wire net6715;
wire net3427;
wire net3542;
wire net9328;
wire net3423;
wire net3419;
wire net4987;
wire net3688;
wire net171;
wire net4354;
wire net3638;
wire net8536;
wire net3411;
wire net2884;
wire net3410;
wire net3408;
wire net1343;
wire net10555;
wire net10350;
wire net6850;
wire net3547;
wire net3406;
wire net8189;
wire net135;
wire net3401;
wire net7616;
wire net3396;
wire net3210;
wire net3394;
wire net3387;
wire net5745;
wire net3384;
wire net3382;
wire net3380;
wire net3377;
wire net7513;
wire net6701;
wire net9292;
wire net3376;
wire net3366;
wire net3370;
wire net7428;
wire net3369;
wire net7485;
wire net3368;
wire net9124;
wire net3367;
wire net3363;
wire net1951;
wire net7285;
wire net9115;
wire net3360;
wire net621;
wire net5422;
wire net3354;
wire net1870;
wire net3350;
wire net3345;
wire net5930;
wire net9854;
wire net4533;
wire net3634;
wire net3341;
wire net7183;
wire net3339;
wire net5845;
wire net3336;
wire net354;
wire net3330;
wire net3327;
wire net1054;
wire net10212;
wire net6551;
wire net3326;
wire net3325;
wire net9148;
wire net3323;
wire net5533;
wire net3318;
wire net7804;
wire net4881;
wire net3316;
wire net1321;
wire net3314;
wire net1702;
wire net3302;
wire net3294;
wire net9273;
wire net3288;
wire net3286;
wire net3284;
wire net581;
wire net7415;
wire net3921;
wire net3280;
wire net2894;
wire net3589;
wire net3691;
wire net5590;
wire net8038;
wire net3278;
wire net2687;
wire net3277;
wire net3275;
wire net4097;
wire net9541;
wire net3658;
wire net10499;
wire net3257;
wire net2284;
wire net7220;
wire net3252;
wire net3246;
wire net3234;
wire net3240;
wire net3239;
wire net5808;
wire net7269;
wire in24;
wire net4645;
wire net7416;
wire net3235;
wire net6464;
wire net3232;
wire net3230;
wire net532;
wire net5925;
wire net3228;
wire net3149;
wire net3227;
wire net5044;
wire net3225;
wire net3224;
wire net3438;
wire net7695;
wire net1451;
wire net8793;
wire net3219;
wire net3218;
wire net5214;
wire net5183;
wire net3211;
wire net3352;
wire net8336;
wire net5697;
wire net7075;
wire net3207;
wire net2852;
wire net9919;
wire net7286;
wire net3198;
wire net3193;
wire net6500;
wire net3191;
wire net3186;
wire net3184;
wire net4949;
wire net3180;
wire net7267;
wire net3647;
wire net3177;
wire net3173;
wire net7727;
wire net3169;
wire net9972;
wire net9810;
wire net1060;
wire net3165;
wire net3498;
wire net3157;
wire net8833;
wire net3375;
wire net8472;
wire net147;
wire net3145;
wire net3143;
wire net3141;
wire net3140;
wire net3137;
wire net3134;
wire net3130;
wire net3126;
wire net8771;
wire net2091;
wire net533;
wire net5789;
wire net6923;
wire net7018;
wire net3160;
wire net6275;
wire net3121;
wire net1918;
wire net3112;
wire net126;
wire net3111;
wire net8663;
wire net7511;
wire net3067;
wire net2981;
wire net8839;
wire net3110;
wire net5123;
wire net3109;
wire net3102;
wire net224;
wire net836;
wire net5999;
wire net5375;
wire net3097;
wire net9684;
wire net3321;
wire net3096;
wire net8542;
wire net8464;
wire net749;
wire net2783;
wire net7998;
wire net3459;
wire net5815;
wire net7006;
wire net3088;
wire net7242;
wire net7567;
wire net3125;
wire net3526;
wire net7927;
wire net5683;
wire net3085;
wire net1175;
wire net2560;
wire net3083;
wire net8215;
wire net2435;
wire net3808;
wire net3698;
wire net3082;
wire net3081;
wire net2565;
wire net3076;
wire net3215;
wire net7151;
wire net3071;
wire net9382;
wire net3949;
wire net3070;
wire net3068;
wire net4842;
wire net6767;
wire net3600;
wire net7306;
wire net3058;
wire net2138;
wire net3057;
wire net2211;
wire net9129;
wire net574;
wire net3431;
wire net3055;
wire net3492;
wire net3053;
wire net5876;
wire net3049;
wire net3047;
wire net8532;
wire net7244;
wire net9217;
wire net3042;
wire net3039;
wire net6528;
wire net9214;
wire net3036;
wire net3035;
wire net3099;
wire net1258;
wire net3034;
wire net3032;
wire net3030;
wire net10023;
wire net7524;
wire net1080;
wire net3029;
wire net10308;
wire net3028;
wire net3023;
wire net2962;
wire net3021;
wire net3017;
wire net1663;
wire net3016;
wire net9355;
wire net5554;
wire net8932;
wire net3015;
wire net847;
wire net3014;
wire net4414;
wire net9450;
wire net3011;
wire net3077;
wire net3010;
wire net5794;
wire net8649;
wire net3006;
wire net411;
wire net10372;
wire net6852;
wire net3005;
wire net3004;
wire net3003;
wire net1704;
wire net9064;
wire net3002;
wire net3000;
wire net2996;
wire net3158;
wire net7131;
wire net1525;
wire net916;
wire net2989;
wire net9767;
wire net3187;
wire net2022;
wire net5200;
wire net6740;
wire net1830;
wire net6770;
wire net6251;
wire net2979;
wire net2978;
wire net159;
wire net2975;
wire net2972;
wire net2730;
wire net326;
wire net10263;
wire net6700;
wire net7684;
wire net2971;
wire net4955;
wire net3562;
wire net4191;
wire net2969;
wire net3481;
wire net2968;
wire net2967;
wire net1022;
wire net287;
wire net3059;
wire net3118;
wire net7176;
wire net2954;
wire net2863;
wire net10360;
wire net9247;
wire net2509;
wire net6044;
wire net2950;
wire net2058;
wire net5520;
wire net3458;
wire net2949;
wire net792;
wire net2946;
wire net2714;
wire net2681;
wire net6721;
wire net2941;
wire net2940;
wire net8251;
wire net2939;
wire net2938;
wire net2936;
wire net7894;
wire net753;
wire net2932;
wire net2930;
wire net6782;
wire net6858;
wire net2928;
wire net9245;
wire net5767;
wire net2923;
wire net2921;
wire net2918;
wire net2917;
wire net2915;
wire net1442;
wire net3679;
wire net6584;
wire net2913;
wire net3859;
wire net7155;
wire net5225;
wire net8964;
wire net4032;
wire net2908;
wire net4094;
wire net2903;
wire net4135;
wire net2902;
wire net9122;
wire net2436;
wire net5492;
wire net7918;
wire net4096;
wire net5265;
wire net534;
wire net10421;
wire net3616;
wire net3533;
wire net2891;
wire net6354;
wire net2886;
wire net5222;
wire net1664;
wire net2878;
wire net2195;
wire net1705;
wire net2877;
wire net8923;
wire net8514;
wire net6667;
wire net6895;
wire net2875;
wire net1256;
wire net3074;
wire net2872;
wire net7250;
wire net10032;
wire net2870;
wire net4238;
wire net2869;
wire net4437;
wire net4475;
wire net4560;
wire net2595;
wire net8610;
wire net2516;
wire net1992;
wire net9085;
wire net6657;
wire net2847;
wire net461;
wire net6897;
wire net2836;
wire net35;
wire net5199;
wire net4652;
wire net5548;
wire net2988;
wire net2871;
wire net2834;
wire net8262;
wire net2832;
wire net2831;
wire net4978;
wire net7309;
wire net2829;
wire net3447;
wire net2752;
wire net9097;
wire net5368;
wire net2826;
wire net2818;
wire net3714;
wire net6357;
wire net2817;
wire net4128;
wire net7971;
wire net2811;
wire net3116;
wire net2807;
wire net5561;
wire net7900;
wire net5735;
wire net2806;
wire net6496;
wire net3467;
wire net8494;
wire net2705;
wire net2801;
wire net2800;
wire net5443;
wire net9203;
wire net2798;
wire net2796;
wire net9813;
wire net3655;
wire net2793;
wire net9567;
wire net3342;
wire net7107;
wire net2790;
wire net8379;
wire net1631;
wire net3710;
wire net1568;
wire net4512;
wire net3995;
wire net3133;
wire net7310;
wire net2784;
wire net2781;
wire net8907;
wire net3831;
wire net4138;
wire net2402;
wire net2777;
wire net3162;
wire net2145;
wire net9270;
wire net146;
wire net2952;
wire net802;
wire net2767;
wire net2766;
wire net5588;
wire net3306;
wire net9639;
wire net6689;
wire net9577;
wire net6806;
wire net2763;
wire net945;
wire net4085;
wire net5372;
wire net5432;
wire net2758;
wire net2756;
wire net2749;
wire net923;
wire net3961;
wire net2747;
wire net9465;
wire net9267;
wire net690;
wire net3203;
wire net9249;
wire net1601;
wire net2743;
wire net3950;
wire net6240;
wire net5193;
wire net6601;
wire net2742;
wire net4666;
wire net8620;
wire net5801;
wire net6272;
wire net3388;
wire net2368;
wire net3528;
wire net585;
wire net3212;
wire net5397;
wire net2738;
wire net2495;
wire net1173;
wire net4323;
wire net7324;
wire net2733;
wire net6028;
wire net7701;
wire net2000;
wire net3276;
wire net7372;
wire net2723;
wire net8912;
wire net2722;
wire net2720;
wire net10573;
wire net1215;
wire net5480;
wire net2707;
wire net5675;
wire net6569;
wire net2700;
wire net777;
wire net3980;
wire net2694;
wire net3516;
wire net1508;
wire net9965;
wire net2622;
wire net7354;
wire net1197;
wire net2691;
wire net2689;
wire out4;
wire net795;
wire net2684;
wire net10196;
wire net8508;
wire net2680;
wire net3348;
wire net2497;
wire net2679;
wire net2674;
wire net1459;
wire net2873;
wire net2760;
wire net2666;
wire net10034;
wire net3612;
wire net3221;
wire net5313;
wire net2663;
wire net3811;
wire net9426;
wire net105;
wire net2659;
wire net2658;
wire net10026;
wire net407;
wire net3268;
wire net4808;
wire net2657;
wire net2653;
wire net2381;
wire net2652;
wire net2650;
wire net1934;
wire net2649;
wire net9023;
wire net2648;
wire net1786;
wire net1037;
wire net2791;
wire net2642;
wire net454;
wire net4528;
wire net2634;
wire net4608;
wire net2631;
wire net2626;
wire net2772;
wire net2625;
wire net6280;
wire net6302;
wire net3202;
wire net4113;
wire net10351;
wire net6979;
wire net4964;
wire net9620;
wire net2620;
wire net9745;
wire net3199;
wire net2618;
wire net626;
wire net6673;
wire net1800;
wire net3346;
wire net231;
wire net3251;
wire net3964;
wire net7034;
wire net9446;
wire net6600;
wire net9137;
wire net2782;
wire net2610;
wire net2603;
wire net361;
wire net4086;
wire net2601;
wire net2600;
wire net662;
wire net8778;
wire net2596;
wire net3802;
wire net2591;
wire net9530;
wire net276;
wire net8828;
wire net2588;
wire net4819;
wire net2586;
wire net2014;
wire net9451;
wire net2232;
wire net2375;
wire net6123;
wire net2583;
wire net2581;
wire net3775;
wire in17;
wire net9990;
wire net4650;
wire net2579;
wire net2695;
wire net5839;
wire net7961;
wire net3579;
wire net2960;
wire net2576;
wire net2574;
wire net9799;
wire net6922;
wire net2571;
wire net2569;
wire net9491;
wire net3031;
wire net2568;
wire net1575;
wire net7799;
wire net3153;
wire net10540;
wire net2655;
wire net4907;
wire net8765;
wire net7623;
wire net6843;
wire net2566;
wire net2563;
wire net5332;
wire net2561;
wire net6644;
wire net7476;
wire net2557;
wire net2555;
wire net1597;
wire net6793;
wire net2543;
wire net2672;
wire net2542;
wire net2541;
wire net1241;
wire net7612;
wire net5883;
wire net2538;
wire net1544;
wire net5457;
wire net8325;
wire net2536;
wire net7801;
wire net5933;
wire net2535;
wire net1563;
wire net5098;
wire net10405;
wire net2534;
wire net2532;
wire net2208;
wire net2527;
wire net9904;
wire net1688;
wire net7965;
wire net3624;
wire net7898;
wire net2524;
wire net8891;
wire net4747;
wire net6618;
wire net6545;
wire net2521;
wire net2520;
wire net4532;
wire net2519;
wire net2518;
wire net2241;
wire net2517;
wire net3586;
wire net2504;
wire net3247;
wire net1203;
wire net2502;
wire net2500;
wire net2499;
wire net3581;
wire net8543;
wire net3392;
wire net5312;
wire net2491;
wire net2487;
wire net2482;
wire net2956;
wire net5093;
wire net9733;
wire net3560;
wire net6660;
wire net5692;
wire net6542;
wire net2480;
wire net2479;
wire net2478;
wire net7750;
wire net2476;
wire net1592;
wire net8987;
wire net65;
wire net2645;
wire net5245;
wire net1613;
wire net5690;
wire net6619;
wire net5238;
wire net9687;
wire net8485;
wire net2469;
wire net2115;
wire net2896;
wire net734;
wire net2460;
wire net2459;
wire net7302;
wire net2453;
wire net2452;
wire net5022;
wire net2448;
wire net1460;
wire net2660;
wire net8711;
wire net2444;
wire net7938;
wire net2442;
wire net2233;
wire net2440;
wire net2439;
wire net8935;
wire net2438;
wire net3470;
wire net2842;
wire net2951;
wire net2498;
wire net2033;
wire net2431;
wire net8457;
wire net1888;
wire net8948;
wire net870;
wire net2429;
wire net6532;
wire net2810;
wire net4108;
wire net2425;
wire net2424;
wire net2422;
wire net8825;
wire net4444;
wire net3155;
wire net208;
wire net4180;
wire net8614;
wire net2421;
wire net604;
wire net3300;
wire net178;
wire net6745;
wire net2416;
wire net2525;
wire net5067;
wire net2413;
wire net1446;
wire net2412;
wire net2411;
wire net7182;
wire net2408;
wire net7972;
wire net2407;
wire net1914;
wire net912;
wire net2404;
wire net2401;
wire net2400;
wire net4607;
wire net6249;
wire net2399;
wire net2397;
wire net2391;
wire net1477;
wire net2390;
wire net10055;
wire net2389;
wire net2388;
wire net6522;
wire net2386;
wire net2385;
wire net10294;
wire net5806;
wire net1181;
wire net2379;
wire net2378;
wire net1848;
wire net2377;
wire net3619;
wire net2840;
wire net2271;
wire net1611;
wire net7895;
wire net6720;
wire net2370;
wire net2364;
wire net8578;
wire net1520;
wire net10417;
wire net2362;
wire net4204;
wire net2361;
wire net3850;
wire net7431;
wire net2356;
wire net2353;
wire net2724;
wire net10508;
wire net3803;
wire net2352;
wire net3148;
wire net1139;
wire net10223;
wire net2351;
wire net9104;
wire net6705;
wire net9714;
wire net2349;
wire net7085;
wire net8293;
wire net2718;
wire net8501;
wire net2347;
wire net2383;
wire net2345;
wire net2858;
wire net2344;
wire net2343;
wire net4250;
wire net8756;
wire net7387;
wire net2338;
wire net5430;
wire net2335;
wire net2334;
wire net9368;
wire net3163;
wire net9425;
wire net2006;
wire net1463;
wire net8465;
wire net3541;
wire net8033;
wire net7738;
wire net7281;
wire net9782;
wire net2326;
wire net9041;
wire net2325;
wire net2317;
wire net5091;
wire net1747;
wire net10289;
wire net8990;
wire net8169;
wire net138;
wire net365;
wire net2312;
wire net9060;
wire net2309;
wire net3413;
wire net7009;
wire net1640;
wire net3668;
wire net4457;
wire net2302;
wire net1118;
wire net390;
wire net2528;
wire net2296;
wire net10302;
wire net1738;
wire net1030;
wire net10507;
wire net2292;
wire net10261;
wire net3124;
wire net2291;
wire net6097;
wire net2290;
wire net762;
wire net5890;
wire net6968;
wire net2307;
wire net6281;
wire net2287;
wire net8361;
wire net5202;
wire net9096;
wire net1909;
wire net3885;
wire net133;
wire net216;
wire net1261;
wire net7417;
wire net2716;
wire net2280;
wire net2846;
wire net2279;
wire net2426;
wire net164;
wire net8067;
wire net2830;
wire net2275;
wire net4011;
wire net2274;
wire net2719;
wire net3269;
wire net5030;
wire net3623;
wire net2276;
wire net2272;
wire net3305;
wire net6714;
wire net2269;
wire net1596;
wire net2735;
wire net3307;
wire net2263;
wire net5075;
wire net5670;
wire net2904;
wire net4118;
wire net2262;
wire net2259;
wire net7193;
wire net2252;
wire net2251;
wire net2249;
wire net5984;
wire net2248;
wire net4790;
wire net2247;
wire net1116;
wire net2245;
wire net2765;
wire net2244;
wire net2243;
wire net6625;
wire net2242;
wire net2240;
wire net3295;
wire net1713;
wire net2238;
wire net2237;
wire net7221;
wire net8789;
wire net179;
wire net1571;
wire net2230;
wire net2229;
wire net8930;
wire net4272;
wire net2277;
wire net7690;
wire net5572;
wire net3066;
wire net5626;
wire net3554;
wire net2226;
wire net4116;
wire net5499;
wire net3310;
wire net2224;
wire net10476;
wire net2222;
wire net1865;
wire net6178;
wire net2219;
wire net10483;
wire net8504;
wire net2313;
wire net4206;
wire net1822;
wire net6485;
wire net1975;
wire net2204;
wire net3527;
wire net4196;
wire net5105;
wire net2192;
wire net2191;
wire net2187;
wire net4006;
wire net2184;
wire net5908;
wire net7483;
wire net2182;
wire net2741;
wire net7975;
wire net327;
wire net9065;
wire net3103;
wire net3291;
wire net4844;
wire net2174;
wire net2172;
wire net3836;
wire net7300;
wire net10198;
wire net3522;
wire net2171;
wire net2165;
wire net2164;
wire net2163;
wire net4775;
wire net2162;
wire net5017;
wire net2161;
wire net1340;
wire net9274;
wire net5607;
wire net6579;
wire net2160;
wire net1208;
wire net9312;
wire net2157;
wire in5;
wire net396;
wire net2154;
wire net7899;
wire net7231;
wire net7184;
wire net2152;
wire net2151;
wire net3890;
wire net2149;
wire net2144;
wire net10357;
wire net7358;
wire net9482;
wire net2493;
wire net6435;
wire net2142;
wire net9554;
wire net8370;
wire net6595;
wire net2135;
wire net2134;
wire net9017;
wire net7551;
wire net853;
wire net8461;
wire net3250;
wire net5382;
wire net8645;
wire net8467;
wire net2354;
wire net2822;
wire net2693;
wire net8403;
wire net5638;
wire net2137;
wire net3643;
wire net2129;
wire net4315;
wire net10158;
wire net9890;
wire net3120;
wire net2126;
wire net5891;
wire net2125;
wire net3436;
wire net1876;
wire net1741;
wire net2123;
wire net219;
wire net2120;
wire net3752;
wire net794;
wire net4363;
wire net1069;
wire net8957;
wire net1365;
wire net6606;
wire net7866;
wire net2114;
wire net2113;
wire net2111;
wire net2108;
wire net2106;
wire net2710;
wire net343;
wire net2105;
wire net8120;
wire net2270;
wire net1809;
wire net10556;
wire net2102;
wire net292;
wire net2881;
wire net3496;
wire net9994;
wire net2101;
wire net2959;
wire net2097;
wire net2708;
wire net2096;
wire net330;
wire net1219;
wire net5507;
wire net2474;
wire net2094;
wire net9557;
wire net6868;
wire net9956;
wire net2088;
wire net2086;
wire net8380;
wire net3267;
wire net8960;
wire net2508;
wire net10500;
wire net2085;
wire net2215;
wire net6537;
wire net2570;
wire net655;
wire net2084;
wire net2041;
wire net503;
wire net2078;
wire net6248;
wire net2180;
wire net3989;
wire net9523;
wire net8730;
wire net6946;
wire net3237;
wire net2073;
wire net2393;
wire net2072;
wire net2970;
wire net2068;
wire net2064;
wire net5702;
wire net9929;
wire net212;
wire net2061;
wire net9034;
wire net7853;
wire net2060;
wire net4319;
wire net9520;
wire net3308;
wire net2057;
wire net3626;
wire net8627;
wire net2054;
wire net425;
wire net3381;
wire net2769;
wire net1796;
wire net2010;
wire net4329;
wire net2859;
wire net2048;
wire net515;
wire net2045;
wire net2265;
wire net6350;
wire net6908;
wire net2042;
wire net7969;
wire net2039;
wire net2037;
wire net1958;
wire net2032;
wire net2246;
wire net1155;
wire net1429;
wire net7716;
wire net2026;
wire net1170;
wire net4754;
wire net2023;
wire net2725;
wire net177;
wire net2021;
wire net10100;
wire net2210;
wire net1368;
wire net7968;
wire net4415;
wire net6395;
wire net10076;
wire net7867;
wire net2019;
wire net6594;
wire net2018;
wire net2016;
wire net2332;
wire net211;
wire net6226;
wire net2015;
wire net2776;
wire net8445;
wire net7359;
wire net2007;
wire net9162;
wire net2005;
wire net3248;
wire net2001;
wire net430;
wire net2098;
wire net1998;
wire net1997;
wire net1853;
wire net750;
wire net5278;
wire net2948;
wire net6708;
wire net1994;
wire net3762;
wire net6194;
wire net2040;
wire net1993;
wire net2009;
wire net310;
wire net10150;
wire net8311;
wire net6727;
wire net2506;
wire net1991;
wire net6892;
wire net2104;
wire net763;
wire net3738;
wire net1190;
wire net1989;
wire net6776;
wire net4922;
wire net3080;
wire net1985;
wire net8392;
wire net744;
wire net9941;
wire net1984;
wire net350;
wire net3726;
wire net8951;
wire net4254;
wire net1983;
wire net1291;
wire net3955;
wire net1977;
wire net1308;
wire net1974;
wire net1754;
wire net4034;
wire net8174;
wire net255;
wire net2792;
wire net5576;
wire net2255;
wire net2572;
wire net1466;
wire net2890;
wire net3967;
wire net2505;
wire net5367;
wire net5369;
wire net1967;
wire net1964;
wire net2985;
wire net1961;
wire net2845;
wire net1960;
wire net9481;
wire net6332;
wire net1959;
wire net1956;
wire net2197;
wire net2471;
wire net3416;
wire net6025;
wire net10278;
wire net9173;
wire net2974;
wire net4137;
wire net1948;
wire net1946;
wire net2510;
wire net1945;
wire net2567;
wire net1943;
wire net1942;
wire net1940;
wire net1939;
wire net6218;
wire net9624;
wire net8447;
wire net2841;
wire net1937;
wire net4937;
wire net861;
wire net9036;
wire net3338;
wire net2823;
wire net2545;
wire net1931;
wire net5031;
wire net9417;
wire net6115;
wire net8134;
wire net5493;
wire net6598;
wire net1923;
wire net1922;
wire net970;
wire net1921;
wire net9485;
wire net5558;
wire net6316;
wire net2214;
wire net1913;
wire net1912;
wire net7378;
wire net4812;
wire net1767;
wire net2933;
wire net8654;
wire net2888;
wire net1903;
wire net8925;
wire net1899;
wire net1897;
wire net8327;
wire net999;
wire net6429;
wire net1896;
wire net3705;
wire net1555;
wire net4107;
wire net1895;
wire net3090;
wire net1894;
wire net10052;
wire net1889;
wire net6166;
wire net2257;
wire net7606;
wire net7259;
wire net3337;
wire net2585;
wire net1293;
wire net8608;
wire net3279;
wire net2036;
wire net1887;
wire net10399;
wire net4647;
wire net2398;
wire net1884;
wire net1883;
wire net294;
wire net5749;
wire net1864;
wire net1861;
wire net500;
wire net1857;
wire net1856;
wire net1855;
wire net172;
wire net9028;
wire net4174;
wire net3681;
wire net1854;
wire net2599;
wire net1850;
wire net4570;
wire net4948;
wire net2337;
wire net1849;
wire net10393;
wire net10206;
wire net686;
wire net7290;
wire net3371;
wire net1846;
wire net904;
wire net442;
wire net10319;
wire net5192;
wire net1842;
wire net1841;
wire net3209;
wire net4044;
wire net1908;
wire net1840;
wire net6462;
wire net1838;
wire net7573;
wire net1851;
wire net1837;
wire net2503;
wire net5678;
wire net6907;
wire net8994;
wire net1835;
wire net8773;
wire net4422;
wire net1826;
wire net6058;
wire net1556;
wire net5253;
wire net5612;
wire net10281;
wire net1819;
wire net1817;
wire net3530;
wire net340;
wire net3194;
wire net1813;
wire net3652;
wire net3378;
wire net3084;
wire net1501;
wire net5756;
wire net2261;
wire net3242;
wire net4839;
wire net2110;
wire net1029;
wire net4802;
wire net3884;
wire net4846;
wire net1811;
wire net313;
wire net4172;
wire net3317;
wire net2076;
wire net1806;
wire net5508;
wire net2628;
wire net776;
wire net10491;
wire net2740;
wire net2575;
wire net1802;
wire net5989;
wire net10197;
wire net6467;
wire net3349;
wire net9497;
wire net2494;
wire net1795;
wire net1318;
wire net6297;
wire net2305;
wire net1792;
wire net9409;
wire net8430;
wire net977;
wire net1791;
wire net2761;
wire net4700;
wire net335;
wire net9367;
wire net6934;
wire net4229;
wire net5823;
wire net5924;
wire net3105;
wire net5556;
wire net7922;
wire net4684;
wire net4863;
wire net7955;
wire net6555;
wire net2704;
wire net9787;
wire net6159;
wire net8151;
wire net1780;
wire net1775;
wire net6976;
wire net3593;
wire net3195;
wire net1654;
wire net1774;
wire net9636;
wire net3503;
wire net2754;
wire net1987;
wire net5674;
wire net1771;
wire net7335;
wire net1770;
wire net3362;
wire net1769;
wire net5172;
wire net1768;
wire net8830;
wire net6197;
wire net6960;
wire net8356;
wire net1766;
wire net9800;
wire net1763;
wire net10452;
wire net2816;
wire net2329;
wire net1759;
wire net9143;
wire net4236;
wire net1757;
wire net2481;
wire net2874;
wire net2753;
wire net3233;
wire net1749;
wire net7374;
wire net5621;
wire net4618;
wire net6531;
wire net2295;
wire net1372;
wire net8170;
wire net114;
wire net8111;
wire net5914;
wire net1742;
wire net5768;
wire net1739;
wire net6451;
wire net4815;
wire net9517;
wire net6574;
wire net3462;
wire net1734;
wire net1733;
wire net2640;
wire net1732;
wire net483;
wire net7916;
wire net1731;
wire net6664;
wire net5288;
wire net1730;
wire net8840;
wire net4280;
wire net4813;
wire net1729;
wire net2731;
wire net1726;
wire net5147;
wire net1725;
wire net4803;
wire net1724;
wire net9942;
wire net5446;
wire net9494;
wire net1723;
wire net116;
wire net28;
wire net1722;
wire net22;
wire net6838;
wire net7744;
wire net1721;
wire net9272;
wire net8602;
wire net8086;
wire net2892;
wire net1720;
wire net1716;
wire net578;
wire net1179;
wire net8070;
wire net5858;
wire net5816;
wire net1040;
wire net3220;
wire net246;
wire net783;
wire net1828;
wire net43;
wire net541;
wire net6604;
wire net4828;
wire net3693;
wire net3037;
wire net8107;
wire net2253;
wire net1941;
wire net6651;
wire net772;
wire net7059;
wire net2643;
wire net761;
wire net8952;
wire net478;
wire net15;
wire net8383;
wire net4301;
wire net9397;
wire net5025;
wire net746;
wire net168;
wire net2827;
wire net6160;
wire net738;
wire net1938;
wire net5560;
wire net3204;
wire net9435;
wire net9285;
wire net1638;
wire net737;
wire net1125;
wire net2879;
wire net3293;
wire net5458;
wire net4904;
wire net7327;
wire net9993;
wire net736;
wire net1785;
wire net414;
wire net5344;
wire net1122;
wire net2696;
wire net7078;
wire net2559;
wire net7462;
wire net730;
wire net4917;
wire net3146;
wire net728;
wire net3599;
wire net406;
wire net9396;
wire net5624;
wire net1999;
wire net4156;
wire net725;
wire net4517;
wire net808;
wire net2732;
wire net2392;
wire net724;
wire net6546;
wire net1526;
wire net2787;
wire net2220;
wire net721;
wire net9889;
wire net7315;
wire net3632;
wire net7661;
wire net1315;
wire net1814;
wire net797;
wire net7548;
wire net1502;
wire net4756;
wire net1475;
wire net715;
wire net1100;
wire net1689;
wire net4316;
wire net9461;
wire net1178;
wire net4708;
wire net3046;
wire net703;
wire net1519;
wire net679;
wire net9550;
wire net1265;
wire net9928;
wire net3552;
wire net700;
wire net4170;
wire net3666;
wire net699;
wire net1075;
wire net706;
wire net4789;
wire net596;
wire net25;
wire net691;
wire net1488;
wire net5351;
wire net2906;
wire net10037;
wire net676;
wire net3078;
wire net7683;
wire net2258;
wire net6107;
wire net1051;
wire net960;
wire net8894;
wire net8274;
wire net2887;
wire net6641;
wire net693;
wire net2515;
wire net914;
wire net1264;
wire net7379;
wire net2446;
wire net670;
wire net7672;
wire net397;
wire net5387;
wire net7054;
wire net6940;
wire net2668;
wire net1218;
wire net6954;
wire net1656;
wire net4962;
wire net1660;
wire net1773;
wire net648;
wire net842;
wire net153;
wire net644;
wire net1418;
wire net5248;
wire net3008;
wire net1373;
wire net640;
wire net4841;
wire net1827;
wire net5348;
wire net5070;
wire net3389;
wire net1797;
wire net282;
wire net6311;
wire net10541;
wire net7166;
wire net637;
wire net2692;
wire net3977;
wire net2038;
wire net1947;
wire net7261;
wire net238;
wire net1383;
wire net7349;
wire net3024;
wire net579;
wire net2604;
wire net713;
wire net4766;
wire net2083;
wire net707;
wire net559;
wire net5884;
wire net632;
wire net8299;
wire net770;
wire net8949;
wire net2188;
wire net3409;
wire net1331;
wire net4499;
wire net2578;
wire net2651;
wire net631;
wire net611;
wire net9793;
wire net4899;
wire net1146;
wire net617;
wire net986;
wire net1615;
wire net6368;
wire net6816;
wire net7109;
wire net817;
wire net4176;
wire net3504;
wire net3355;
wire net2409;
wire net2544;
wire net603;
wire net9202;
wire net4290;
wire net3063;
wire net1153;
wire net599;
wire net8439;
wire net328;
wire net766;
wire net6707;
wire net3454;
wire net7026;
wire net1573;
wire net2608;
wire net591;
wire net996;
wire net6373;
wire net2260;
wire net2973;
wire net4591;
wire net1113;
wire net2475;
wire net587;
wire net934;
wire net1863;
wire net3920;
wire net9401;
wire net1415;
wire net7698;
wire net6205;
wire net8419;
wire net3608;
wire net5881;
wire net7868;
wire net1560;
wire net650;
wire net7877;
wire net6824;
wire net58;
wire net8484;
wire net3217;
wire net9241;
wire net8843;
wire net5268;
wire net85;
wire net3027;
wire net4266;
wire net9615;
wire net4927;
wire net4347;
wire net7363;
wire net4143;
wire net186;
wire net8259;
wire net3073;
wire net1882;
wire net1393;
wire net9853;
wire net4348;
wire net710;
wire net3249;
wire net4529;
wire net1976;
wire net612;
wire net1010;
wire net957;
wire net5236;
wire net573;
wire net864;
wire net4998;
wire net3060;
wire net4745;
wire net3056;
wire net357;
wire net1965;
wire net768;
wire net1014;
wire net1681;
wire net8977;
wire net247;
wire net1687;
wire net5889;
wire net4282;
wire net564;
wire net3914;
wire net4577;
wire net6879;
wire net2020;
wire net1772;
wire net4498;
wire net189;
wire net5191;
wire net383;
wire net2788;
wire net1673;
wire net3782;
wire net555;
wire net1379;
wire net3737;
wire net553;
wire net2205;
wire net6826;
wire net9044;
wire net2636;
wire net7294;
wire net551;
wire net10407;
wire net8130;
wire net4390;
wire net1063;
wire net549;
wire net10258;
wire net3595;
wire net1428;
wire net6792;
wire net6363;
wire net546;
wire net2580;
wire net6680;
wire net5961;
wire net544;
wire net6353;
wire net3262;
wire net9410;
wire net4896;
wire net3661;
wire net1;
wire net7385;
wire net2602;
wire in3;
wire net1270;
wire net4584;
wire net2584;
wire net896;
wire net7402;
wire net2029;
wire net535;
wire net3168;
wire net1552;
wire net9453;
wire net2729;
wire net2726;
wire net642;
wire net2159;
wire net659;
wire net830;
wire net3610;
wire net4431;
wire net729;
wire net3379;
wire net823;
wire net1250;
wire net2117;
wire net1695;
wire net3860;
wire net1886;
wire net1468;
wire net7830;
wire net3445;
wire net98;
wire net524;
wire net4001;
wire net876;
wire net1052;
wire net3587;
wire net3333;
wire net5180;
wire net2079;
wire net9509;
wire net2953;
wire net297;
wire net10006;
wire net8729;
wire net5055;
wire net516;
wire net2779;
wire net1472;
wire net1793;
wire net6982;
wire net8290;
wire net7552;
wire net514;
wire net8942;
wire net511;
wire net4685;
wire net3618;
wire net1335;
wire net5148;
wire net4151;
wire net685;
wire net107;
wire net2539;
wire net3881;
wire net269;
wire net9652;
wire net346;
wire net8575;
wire net510;
wire net7122;
wire net1233;
wire net1025;
wire net506;
wire net927;
wire net3100;
wire net333;
wire net9466;
wire net3062;
wire net3214;
wire net1927;
wire net975;
wire net1952;
wire net505;
wire net2864;
wire net9804;
wire net8629;
wire net8256;
wire net3550;
wire net6150;
wire net1376;
wire net2630;
wire net1409;
wire net3696;
wire net1437;
wire net1829;
wire net1032;
wire net9595;
wire net8255;
wire net3086;
wire net501;
wire net2931;
wire net3407;
wire net1481;
wire net652;
wire net495;
wire net7364;
wire net494;
wire net988;
wire net492;
wire net2143;
wire net489;
wire net485;
wire net2745;
wire net985;
wire net488;
wire net646;
wire net838;
wire net5396;
wire net2170;
wire net475;
wire net6502;
wire net8275;
wire net2209;
wire net639;
wire net674;
wire net525;
wire net3400;
wire net7875;
wire net474;
wire net3094;
wire net4975;
wire net1867;
wire net8834;
wire net473;
wire net6157;
wire net2955;
wire net1145;
wire net4658;
wire net472;
wire net3331;
wire net3340;
wire net1347;
wire net3101;
wire net3958;
wire net3707;
wire net2616;
wire net3061;
wire net2331;
wire net967;
wire net5346;
wire net6035;
wire net3646;
wire net7051;
wire net1057;
wire net2675;
wire net1567;
wire net1272;
wire net2176;
wire net10410;
wire net4372;
wire net8014;
wire net780;
wire net7202;
wire net364;
wire net3395;
wire net1266;
wire net8121;
wire net7904;
wire net5097;
wire net6057;
wire net4099;
wire net5582;
wire net283;
wire net6856;
wire net9353;
wire net3289;
wire net10208;
wire net6002;
wire net2737;
wire net3127;
wire net1114;
wire net9066;
wire net3972;
wire net1295;
wire net10444;
wire net2056;
wire net3832;
wire net9408;
wire net3965;
wire net3159;
wire net459;
wire net545;
wire net6003;
wire net4225;
wire net453;
wire net624;
wire net629;
wire net731;
wire net450;
wire net7946;
wire net448;
wire net5559;
wire net1196;
wire net2122;
wire net5363;
wire net5;
wire net8898;
wire net1012;
wire net4443;
wire net3285;
wire net3944;
wire net9006;
wire net1074;
wire net2216;
wire net3704;
wire net561;
wire net444;
wire net8656;
wire net2638;
wire net2071;
wire net1374;
wire net3621;
wire net10389;
wire net8950;
wire net8904;
wire net504;
wire net2997;
wire net336;
wire net280;
wire net8881;
wire net969;
wire net437;
wire net4483;
wire net7764;
wire net3064;
wire net3631;
wire net8926;
wire net162;
wire net1017;
wire net4787;
wire net10315;
wire net718;
wire net6725;
wire net2430;
wire net4893;
wire net3095;
wire net5764;
wire net3900;
wire net10383;
wire net8612;
wire net432;
wire net1761;
wire net5294;
wire net8706;
wire net2118;
wire net1645;
wire net428;
wire net774;
wire net556;
wire net3312;
wire net2706;
wire net7487;
wire net771;
wire net5184;
wire net5648;
wire net928;
wire net1336;
wire net1220;
wire net5235;
wire net3033;
wire net293;
wire net2324;
wire net2107;
wire net5829;
wire net689;
wire net7218;
wire net422;
wire net1743;
wire clk;
wire net5308;
wire net2637;
wire net3122;
wire net6691;
wire net3576;
wire net4327;
wire net382;
wire net563;
wire net5841;
wire net1188;
wire net3663;
wire net5465;
wire net758;
wire net8650;
wire net2746;
wire net1625;
wire net417;
wire net901;
wire net10547;
wire net2030;
wire net3791;
wire net415;
wire net4389;
wire net5217;
wire net3142;
wire net4781;
wire net412;
wire net748;
wire net1224;
wire net2299;
wire net9118;
wire net702;
wire net5077;
wire net7425;
wire net634;
wire net1981;
wire net3838;
wire net7610;
wire net5879;
wire net554;
wire net4216;
wire net9725;
wire net1192;
wire net6786;
wire net7583;
wire net2597;
wire net3939;
wire net8071;
wire net3026;
wire net3721;
wire net4454;
wire net680;
wire net2677;
wire net6442;
wire net6797;
wire net403;
wire net4296;
wire net2066;
wire net2943;
wire net4852;
wire net8878;
wire net7053;
wire net1330;
wire net3216;
wire net3274;
wire net9128;
wire net5131;
wire net854;
wire net8922;
wire net2656;
wire net4833;
wire net5512;
wire net8320;
wire net1678;
wire net1236;
wire net3397;
wire net166;
wire net1621;
wire net6466;
wire net388;
wire net402;
wire net387;
wire net2924;
wire net1097;
wire net3565;
wire net4489;
wire net4243;
wire net1874;
wire net385;
wire in21;
wire net10304;
wire net9818;
wire net5303;
wire net2825;
wire net384;
wire net2050;
wire net2456;
wire net885;
wire net2234;
wire net3639;
wire net2156;
wire net8655;
wire net207;
wire net317;
wire net7528;
wire net3273;
wire net1089;
wire net4610;
wire net5482;
wire net6548;
wire net10078;
wire net1666;
wire net4400;
wire net1277;
wire net2298;
wire net155;
wire net1087;
wire net2070;
wire net3858;
wire net3344;
wire net3568;
wire net5048;
wire net2934;
wire net1034;
wire in8;
wire net4370;
wire net4449;
wire net10361;
wire net4818;
wire net6296;
wire net759;
wire net1518;
wire net2089;
wire net3399;
wire net5358;
wire net152;
wire net139;
wire net5987;
wire net895;
wire net1249;
wire net3651;
wire net742;
wire net8947;
wire net2759;
wire net2893;
wire net4689;
wire net9642;
wire net5682;
wire net2533;
wire net3680;
wire net2025;
wire net132;
wire net7713;
wire net1221;
wire net862;
wire net131;
wire net6498;
wire net733;
wire net2673;
wire net129;
wire net2529;
wire net4453;
wire net5780;
wire net10513;
wire net7044;
wire net3418;
wire net633;
wire net318;
wire net2304;
wire net9486;
wire net8772;
wire net7029;
wire net810;
wire net6735;
wire net6853;
wire net6986;
wire net258;
wire net10207;
wire net2789;
wire net3115;
wire net5563;
wire net123;
wire net592;
wire net7466;
wire net117;
wire net3973;
wire net9553;
wire net121;
wire net5976;
wire net1297;
wire net0;
wire net3167;
wire net4303;
wire net8985;
wire net1982;
wire net10130;
wire net3403;
wire net462;
wire net653;
wire net3682;
wire net5759;
wire net1617;
wire net4306;
wire net285;
wire net600;
wire net5877;
wire net1234;
wire net7821;
wire net2236;
wire net1043;
wire net8020;
wire net4579;
wire net2995;
wire net9936;
wire net73;
wire net4401;
wire net825;
wire net4402;
wire net10019;
wire net1765;
wire net113;
wire net2550;
wire net6089;
wire net752;
wire net3290;
wire net1332;
wire net309;
wire net791;
wire net4218;
wire net7370;
wire net538;
wire net833;
wire net8592;
wire in13;
wire net10065;
wire net4239;
wire net311;
wire net362;
wire net1226;
wire net978;
wire net2712;
wire net110;
wire net949;
wire net886;
wire net8618;
wire net2374;
wire net890;
wire net4075;
wire net2709;
wire net6153;
wire net69;
wire net8502;
wire net793;
wire net2167;
wire net9779;
wire net846;
wire net1569;
wire net4041;
wire net10374;
wire net627;
wire net59;
wire net717;
wire net3443;
wire net874;
wire net7622;
wire net695;
wire net7467;
wire net1658;
wire net5258;
wire net513;
wire net9946;
wire net6147;
wire net3372;
wire net3113;
wire net6652;
wire net463;
wire net751;
wire net1551;
wire net915;
wire net7145;
wire net103;
wire net5609;
wire net2848;
wire net44;
wire net849;
wire net100;
wire net97;
wire net2964;
wire net4411;
wire net6095;
wire net1878;
wire net394;
wire net4866;
wire net4993;
wire net3311;
wire net8537;
wire net787;
wire net2819;
wire net239;
wire net10002;
wire net27;
wire net195;
wire net1929;
wire net657;
wire net3945;
wire net94;
wire net1185;
wire net8487;
wire net2067;
wire net6663;
wire in12;
wire net9402;
wire net409;
wire net482;
wire net264;
wire net209;
wire net4683;
wire net582;
wire net3332;
wire net2646;
wire net8694;
wire net6530;
wire net5379;
wire net971;
wire net6921;
wire net88;
wire net1900;
wire net4553;
wire net9403;
wire net3164;
wire net5893;
wire net5243;
wire net735;
wire net99;
wire net3505;
wire net925;
wire net9984;
wire net7880;
wire net5406;
wire net2485;
wire net826;
wire net3179;
wire net199;
wire net2318;
wire net458;
wire net6760;
wire net678;
wire net262;
wire net1287;
wire net4759;
wire net3633;
wire net3571;
wire net1789;
wire net5407;
wire net87;
wire net7177;
wire net5568;
wire net290;
wire net66;
wire net8963;
wire net5473;
wire net6737;
wire net5112;
wire net1710;
wire net486;
wire net9969;
wire net9012;
wire net7278;
wire net2357;
wire net1046;
wire net10550;
wire net6360;
wire net857;
wire net81;
wire net3298;
wire net9420;
wire net3420;
wire net2264;
wire net2514;
wire net7216;
wire net6596;
wire net9962;
wire net202;
wire net5040;
wire net2339;
wire net572;
wire net3795;
wire net7728;
wire net1212;
wire net1545;
wire net2428;
wire net11;
wire net3322;
wire net1448;
wire in7;
wire net374;
wire net9296;
wire net4447;
wire net799;
wire net1486;
wire net1707;
wire net4162;
wire net7982;
wire net6356;
wire net2074;
wire net2100;
wire net889;
wire net8835;
wire net877;
wire net490;
wire net1064;
wire net2647;
wire net8640;
wire net298;
wire net467;
wire net241;
wire net851;
wire net9;
wire net1028;
wire net6017;
wire net998;
wire net9943;
wire net3166;
wire net4373;
wire net160;
wire net1223;
wire net765;
wire net2853;
wire net252;
wire net10101;
wire net8287;
wire net7470;
wire net1603;
wire net31;
wire net288;
wire net2200;
wire net441;
wire net673;
wire net1314;
wire net3402;
wire net2155;
wire net6957;
wire net3236;
wire net2283;
wire net3686;
wire net773;
wire net3391;
wire net4653;
wire net7092;
wire net3303;
wire in6;
wire net4619;
wire net167;
wire net1414;
wire net9712;
wire net2876;
wire net2750;
wire net2189;
wire net9255;
wire net7320;
wire net2330;
wire net891;
wire net5617;
wire net8221;
wire net3304;
wire net8422;
wire net6381;
wire net75;
wire net2053;
wire net2513;
wire net8308;
wire net523;
wire net9082;
wire net2983;
wire net45;
wire net5488;
wire net3171;
wire net4979;
wire net935;
wire net3468;
wire net5603;
wire net4;
wire net9110;
wire net334;
wire net2268;
wire net477;
wire net9844;
wire net1489;
wire net2522;
wire net481;
wire net3299;
wire net6;
wire net8531;
wire net5913;
wire net665;
wire net2371;
wire net9609;
wire net1788;
wire net9093;
wire net4362;
wire net5602;
wire net379;
wire net197;
wire net6612;
wire net1387;
wire net10380;
wire net779;
wire net10467;
wire net3414;
wire net106;
wire net8896;
wire net6509;
wire net5350;
wire net995;
wire net7575;
wire net3876;
wire net2451;
wire net566;
wire net1210;
wire net1172;
wire net1498;
wire net7788;
wire net2621;
wire net1419;
wire net2670;
wire net68;
wire net6400;
wire net1405;
wire net7406;
wire net723;
wire net1177;
wire net6344;
wire net1110;
wire net696;
wire net4074;
wire net2008;
wire net8511;
wire net1632;
wire net7069;
wire net8177;
wire net7825;
wire net245;
wire net3192;
wire net1834;
wire net2839;
wire net2396;
wire net6079;
wire net3592;
wire net667;
wire net3452;
wire net18;
wire net1214;
wire net7061;
wire net90;
wire net10165;
wire net5947;
wire net1425;
wire net8;
wire net8609;
wire net1677;
wire net1727;
wire net3460;
wire net2849;
wire net2688;
wire net2804;
wire net2082;
wire net1443;
wire in23;
wire net3558;
wire net5866;
wire net7907;
wire net7630;
wire net4017;
wire net9646;
wire net9608;
wire net163;
wire net3170;
wire net7414;
wire net51;
wire net5680;
wire net10371;
wire net2034;
wire net5800;
wire net2285;
wire net726;
wire net1165;
wire net5577;
wire net5748;
wire net7132;
wire net10496;
wire net7800;
wire net347;
wire net5090;
wire net1007;
wire net1408;
wire net6909;
wire net2526;
wire net9637;
wire net4910;
wire net84;
wire net2577;
wire net2667;
wire net6122;
wire net398;
wire net1610;
wire net2363;
wire net7966;
wire net6188;
wire net3128;
wire in4;
wire net3309;
wire net1971;
wire net9526;
wire net240;
wire net9379;
wire net4799;
wire net1885;
wire net175;
wire net682;
wire net570;
wire net1777;
wire net7805;
wire net274;
wire in16;
wire net1549;
wire net4497;
wire net5886;
wire net2308;
wire net1252;
wire net1503;
wire net1676;
wire net5216;
wire net2633;
wire net496;
wire net1055;
wire net426;
wire net8441;
wire net348;
wire net1668;
wire net962;
wire net10420;
wire net36;
wire net4441;
wire net507;
wire net5673;
wire net1338;
wire net2201;
wire net671;
wire net7381;
wire net7491;
wire net3383;
wire net8595;
wire net21;
wire net143;
wire net609;
wire net1421;
wire net920;
wire net6911;
wire net3450;
wire net625;
wire net393;
wire net522;
wire net2463;
wire net1745;
wire in20;
wire net491;
wire net818;
wire net4988;
wire net300;
wire net157;
wire net2081;
wire net10336;
wire net1935;
wire net95;
wire net7596;
wire net79;
wire net835;
wire net20;
wire net4002;
wire net10079;
wire net86;
wire net601;
wire net2256;
wire net3361;
wire net1530;
wire net3983;
wire net154;
wire net1006;
wire net9930;
wire net4260;
wire net6706;
wire net7658;
wire net1893;
wire net251;
wire net1420;
wire net5449;
wire in18;
wire net6484;
wire net775;
wire net10527;
wire net3364;
wire net254;
wire net7646;
wire net64;
wire net8013;
wire net408;
wire net4063;
wire net2530;
wire net2049;
wire net951;
wire net12;
wire net536;
wire net7897;
wire net83;
wire net33;
wire net4167;
wire net1011;
wire net9873;
wire net2150;
wire net185;
wire net5637;
wire net10347;
wire net4738;
wire net5792;
wire net3200;
wire net1820;
wire net5699;
wire net638;
wire net8755;
wire net128;
wire net5392;
wire net3176;
wire net2866;
wire net7818;
wire net2980;
wire net4326;
wire net1205;
wire net37;
wire net2384;
wire net7124;
wire net4184;
wire net530;
wire net9391;
wire net5117;
wire net6156;
wire net1511;
wire net38;
wire net3569;
wire net3630;
wire net127;
wire net7257;
wire net1346;
wire net2814;
wire net569;
wire net502;
wire net158;
wire net6458;
wire net6724;
wire net3428;
wire net145;
wire net8194;
wire net213;
wire net5936;
wire net7834;
wire net499;
wire net6278;
wire net50;
wire net2128;
wire net6069;
wire net2103;
wire net4945;
wire net7355;
wire net229;
wire net732;
wire net4869;
wire net457;
wire net645;
wire net4668;
wire net1636;
wire net479;
wire net149;
wire net10316;
wire net57;
wire net6006;
wire net984;
wire net8126;
wire net3495;
wire net2838;
wire net3845;
wire net3172;
wire net9284;
wire net137;
wire net2203;
wire net3182;
wire net4960;
wire net7494;
wire net5024;
wire net5436;
wire net5481;
wire net9480;
wire net6303;
wire net1586;
wire net3843;
wire net1148;
wire net1168;
wire net10460;
wire net2346;
wire net380;
wire net3197;
wire net359;
wire net993;
wire net191;
wire net755;
wire net47;
wire net5013;
wire net3625;
wire net1104;
wire net5834;
wire net512;
wire net7282;
wire net3052;
wire net2415;
wire net8743;
wire net7074;
wire net1305;
wire net13;
wire net3899;
wire net3001;
wire net3421;
wire net89;
wire net2942;
wire net741;
wire net3534;
wire net10063;
wire net3446;
wire net6818;
wire net944;
wire net1714;
wire net5177;
wire net5267;
wire net9489;
wire net3465;
wire net6885;
wire net1213;
wire net1410;
wire net3188;
wire net395;
wire net6733;
wire net2992;
wire net2387;
wire net49;
wire net6702;
wire net7021;
wire net664;
wire net9866;
wire net7618;
wire net296;
wire net10171;
wire net855;
wire net55;
wire net134;
wire net3474;
wire net3585;
wire net1182;
wire net4054;
wire net5928;
wire net6941;
wire net6717;
wire net2212;
wire in1;
wire net74;
wire net4692;
wire net2617;
wire out9;
wire net2077;
wire net210;
wire net3254;
wire net4098;
wire net1954;
wire net4211;
wire net1237;
wire net10220;
wire net1317;
wire net9119;
wire net7331;
wire net5977;
wire net176;
wire net80;
wire net756;
wire net1970;
wire net1858;
wire net9277;
wire net1243;
wire net1284;
wire net2857;
wire net5306;
wire net1639;
wire net852;
wire net3683;
wire net1465;
wire net6064;
wire net3642;
wire net445;
wire net7490;
wire net3785;
wire net5053;
wire net5661;
wire net9686;
wire net8617;
wire net70;
wire net2193;
wire net279;
wire net3453;
wire net2;
wire net2468;
wire net192;
wire net594;
wire net174;
wire net6092;
wire net560;
wire net1755;
wire net225;
wire net1653;
wire net7705;
wire net265;
wire net6474;
wire net9186;
wire net1804;
wire net2437;
wire net96;
wire net8230;
wire net3513;
wire net4939;
wire in2;
wire net610;
wire net180;
wire net4252;
wire net550;
wire net4520;
wire net3694;
wire net1542;
wire net3434;
wire net4153;
wire net5132;
wire net1447;
wire net9582;
wire net101;
wire net3784;
wire net3711;
wire net281;
wire net181;
wire net698;
wire net3510;
wire net1986;
wire net2278;
wire net182;
wire net3201;
wire net641;
wire net7604;
wire net6990;
wire net1033;
wire net7613;
wire net785;
wire net701;
wire net286;
wire net5221;
wire net8742;
wire net2547;
wire net3139;
wire net476;
wire net3393;
wire net722;
wire net1095;
wire net4832;
wire net1803;
wire net301;
wire net1683;
wire net3315;
wire net8573;
wire net2427;
wire net345;
wire net3461;
wire net537;
wire net1881;
wire net10342;
wire net5373;
wire net8759;
wire net7429;
wire net2703;
wire net4460;
wire net966;
wire net4924;
wire net2333;
wire net1016;
wire net8099;
wire net193;
wire net1348;
wire net7042;
wire net48;
wire net8774;
wire net2627;
wire net194;
wire net3927;
wire net4337;
wire net5628;
wire net198;
wire net360;
wire net2833;
wire net2012;
wire net8841;
wire net6549;
wire net6881;
wire net236;
wire net9445;
wire net320;
wire net4304;
wire net295;
wire net204;
wire net3620;
wire net8824;
wire net3174;
wire net3613;
wire net7942;
wire net7692;
wire net3747;
wire net589;
wire net53;
wire net583;
wire net214;
wire net3665;
wire net9882;
wire net6994;
wire net7441;
wire net1262;
wire net8010;
wire net767;
wire net3797;
wire net7147;
wire net237;
wire net4255;
wire net9848;
wire net480;
wire net5681;
wire net8282;
wire net1901;
wire net924;
wire net9127;
wire net2701;
wire net3898;
wire net3320;
wire net233;
wire net6744;
wire net8482;
wire net3718;
wire net220;
wire net6131;
wire net520;
wire net981;
wire net3892;
wire net7440;
wire net366;
wire net607;
wire net7080;
wire net651;
wire net7768;
wire net620;
wire net6997;
wire net939;
wire net3347;
wire net10454;
wire net4586;
wire net3773;
wire net5152;
wire net1614;
wire net2486;
wire net452;
wire net2372;
wire net2592;
wire net63;
wire net2227;
wire net7139;
wire net10264;
wire net1371;
wire net613;
wire net6914;
wire net760;
wire net7303;
wire net223;
wire net5362;
wire net4996;
wire net897;
wire net908;
wire net438;
wire net10362;
wire net9134;
wire net2994;
wire net2678;
wire net10074;
wire net6517;
wire net8690;
wire net227;
wire net3611;
wire net9021;
wire net7346;
wire in9;
wire net660;
wire net6036;
wire net6414;
wire net542;
wire net2702;
wire net1326;
wire net628;
wire net2914;
wire net9184;
wire net5518;
wire net1748;
wire net526;
wire net1495;
wire net2573;
wire net4605;
wire net10309;
wire net230;
wire net1492;
wire net3755;
wire net3297;
wire net5186;
wire net577;
wire net5095;
wire net661;
wire net1910;
wire net1467;
wire net10049;
wire net7469;
wire net4773;
wire net3147;
wire net8167;
wire net2202;
wire net8398;
wire net5061;
wire net4774;
wire net418;
wire net323;
wire net10245;
wire net552;
wire net2899;
wire net244;
wire net3701;
wire net7782;
wire net7219;
wire net2773;
wire net905;
wire net338;
wire net672;
wire net3098;
wire net4273;
wire net2865;
wire net1790;
wire net24;
wire net1602;
wire net3640;
wire net801;
wire net2147;
wire net5087;
wire net249;
wire net8436;
wire net7550;
wire net5218;
wire net8132;
wire net1593;
wire net9246;
wire net3417;
wire net5943;
wire net9619;
wire net6070;
wire net5696;
wire net2132;
wire net10134;
wire net9257;
wire net3915;
wire net5610;
wire net8859;
wire net3463;
wire net518;
wire net3848;
wire net10356;
wire net1499;
wire net2911;
wire net7792;
wire net3605;
wire net5952;
wire net6198;
wire net183;
wire net1434;
wire net272;
wire net1558;
wire net902;
wire net200;
wire net635;
wire net8829;
wire net8243;
wire net5195;
wire net6256;
wire net3771;
wire net234;
wire net4545;
wire net598;
wire net1538;
wire net4130;
wire net4798;
wire net961;
wire net884;
wire net6277;
wire net487;
wire net6743;
wire net261;
wire net7515;
wire net1253;
wire net315;
wire net9775;
wire net1137;
wire net3441;
wire net1426;
wire net5586;
wire net7680;
wire net493;
wire net263;
wire net2221;
wire net4384;
wire net10059;
wire net8594;
wire net8359;
wire net112;
wire net3923;
wire net6094;
wire net1396;
wire net8906;
wire net2916;
wire net2477;
wire net4120;
wire net2654;
wire net2199;
wire net6423;
wire net5460;
wire net6647;
wire net8386;
wire net663;
wire net1821;
wire net6421;
wire net372;
wire net8277;
wire net2419;
wire net10156;
wire net7396;
wire net443;
wire net17;
wire net270;
wire net8616;
wire net7820;
wire net3689;
wire net757;
wire net9635;
wire net1384;
wire net6951;
wire net997;
wire net7962;
wire net5309;
wire net3;
wire net2293;
wire net4636;
wire net727;
wire net344;
wire net9259;
wire net6063;
wire net9380;
wire net3770;
wire net5906;
wire net9903;
wire net3475;
wire net4763;
wire net1643;
wire net2778;
wire net5341;
wire net878;
wire net593;
wire net278;
wire net7700;
wire net3685;
wire net1163;
wire in10;
wire net4961;
wire net436;
wire net2140;
wire net3374;
wire net4930;
wire net1001;
wire net4179;
wire net7084;
wire net2861;
wire net161;
wire net7544;
wire net5639;
wire net291;
wire net9098;
wire net5966;
wire net9880;
wire net1595;
wire net1836;
wire net588;
wire net529;
wire net376;
wire net1359;
wire net10122;
wire net4317;
wire net370;
wire net3617;
wire net19;
wire net4884;
wire net5159;
wire net306;
wire net4944;
wire net1717;
wire net1778;
wire net8914;
wire net1026;
wire net10327;
wire net1009;
wire net446;
wire net141;
wire net9940;
wire net8909;
wire net7162;
wire net3009;
wire net1684;
wire net784;
wire net1696;
wire net7775;
wire net3245;
wire net10514;
wire net5108;
wire net1862;
wire net130;
wire net1204;
wire net4821;
wire net9658;
wire net932;
wire net7156;
wire net217;
wire net312;
wire net1018;
wire net332;
wire net1158;
wire net93;
wire net9949;
wire net5315;
wire net7;
wire net10;
wire net2327;
wire net9235;
wire net8734;
wire in22;
wire net2935;
wire net7127;
wire net3007;
wire net2365;
wire net4868;
wire net9317;
wire net3531;
wire net455;
wire net2855;
wire net423;
wire net958;
wire net3185;
wire net976;
wire net4633;
wire net8503;
wire net2289;
wire net72;
wire net3132;
wire net7858;
wire net221;
wire net965;
wire net337;
wire net4568;
wire net968;
wire net7246;
wire net4507;
wire net7408;
wire net9318;
wire net3577;
wire net1452;
wire net5965;
wire net3676;
wire net2554;
wire net3667;
wire net3270;
wire net3573;
wire net1440;
wire net367;
wire net2821;
wire net597;
wire net3229;
wire net704;
wire net349;
wire net8399;
wire net2556;
wire net1200;
wire net2002;
wire net5497;
wire net9676;
wire net2552;
wire net2805;
wire net4455;
wire net464;
wire net6712;
wire net1635;
wire net356;
wire net9177;
wire net2815;
wire net8463;
wire net2093;
wire net1823;
wire net9478;
wire net1693;
wire net8054;
wire net2764;
wire net4213;
wire net371;
wire net1756;
wire net859;
wire net4750;
wire net6490;
wire net4451;
wire net3969;
wire net373;
wire net7936;
wire net4202;
wire net800;
wire net9149;
wire net3628;
wire net2629;
wire net3913;
wire net807;
wire net811;
wire net8505;
wire net812;
wire net9722;
wire net5953;
wire net1059;
wire net813;
wire net5326;
wire net1588;
wire net275;
wire net6019;
wire net7361;
wire net5292;
wire net196;
wire net1925;
wire net3119;
wire net10121;
wire net4840;
wire net6580;
wire net816;
wire net6703;
wire net8591;
wire net2473;
wire net1310;
wire net819;
wire net3745;
wire net822;
wire net1528;
wire net3238;
wire net824;
wire net3769;
wire net2639;
wire net1462;
wire net6441;
wire net2736;
wire net3435;
wire net6307;
wire net4696;
wire net831;
wire net3760;
wire net832;
wire net3856;
wire net7368;
wire net9926;
wire net7072;
wire net3702;
wire net2069;
wire in25;
wire net4542;
wire net102;
wire net5349;
wire net841;
wire net1369;
wire net843;
wire net844;
wire net5536;
wire net2231;
wire net71;
wire net2235;
wire net845;
wire net4330;
wire net7245;
wire net839;
wire net3356;
wire net894;
wire net1068;
wire net6237;
wire net1892;
wire net5882;
wire net1832;
wire net368;
wire net1159;
wire net7031;
wire net1839;
wire net856;
wire net10097;
wire net3244;
wire net809;
wire net858;
wire net2728;
wire net1449;
wire net1021;
wire net4190;
wire net1736;
wire net860;
wire net972;
wire net2813;
wire net863;
wire net5712;
wire net4737;
wire net3908;
wire net7967;
wire net2507;
wire net1482;
wire net3471;
wire net2062;
wire net866;
wire net868;
wire net10056;
wire net5279;
wire net2031;
wire net4500;
wire net1507;
wire net5525;
wire net869;
wire net5084;
wire net5399;
wire net6088;
wire net1450;
wire net6799;
wire net871;
wire net1968;
wire net1367;
wire net873;
wire net2698;
wire net5874;
wire net989;
wire net7260;
wire net2458;
wire net6832;
wire net3561;
wire net10119;
wire net4972;
wire net879;
wire net8770;
wire net3852;
wire net9327;
wire net5010;
wire net6861;
wire net3398;
wire net1401;
wire net1083;
wire net259;
wire net1065;
wire net881;
wire net5335;
wire net2927;
wire net1930;
wire net1973;
wire net6948;
wire net887;
wire net656;
wire net5993;
wire net892;
wire net7872;
wire net4487;
wire net893;
wire net10344;
wire net7326;
wire net6149;
wire net898;
wire net6404;
wire net3266;
wire net6956;
wire net903;
wire net4521;
wire net2889;
wire net5283;
wire net1259;
wire net7798;
wire net3753;
wire net906;
wire net9824;
wire net378;
wire net4111;
wire net955;
wire net6170;
wire net910;
wire net8557;
wire net3432;
wire net1329;
wire net5019;
wire net911;
wire net2697;
wire net4309;
wire net608;
wire net913;
wire net4855;
wire net2447;
wire net714;
wire net922;
wire net3873;
wire net2457;
wire net4973;
wire net2311;
wire net1207;
wire net10050;
wire net926;
wire net5864;
wire net7249;
wire net9365;
wire net616;
wire net1608;
wire net6566;
wire net584;
wire net7314;
wire net930;
wire net2131;
wire net5946;
wire net3089;
wire net5833;
wire net2323;
wire net933;
wire net2593;
wire net4933;
wire net2294;
wire net4104;
wire net4124;
wire net5741;
wire net1509;
wire net4535;
wire net1298;
wire net936;
wire net788;
wire net3654;
wire net8416;
wire net1955;
wire net6145;
wire net8910;
wire net1339;
wire net4338;
wire net938;
wire net940;
wire net3761;
wire net3813;
wire net7178;
wire net3405;
wire net3979;
wire net8790;
wire net1147;
wire net5633;
wire net9952;
wire net1093;
wire net941;
wire net1737;
wire net943;
wire net4220;
wire net1657;
wire net990;
wire net7677;
wire net946;
wire net1980;
wire net3189;
wire net1907;
wire net6461;
wire net7896;
wire net1364;
wire net1191;
wire net1136;
wire net6214;
wire net8267;
wire net3093;
wire net948;
wire net614;
wire net5026;
wire net2414;
wire net6419;
wire net1969;
wire net8313;
wire net5403;
wire net1024;
wire net3226;
wire net4409;
wire net8041;
wire net953;
wire net3329;
wire net5784;
wire net954;
wire net2223;
wire net1183;
wire net959;
wire net248;
wire net6128;
wire net7901;
wire net4076;
wire net2609;
wire net5354;
wire net5814;
wire net170;
wire net1194;
wire net391;
wire net1407;
wire net331;
wire net78;
wire net963;
wire net521;
wire net4931;
wire net5700;
wire net9913;
wire net1027;
wire net8818;
wire net1816;
wire net1661;
wire net974;
wire net6288;
wire net5583;
wire net2004;
wire net979;
wire net980;
wire out16;
wire net1700;
wire net6723;
wire net4557;
wire net983;
wire net3282;
wire net8506;
wire net815;
wire net991;
wire net203;
wire net2267;
wire net1299;
wire net1928;
wire net6476;
wire net2856;
wire net1776;
wire net1000;
wire net3150;
wire net1003;
wire net466;
wire net2854;
wire net4139;
wire net789;
wire net1005;
wire net1008;
wire net3591;
wire net6654;
wire net2897;
wire net1427;
wire net8229;
wire net3604;
wire net8088;
wire net2662;
wire net1013;
wire net882;
wire net3343;
wire net3208;
wire net10370;
wire net1629;
wire net416;
wire net4440;
wire net1023;
wire net2537;
wire net498;
wire net4856;
wire net1541;
wire net528;
wire net6203;
wire net1115;
wire net6766;
wire net10205;
wire net2198;
wire net5411;
wire net1031;
wire net1694;
wire net2799;
wire net4429;
wire net1035;
wire net7883;
wire net4482;
wire net5263;
wire net284;
wire net5660;
wire net1510;
wire net29;
wire net4527;
wire net606;
wire net4646;
wire net7957;
wire net1036;
wire net3263;
wire net4394;
wire net1871;
wire net9302;
wire net694;
wire net2770;
wire net1042;
wire net4513;
wire net9744;
wire net7345;
wire net9510;
wire net3703;
wire net567;
wire net1044;
wire net630;
wire net3048;
wire net7793;
wire net5668;
wire net1152;
wire net2895;
wire net5524;
wire net4010;
wire net2316;
wire net1045;
wire net2297;
wire net7637;
wire net1711;
wire net1400;
wire net5167;
wire net4267;
wire net1269;
wire net250;
wire net4990;
wire net2531;
wire net2613;
wire net5519;
wire net1048;
wire net6465;
wire net2755;
wire net1422;
wire net1879;
wire net10432;
wire net8420;
wire net1020;
wire net2492;
wire net1056;
wire net10314;
wire net2501;
wire net4425;
wire net5262;
wire net6697;
wire net6813;
wire net4601;
wire net5538;
wire net2454;
wire net5305;
wire net10434;
wire net602;
wire net1744;
wire net1062;
wire net9229;
wire net3751;
wire net10250;
wire net2614;
wire net1066;
wire net1067;
wire net6671;
wire net1071;
wire net42;
wire net5064;
wire net1072;
wire net4971;
wire net8967;
wire net8211;
wire net2780;
wire net1642;
wire net3231;
wire net9819;
wire net1622;
wire net2055;
wire net1630;
wire net7563;
wire net1073;
wire net1227;
wire net1076;
wire net1361;
wire net1150;
wire net9551;
wire net5038;
wire net2301;
wire net6455;
wire net9730;
wire net6267;
wire net1868;
wire net1079;
wire net5272;
wire net2472;
wire net92;
wire net2809;
wire net3886;
wire net1500;
wire net3962;
wire net9643;
wire net6434;
wire net880;
wire net6764;
wire net5410;
wire net739;
wire net1081;
wire net386;
wire net5669;
wire net2757;
wire net1094;
wire net1323;
wire net7223;
wire net142;
wire net2011;
wire net5447;
wire net2612;
wire net389;
wire net7481;
wire net1098;
wire net9150;
wire net1406;
wire net273;
wire net1099;
wire net1493;
wire net1101;
wire net1103;
wire net10568;
wire net9814;
wire net7102;
wire net1105;
wire net3152;
wire net5284;
wire net2405;
wire net6684;
wire net8133;
wire net16;
wire net2206;
wire net2455;
wire net4515;
wire net1108;
wire net3835;
wire net9584;
wire net5229;
wire net1978;
wire net3768;
wire net3069;
wire net1634;
wire net1665;
wire net1039;
wire net9440;
wire net4026;
wire net3072;
wire net5963;
wire net1112;
wire net1119;
wire net314;
wire net1090;
wire net1120;
wire net1523;
wire net4023;
wire net1126;
wire net7192;
wire net3365;
wire net1818;
wire net1127;
wire net1712;
wire net8440;
wire net1129;
wire net4336;
wire net5415;
wire net5455;
wire net1130;
wire net1131;
wire net4742;
wire net5210;
wire net3065;
wire net684;
wire net1132;
wire out23;
wire net1589;
wire net7589;
wire net1133;
wire net8340;
wire net3292;
wire net7095;
wire net3054;
wire net2644;
wire net6872;
wire net6225;
wire net2564;
wire net5165;
wire net6980;
wire net619;
wire net1141;
wire net2133;
wire net2594;
wire net4915;
wire net2488;
wire net5394;
wire out15;
wire net1144;
wire net4439;
wire net8767;
wire net1149;
wire net1077;
wire net456;
wire net7137;
wire net392;
wire net6234;
wire net10560;
wire net1230;
wire net9121;
wire net1652;
wire net1411;
wire net3602;
wire net2121;
wire net8599;
wire net1160;
wire net4060;
wire net2795;
wire net2976;
wire net2937;
wire net9707;
wire net2320;
wire net1161;
wire net6677;
wire net2715;
wire net2512;
wire net1164;
wire net1303;
wire net7239;
wire net2112;
wire net3499;
wire net1996;
wire net9101;
wire net6324;
wire net62;
wire net1171;
wire net2434;
wire net2540;
wire net5069;
wire net9521;
wire net3075;
wire net1174;
wire net6228;
wire net5421;
wire net201;
wire net9556;
wire net9092;
wire net1906;
wire net3566;
wire net2944;
wire net1180;
wire net5464;
wire net7319;
wire net2920;
wire net2139;
wire net2359;
wire net4908;
wire net3430;
wire net615;
wire net5820;
wire net460;
wire net6877;
wire net1184;
wire net2867;
wire net2239;
wire net8590;
wire net1799;
wire net1186;
wire net9626;
wire net821;
wire net9792;
wire net2449;
wire net9388;
wire net34;
wire net5867;
wire net9442;
wire net358;
wire net1516;
wire net4110;
wire net6761;
wire net8817;
wire net1281;
wire net3603;
wire net9662;
wire net8310;
wire net76;
wire net3887;
wire net1199;
wire net1268;
wire net1311;
wire net1201;
wire net1202;
wire net10166;
wire net4551;
wire net7702;
wire net4609;
wire net9776;
wire net3424;
wire net8662;
wire net6876;
wire net1206;
wire net3044;
wire net2090;
wire net558;
wire net4671;
wire net668;
wire net3422;
wire net1578;
wire net5838;
wire net1209;
wire net7328;
wire net9218;
wire net226;
wire net7638;
wire net1604;
wire net3138;
wire net1313;
wire net8698;
wire net1217;
wire net2403;
wire net4154;
wire net4313;
wire net120;
wire net2605;
wire net4493;
wire net1267;
wire net5645;
wire net2394;
wire net2099;
wire net1222;
wire net1491;
wire net1225;
wire net6591;
wire net1228;
wire net2369;
wire net2489;
wire net9921;
wire net2046;
wire net883;
wire net5483;
wire net964;
wire net5827;
wire net1232;
wire net256;
wire net1238;
wire net6636;
wire net2803;
wire net3091;
wire net2376;
wire net8563;
wire net8056;
wire net1240;
wire net8228;
wire net888;
wire net747;
wire net3520;
wire net1244;
wire net9414;
wire net5271;
wire net1718;
wire net5166;
wire net5974;
wire net215;
wire net1245;
wire net3627;
wire net6431;
wire net7465;
wire net3114;
wire net1248;
wire net2228;
wire net1251;
wire net4849;
wire net2794;
wire net3258;
wire net3104;
wire net1231;
wire net2868;
wire net140;
wire net1255;
wire net8674;
wire net2146;
wire net1162;
wire net3429;
wire net9049;
wire net1257;
wire net2991;
wire net4793;
wire net91;
wire net1990;
wire net67;
wire net401;
wire net5257;
wire net3970;
wire net654;
wire net1276;
wire net1278;
wire net8943;
wire net909;
wire net3960;
wire out21;
wire net4231;
wire net9125;
wire net5037;
wire net6927;
wire net1279;
wire net1598;
wire net6526;
wire net5758;
wire net798;
wire net1280;
wire net5724;
wire net8298;
wire net1307;
wire net7681;
wire net5378;
wire net2885;
wire net468;
wire net6398;
wire net421;
wire net1480;
wire net636;
wire net10227;
wire net3092;
wire net1282;
wire net4068;
wire net6221;
wire net6692;
wire net1283;
wire net5194;
wire net5400;
wire net9077;
wire net1357;
wire net1286;
wire net1288;
wire net7597;
wire net5774;
wire net1289;
wire net3551;
wire net1292;
wire net6576;
wire net2699;
wire net1296;
wire net1550;
wire net1911;
wire net10539;
wire net9062;
wire net4215;
wire net1301;
wire net1302;
wire net7353;
wire net688;
wire net1553;
wire net1471;
wire net4748;
wire net7158;
wire net1306;
wire net1585;
wire net8679;
wire net8184;
wire net4958;
wire net5277;
wire net10516;
wire net1316;
wire net2360;
wire net6774;
wire net440;
wire net7492;
wire net4133;
wire net1831;
wire net1522;
wire net1322;
wire net4230;
wire net2802;
wire net2558;
wire net5630;
wire net1327;
wire net5156;
wire net1398;
wire net3107;
wire net3790;
wire net1619;
wire net9117;
wire net1341;
wire net2406;
wire net1342;
wire net1350;
wire net1300;
wire net2464;
wire net5629;
wire net6148;
wire net1260;
wire net1351;
wire net4470;
wire net1355;
wire net5887;
wire net1483;
wire net8931;
wire net2958;
wire net4234;
wire net834;
wire net10262;
wire net5790;
wire net1360;
wire net3935;
wire net7463;
wire net2441;
wire net1627;
wire net1562;
wire net10040;
wire net3183;
wire net643;
wire net1319;
wire net7959;
wire net2169;
wire net1366;
wire net5057;
wire net2589;
wire net4462;
wire net952;
wire net3448;
wire net1580;
wire net6796;
wire net351;
wire net4452;
wire net8090;
wire net848;
wire net7226;
wire net1375;
wire net9872;
wire net3464;
wire net3925;
wire net973;
wire net451;
wire net2734;
wire net7685;
wire net1378;
wire net1092;
wire net6882;
wire net8703;
wire net1380;
wire net7828;
wire net1381;
wire net4387;
wire net10426;
wire net6425;
wire net9614;
wire net1382;
wire net10025;
wire net1389;
wire net2880;
wire net1435;
wire net9829;
wire net2466;
wire net804;
wire net3607;
wire net937;
wire net1385;
wire net1386;
wire net5539;
wire net1388;
wire net3045;
wire in15;
wire net711;
wire net1591;
wire net1784;
wire net7070;
wire net1391;
wire net2080;
wire net10203;
wire net2548;
wire net719;
wire net3572;
wire net1394;
wire net1395;
wire net2721;
wire net6905;
wire net1962;
wire net1399;
wire net8928;
wire net931;
wire net381;
wire net429;
wire net1402;
wire net7015;
wire net1403;
wire net2213;
wire net2982;
wire net484;
wire net2075;
wire net4768;
wire net1085;
wire net1404;
wire net828;
wire net2450;
wire net1413;
wire net321;
wire net4081;
wire net2883;
wire net7450;
wire net2775;
wire net6337;
wire net8775;
wire net405;
wire net10391;
wire net10069;
wire net7504;
wire net1424;
wire net2423;
wire net1431;
wire net6565;
wire net6264;
wire net1944;
wire net1637;
wire net1432;
wire net2929;
wire net1600;
wire net3386;
wire net1433;
wire net1607;
wire net2250;
wire net1157;
wire net8801;
wire net1438;
wire net1441;
wire net5553;
wire net9168;
wire net1344;
wire net1453;
wire net7101;
wire net7276;
wire net6472;
wire net697;
wire net4565;
wire net2999;
wire net433;
wire net6864;
wire net1333;
wire net1457;
wire net899;
wire net3537;
wire net1091;
wire net5837;
wire net1454;
wire net7506;
wire net5360;
wire net1455;
wire net2254;
wire net2641;
wire net1844;
wire net2065;
wire net7475;
wire net3050;
wire net1456;
wire net1458;
wire net2844;
wire net7295;
wire net576;
wire net3043;
wire net10195;
wire net1626;
wire net6971;
wire net2683;
wire net1143;
wire net6038;
wire net6682;
wire net1461;
wire net1579;
wire net3563;
wire net1353;
wire net6229;
wire net1469;
wire net1169;
wire net1084;
wire net7262;
wire net4622;
wire net5027;
wire net5778;
wire net6068;
wire net1470;
wire net3518;
wire net6637;
wire net929;
wire net1473;
wire net447;
wire net1189;
wire net1478;
wire net5009;
wire net7022;
wire net2175;
wire net1271;
wire net5779;
wire net10390;
wire net3154;
wire net1484;
wire net6186;
wire net6975;
wire net7650;
wire net803;
wire net4015;
wire net3144;
wire net3644;
wire net3255;
wire net3019;
wire net1494;
wire net4079;
wire net5062;
wire net1496;
wire net5688;
wire net2966;
wire net9037;
wire net1497;
wire net6114;
wire net7204;
wire net3013;
wire net3181;
wire net1950;
wire net1504;
wire net10191;
wire net8596;
wire net3524;
wire net1670;
wire net4393;
wire net829;
wire net10192;
wire net1506;
wire net6573;
wire net8278;
wire net8268;
wire net14;
wire net8384;
wire net5695;
wire net1512;
wire net5289;
wire net669;
wire net1513;
wire net10463;
wire net1514;
wire net10003;
wire net3549;
wire net1648;
wire net316;
wire net8481;
wire net1618;
wire net2562;
wire net7338;
wire net1916;
wire net1760;
wire net7418;
wire net8716;
wire net8200;
wire net1524;
wire net1833;
wire net709;
wire in14;
wire net9981;
wire net3984;
wire net6730;
wire net8866;
wire net2671;
wire net375;
wire net5647;
wire net1485;
wire net1531;
wire net6607;
wire net1533;
wire net10014;
wire net1536;
wire net3490;
wire net10103;
wire net1584;
wire net5549;
wire net1735;
wire net5614;
wire net122;
wire net1547;
wire net9264;
wire net2178;
wire net1798;
wire net5058;
wire net1548;
wire net3954;
wire net7011;
wire net6924;
wire net115;
wire net7457;
wire net1554;
wire net8108;
wire net6645;
wire net778;
wire net557;
wire net190;
wire net5599;
wire net1557;
wire net3479;
wire net1559;
wire net677;
wire net1570;
wire net1746;
wire net837;
wire net3793;
wire net4847;
wire net5776;
wire net7016;
wire net77;
wire net1843;
wire net956;
wire net796;
wire net6973;
wire net7159;
wire net4035;
wire net4374;
wire net1564;
wire net4072;
wire net2882;
wire net7635;
wire net2549;
wire net8748;
wire net1565;
wire net2116;
wire net3988;
wire net125;
wire net1926;
wire net1574;
wire net1576;
wire net2919;
wire net8064;
wire net4413;
wire net1577;
wire net3283;
wire net1581;
wire net5264;
wire net4039;
wire net1587;
wire net8352;
wire net2087;
wire net1963;
wire net1920;
wire net6989;
wire net1594;
wire net3457;
wire net8204;
wire net7235;
wire net7241;
wire net1285;
wire net1078;
wire net242;
wire net2141;
wire net7082;
wire net9770;
wire net1606;
wire net1924;
wire net7046;
wire net1609;
wire net2523;
wire net308;
wire net2266;
wire net4901;
wire net1167;
wire net2669;
wire net7103;
wire net3805;
wire net2785;
wire net942;
wire net5727;
wire net1572;
wire net7555;
wire net1304;
wire net1620;
wire net257;
wire net1852;
wire net5555;
wire net3415;
wire net9986;
wire net1623;
wire net2355;
wire net1124;
wire net7185;
wire net1697;
wire net3108;
wire net1633;
wire net4148;
wire net8192;
wire net3106;
wire net5579;
wire net5371;
wire net8582;
wire net618;
wire net2690;
wire net1641;
wire net527;
wire net1644;
wire net1646;
wire net1651;
wire net1650;
wire net4710;
wire net2909;
wire net2028;
wire net5440;
wire net4181;
wire net3117;
wire net4620;
wire net1490;
wire net4589;
wire net205;
wire net4058;
wire net4185;
wire net2774;
wire net1479;
wire net6351;
wire net867;
wire net1904;
wire net7945;
wire net1669;
wire net623;
wire net4200;
wire net10534;
wire net1671;
wire net8289;
wire net2686;
wire net2217;
wire net1672;
wire net3358;
wire net921;
wire net6483;
wire net712;
wire net1674;
wire net2824;
wire net3040;
wire net1682;
wire net108;
wire net3196;
wire net7296;
wire net7963;
wire net3241;
wire net9301;
wire net271;
wire net5242;
wire net5746;
wire net1685;
wire net3041;
wire net3933;
wire net1751;
wire net1703;
wire net1686;
wire net10429;
wire net10159;
wire net782;
wire net1690;
wire net52;
wire net1692;
wire net2092;
wire net6640;
wire net1698;
wire net439;
wire net5000;
wire net5950;
wire net605;
wire out3;
wire net2484;
wire net10331;
wire net3296;
wire net6965;
wire net1706;
wire net6039;
wire net7952;
wire net1709;
wire net692;
wire net6385;
wire net3713;
wire net7979;
wire net3716;
wire net4352;
wire net4398;
wire net1667;
wire net3717;
wire net3259;
wire net3719;
wire net1246;
wire net5799;
wire net3720;
wire net543;
wire net3722;
wire net1599;
wire net3772;
wire net9031;
wire net4657;
wire net1247;
wire net5494;
wire net982;
wire net7423;
wire net4796;
wire net3723;
wire net5843;
wire net3725;
wire net5002;
wire net3727;
wire net3728;
wire net6862;
wire net3730;
wire net10054;
wire net9172;
wire net3731;
wire net5967;
wire net3732;
wire net3734;
wire net9042;
wire net3735;
wire net2432;
wire net4071;
wire net2127;
wire net3736;
wire net9254;
wire net3739;
wire net8315;
wire net4087;
wire net8813;
wire net5849;
wire net8031;
wire net1866;
wire net5656;
wire net3740;
wire net3741;
wire net9864;
wire net9070;
wire net9009;
wire net1758;
wire net3743;
wire net9827;
wire net3744;
wire net3222;
wire net260;
wire net3748;
wire net7774;
wire net6023;
wire net3749;
wire net4163;
wire net1356;
wire net3754;
wire net3756;
wire net6639;
wire net1616;
wire net7130;
wire net3757;
wire net3758;
wire net3715;
wire net7458;
wire net1187;
wire net3759;
wire net3763;
wire net3764;
wire net8499;
wire net8446;
wire net3766;
wire net10466;
wire net6661;
wire net3767;
wire net3774;
wire net4178;
wire net3776;
wire net5208;
wire net7120;
wire net5782;
wire net1444;
wire net6655;
wire net3779;
wire net3918;
wire net2336;
wire net3780;
wire net3783;
wire net3786;
wire net8483;
wire net1242;
wire net3787;
wire net3928;
wire net3788;
wire net3789;
wire net3265;
wire net1211;
wire net4874;
wire net6048;
wire net8214;
wire net4014;
wire net6449;
wire net4736;
wire net7576;
wire net3301;
wire net3796;
wire net5173;
wire net4735;
wire net2328;
wire net7142;
wire net3798;
wire net3799;
wire net3800;
wire net3801;
wire net3807;
wire net9977;
wire net6492;
wire net3809;
wire net4665;
wire net1086;
wire net3810;
wire net7347;
wire net3812;
wire net5376;
wire net3814;
wire net6329;
wire net3433;
wire net3817;
wire net7000;
wire net3818;
wire net3819;
wire net6335;
wire net3820;
wire net3821;
wire net10531;
wire net3822;
wire net8233;
wire net3826;
wire net5092;
wire net3827;
wire net10111;
wire net9762;
wire net4103;
wire net3828;
wire net7766;
wire net3829;
wire net3846;
wire net3830;
wire net6473;
wire net3833;
wire net2907;
wire net6026;
wire net3834;
wire net3837;
wire net2986;
wire net6387;
wire net3653;
wire net3839;
wire net3840;
wire net3841;
wire net4782;
wire net5613;
wire net3842;
wire net716;
wire net3844;
wire net7817;
wire net3847;
wire net3824;
wire net4951;
wire net2713;
wire net3849;
wire net40;
wire net6172;
wire net3851;
wire net3853;
wire net3854;
wire net9441;
wire net4408;
wire net3855;
wire net3857;
wire net3861;
wire net3862;
wire net3864;
wire net9531;
wire net3866;
wire net7778;
wire net4510;
wire net3867;
wire net3868;
wire net3869;
wire net9433;
wire net3870;
wire net5140;
wire net3871;
wire net4967;
wire net1195;
wire net6142;
wire net3872;
wire net3874;
wire net5704;
wire net4161;
wire net3437;
wire net3875;
wire net8548;
wire net2922;
wire net1783;
wire net3877;
wire net7940;
wire net3878;
wire net10501;
wire net3879;
wire net3880;
wire net5158;
wire net10057;
wire net7808;
wire net3598;
wire net3882;
wire net1053;
wire net3888;
wire net3629;
wire net3889;
wire net3891;
wire net3893;
wire net8098;
wire net465;
wire net1860;
wire net3894;
wire net3895;
wire net9297;
wire net8664;
wire net2418;
wire net3902;
wire net7444;
wire net3555;
wire net3903;
wire net3904;
wire net7987;
wire net3905;
wire net5080;
wire net3906;
wire net9808;
wire net4016;
wire net3907;
wire net5530;
wire net3909;
wire net4811;
wire net8375;
wire net7773;
wire net3910;
wire net3911;
wire net5649;
wire net3912;
wire net3916;
wire net4733;
wire net6124;
wire net5456;
wire net5496;
wire net6298;
wire net6578;
wire net9219;
wire net3917;
wire net7071;
wire net3919;
wire net3272;
wire net3922;
wire net5664;
wire net6731;
wire net3924;
wire net1354;
wire net3926;
wire net3929;
wire net8804;
wire net3931;
wire net1216;
wire net1750;
wire net1753;
wire net3932;
wire net1532;
wire net6073;
wire net3934;
wire net3936;
wire net5578;
wire net8604;
wire net3937;
wire net9447;
wire net3664;
wire net3938;
wire net3940;
wire net900;
wire net3941;
wire net10112;
wire net1193;
wire net4764;
wire net3943;
wire net3946;
wire net3947;
wire net3948;
wire net3951;
wire net3952;
wire net3953;
wire net3956;
wire net3957;
wire net9477;
wire net3959;
wire net3963;
wire net6043;
wire net3966;
wire net5412;
wire net6787;
wire net3968;
wire net5007;
wire net3971;
wire net419;
wire net3974;
wire net9196;
wire net3975;
wire net4235;
wire net6046;
wire net3978;
wire net1515;
wire net4186;
wire net9345;
wire net5622;
wire net3981;
wire net10536;
wire net3982;
wire net1936;
wire net3985;
wire net3986;
wire net3991;
wire net3992;
wire net7170;
wire net2282;
wire net3993;
wire net3994;
wire net6120;
wire net3996;
wire net3997;
wire net6358;
wire net3998;
wire net7947;
wire net3706;
wire net4089;
wire net3999;
wire net8089;
wire net2828;
wire net4003;
wire net2490;
wire net6403;
wire net4109;
wire net5126;
wire net4005;
wire net6630;
wire net4007;
wire net4008;
wire net9754;
wire net8376;
wire net4012;
wire net46;
wire net4018;
wire net6543;
wire net4020;
wire net7435;
wire net4021;
wire net4926;
wire net4022;
wire net5900;
wire net1135;
wire net4024;
wire net4580;
wire net6072;
wire net8061;
wire net4027;
wire net6510;
wire net539;
wire net5386;
wire net7047;
wire net4028;
wire net4030;
wire net4031;
wire net4033;
wire net4036;
wire net4037;
wire net4820;
wire net6998;
wire net4038;
wire net4040;
wire net4042;
wire net666;
wire net4043;
wire net4276;
wire net4045;
wire net1917;
wire net5743;
wire net9354;
wire net5164;
wire net994;
wire net4046;
wire net4049;
wire net9549;
wire net8630;
wire net7611;
wire net4051;
wire net4052;
wire net6427;
wire net4053;
wire net4055;
wire net8562;
wire net4057;
wire net4059;
wire net8687;
wire net6422;
wire net658;
wire net5503;
wire net4061;
wire net4062;
wire net5685;
wire net7065;
wire net4064;
wire net4084;
wire net8872;
wire net790;
wire net4065;
wire net6176;
wire net7839;
wire net6634;
wire net4066;
wire net565;
wire net4067;
wire net4069;
wire net8334;
wire net2310;
wire net4070;
wire net6541;
wire net4073;
wire net4680;
wire net6322;
wire net4077;
wire net7664;
wire net907;
wire net150;
wire net4078;
wire net4080;
wire net4082;
wire net9566;
wire net4083;
wire net8162;
wire net2623;
wire net4090;
wire net5299;
wire net4091;
wire net10106;
wire net9072;
wire net4719;
wire net4093;
wire net5948;
wire net4095;
wire out24;
wire net4728;
wire net4101;
wire net8008;
wire net4434;
wire net5227;
wire net6448;
wire net5991;
wire net6763;
wire net5088;
wire net4105;
wire net1423;
wire net4106;
wire net4112;
wire net4114;
wire net7230;
wire net4117;
wire net3724;
wire net4119;
wire net4123;
wire net3425;
wire net5469;
wire net5321;
wire net6866;
wire net2358;
wire net4125;
wire net4126;
wire net4127;
wire net10113;
wire net5769;
wire net4129;
wire net4131;
wire net9562;
wire net4132;
wire net4136;
wire net3038;
wire net4140;
wire net7838;
wire net2465;
wire net4141;
wire net4142;
wire net82;
wire net4144;
wire net8533;
wire net1134;
wire net4145;
wire net4146;
wire net4147;
wire net1235;
wire net5116;
wire net2984;
wire net4150;
wire net8059;
wire net4152;
wire net7951;
wire net2786;
wire net5389;
wire net410;
wire net4155;
wire net449;
wire net7344;
wire net4160;
wire net4164;
wire net3087;
wire net4165;
wire net1142;
wire net4168;
wire net3156;
wire net4169;
wire net1417;
wire net2185;
wire net4171;
wire net5230;
wire net4173;
wire net4177;
wire net2511;
wire net4182;
wire net7831;
wire net6506;
wire net10172;
wire net148;
wire net4183;
wire net4187;
wire net5074;
wire net4189;
wire net6649;
wire net9271;
wire net5071;
wire net4192;
wire net3901;
wire net6993;
wire net4193;
wire net497;
wire net4194;
wire net8116;
wire net6255;
wire net7270;
wire net4197;
wire net2027;
wire net4198;
wire net9998;
wire net4199;
wire net10137;
wire net4265;
wire net8424;
wire net6310;
wire net4203;
wire net4205;
wire net4207;
wire net4208;
wire net1701;
wire net4209;
wire net3564;
wire net5302;
wire net5423;
wire net2768;
wire net4212;
wire net4217;
wire net4221;
wire net3328;
wire net4222;
wire net4648;
wire net235;
wire net5990;
wire net4223;
wire net8094;
wire net4224;
wire net917;
wire net4226;
wire net4227;
wire net4228;
wire net4232;
wire net4233;
wire net5207;
wire net3729;
wire net4237;
wire net4240;
wire net4241;
wire net2218;
wire net7189;
wire net4245;
wire net6204;
wire net9656;
wire net4246;
wire net2965;
wire net5198;
wire net4247;
wire net6125;
wire net4248;
wire net6416;
wire net4249;
wire net4251;
wire net6488;
wire net4253;
wire net8657;
wire net4256;
wire net1628;
wire net4258;
wire net6785;
wire net9950;
wire net4259;
wire net5345;
wire net7104;
wire net4262;
wire net8000;
wire net1439;
wire net4263;
wire net3178;
wire net4269;
wire net1566;
wire net4264;
wire net4268;
wire net5434;
wire net4274;
wire net5135;
wire net3243;
wire net342;
wire net4275;
wire net2624;
wire net4278;
wire net54;
wire net4279;
wire net4281;
wire net4631;
wire net4283;
wire net9308;
wire net9262;
wire net4284;
wire net4285;
wire net4286;
wire net4588;
wire net4612;
wire net3319;
wire net4288;
wire net2177;
wire net4289;
wire net4291;
wire net4292;
wire net4294;
wire net4295;
wire net4297;
wire net8135;
wire net4298;
wire net4299;
wire net7079;
wire net4300;
wire net8065;
wire net2587;
wire net4302;
wire net2632;
wire net4826;
wire net1416;
wire net4305;
wire net2024;
wire net5944;
wire net7115;
wire net4311;
wire net6991;
wire net7608;
wire net4314;
wire net8933;
wire net8019;
wire net4491;
wire net4318;
wire net4325;
wire net4625;
wire net4328;
wire net6252;
wire net4331;
wire net7384;
wire net10251;
wire net519;
wire net4157;
wire net4332;
wire net4836;
wire net7256;
wire net4333;
wire net4334;
wire net4335;
wire net6361;
wire net8393;
wire net4339;
wire net7390;
wire net10243;
wire net4340;
wire net3335;
wire net4341;
wire net8141;
wire net5502;
wire net4342;
wire net8797;
wire net4188;
wire net4343;
wire net4970;
wire net4344;
wire net4345;
wire net2322;
wire net5401;
wire net2321;
wire net5049;
wire net10478;
wire net9698;
wire net4349;
wire net4350;
wire net5060;
wire net4351;
wire net7329;
wire net8085;
wire net6504;
wire net4356;
wire net4357;
wire net4358;
wire net2717;
wire net4359;
wire net6894;
wire net5086;
wire net4360;
wire net10554;
wire net7722;
wire net6151;
wire net10462;
wire net4361;
wire net118;
wire net4364;
wire net1121;
wire net4367;
wire net4368;
wire net4369;
wire net4371;
wire net8451;
wire net517;
wire net4375;
wire net7495;
wire net7126;
wire net4376;
wire net6380;
wire net6849;
wire net4377;
wire net1082;
wire net6376;
wire in19;
wire net4379;
wire net4380;
wire net7190;
wire net4381;
wire net7639;
wire net1845;
wire net5429;
wire net4382;
wire net4383;
wire net302;
wire net1740;
wire net4385;
wire net10217;
wire net4000;
wire net4386;
wire net1762;
wire net1679;
wire net4261;
wire net4388;
wire net7815;
wire net5114;
wire net6629;
wire net4392;
wire net4395;
wire net4396;
wire net10512;
wire net4853;
wire net4397;
wire net5100;
wire net5255;
wire net10562;
wire net8171;
wire net4399;
wire net4403;
wire net3897;
wire net6299;
wire net2945;
wire in11;
wire net4405;
wire net4410;
wire net4412;
wire net6539;
wire net4416;
wire net4417;
wire net4418;
wire net4419;
wire net9838;
wire net8285;
wire net6481;
wire net8846;
wire net4421;
wire net2314;
wire net6268;
wire net4423;
wire net4426;
wire net4427;
wire net6436;
wire net4428;
wire net7111;
wire net188;
wire net5529;
wire net4433;
wire net9370;
wire net4436;
wire net10199;
wire net4667;
wire net339;
wire net6821;
wire net4438;
wire net404;
wire out1;
wire net4957;
wire net4442;
wire net369;
wire net2445;
wire net4445;
wire net6758;
wire net4446;
wire net5597;
wire net434;
wire net4448;
wire net4450;
wire net7854;
wire net5388;
wire net6585;
wire net4458;
wire net3482;
wire net4461;
wire net2303;
wire net5589;
wire net1655;
wire net424;
wire net4463;
wire net4464;
wire net7837;
wire net4466;
wire net4467;
wire net4469;
wire net1801;
wire net4471;
wire net4293;
wire net2136;
wire net5912;
wire net1254;
wire net4474;
wire net4476;
wire net4477;
wire net1691;
wire net4478;
wire net4479;
wire net5021;
wire net4481;
wire net5498;
wire net4484;
wire net7430;
wire net4485;
wire net4486;
wire net4490;
wire net5377;
wire net8237;
wire net4492;
wire net6179;
wire net4494;
wire net4496;
wire net173;
wire net4501;
wire net4503;
wire net4637;
wire net3594;
wire net4504;
wire net7382;
wire net4505;
wire net10346;
wire net675;
wire net4506;
wire net5381;
wire net4508;
wire net2551;
wire net5625;
wire net622;
wire net4509;
wire net2947;
wire net4511;
wire net6366;
wire net5926;
wire net4516;
wire net7599;
wire net4522;
wire net4523;
wire net4524;
wire net4525;
wire net8173;
wire net8115;
wire net4526;
wire net2153;
wire net4530;
wire net2306;
wire net4531;
wire net4534;
wire net268;
wire net1534;
wire net5428;
wire net4536;
wire net5347;
wire net4539;
wire net5573;
wire net1487;
wire net4540;
wire net4541;
wire net4543;
wire net5420;
wire net469;
wire net4546;
wire net6560;
wire net4722;
wire net7023;
wire net7332;
wire net4547;
wire net4549;
wire net4550;
wire net4552;
wire net4554;
wire net435;
wire net4555;
wire net5711;
wire net7081;
wire net9599;
wire net4556;
wire net4558;
wire net10077;
wire net508;
wire net4559;
wire net4562;
wire net187;
wire net6668;
wire net4567;
wire net7330;
wire net4569;
wire net6642;
wire net2835;
wire net3206;
wire net4571;
wire net4287;
wire net4572;
wire net4590;
wire net4574;
wire net4575;
wire net7741;
wire net3373;
wire net4576;
wire net4578;
wire net2095;
wire net6916;
wire net1358;
wire net7321;
wire net4581;
wire net5319;
wire net4583;
wire net6245;
wire net9944;
wire net4585;
wire net3823;
wire net4659;
wire net1590;
wire net4587;
wire net3580;
wire net4592;
wire net5728;
wire net1476;
wire net4593;
wire net4594;
wire net4596;
wire net7735;
wire net6534;
wire net4597;
wire net4598;
wire net7356;
wire net4599;
wire net3976;
wire net4600;
wire net4602;
wire net7048;
wire net4604;
wire net5322;
wire net6669;
wire net9886;
wire net2676;
wire net4606;
wire net6958;
wire net30;
wire net4611;
wire net4731;
wire net1890;
wire net4613;
wire net6370;
wire net3781;
wire net4614;
wire net4615;
wire net3709;
wire net4616;
wire net4617;
wire net6732;
wire net10542;
wire net4621;
wire net4626;
wire in0;
wire net6919;
wire net3151;
wire net4627;
wire net6001;
wire net2926;
wire net3777;
wire net6932;
wire net3671;
wire net4628;
wire net1363;
wire net4629;
wire net3645;
wire net4630;
wire net4632;
wire net6084;
wire net4634;
wire net4635;
wire net2417;
wire net4050;
wire net4638;
wire net8045;
wire net4838;
wire net4640;
wire net6930;
wire net4641;
wire net4643;
wire net5043;
wire net1808;
wire net6949;
wire net8586;
wire net6572;
wire net4651;
wire net4654;
wire net4655;
wire net9372;
wire net7964;
wire net4656;
wire net5752;
wire net4660;
wire net8182;
wire net4752;
wire net4661;
wire net7419;
wire net4662;
wire net8181;
wire net4663;
wire net4664;
wire net4669;
wire net6152;
wire net4670;
wire net8072;
wire net222;
wire net4672;
wire net4674;
wire net2797;
wire net4675;
wire net4676;
wire net1915;
wire net4677;
wire net4678;
wire net4679;
wire net1274;
wire net4682;
wire net2288;
wire net4686;
wire net4687;
wire net8676;
wire net4688;
wire net4690;
wire net4691;
wire net4755;
wire net8709;
wire net2990;
wire net4693;
wire net4694;
wire net9348;
wire net3700;
wire net4644;
wire net4695;
wire net9468;
wire net4697;
wire net4698;
wire net9340;
wire net4699;
wire net4701;
wire net7827;
wire net4702;
wire net4703;
wire net7273;
wire net6987;
wire net4705;
wire net992;
wire net4707;
wire net8500;
wire net4711;
wire net4366;
wire net5355;
wire net4712;
wire net4713;
wire net6320;
wire net4714;
wire net1088;
wire net218;
wire net4715;
wire net4257;
wire net4716;
wire net4717;
wire net3264;
wire net5742;
wire net4720;
wire net8807;
wire net2751;
wire net4999;
wire net4721;
wire net7720;
wire net4048;
wire net6839;
wire net5161;
wire net4723;
wire net4724;
wire net4725;
wire net4726;
wire net4727;
wire net7676;
wire net4729;
wire net4730;
wire net3990;
wire net6978;
wire net4732;
wire net4734;
wire net7237;
wire net4739;
wire net4740;
wire net4743;
wire net1933;
wire net2850;
wire net4102;
wire net4744;
wire net4746;
wire net4882;
wire net4166;
wire net4749;
wire net4751;
wire net2998;
wire net4753;
wire net4758;
wire net6067;
wire net4835;
wire net4760;
wire net2606;
wire net4761;
wire net4355;
wire net6393;
wire net4762;
wire net9964;
wire net4765;
wire net9198;
wire net5598;
wire net4767;
wire net1117;
wire net4769;
wire net743;
wire net4770;
wire net6936;
wire net5190;
wire net4771;
wire net4772;
wire net4404;
wire net4432;
wire net6470;
wire net4009;
wire net4776;
wire net4777;
wire net10029;
wire net7995;
wire net7094;
wire net7718;
wire net4778;
wire net4271;
wire net6410;
wire net1106;
wire net4780;
wire net9627;
wire net4783;
wire net4784;
wire net4785;
wire net4430;
wire net4786;
wire net4788;
wire net4791;
wire net4792;
wire net2366;
wire net1543;
wire net4795;
wire net4797;
wire net289;
wire net4800;
wire net2808;
wire net4801;
wire net4805;
wire net4324;
wire net7028;
wire net4806;
wire net4807;
wire net2771;
wire net6437;
wire net740;
wire net4809;
wire net6482;
wire net10354;
wire net470;
wire net4810;
wire net4814;
wire net4816;
wire net4822;
wire net5564;
wire net4823;
wire net4824;
wire net4519;
wire net4825;
wire net4827;
wire net4829;
wire net6016;
wire net4830;
wire net9223;
wire net6438;
wire net4831;
wire net2367;
wire net4834;
wire net6417;
wire net4837;
wire net10115;
wire net4845;
wire net5287;
wire net3161;
wire net5986;
wire net6432;
wire net3690;
wire net4214;
wire net4848;
wire net4850;
wire net4851;
wire net4548;
wire net5384;
wire net8847;
wire net4857;
wire net4858;
wire net4860;
wire net4861;
wire net4862;
wire net1517;
wire net4864;
wire net4865;
wire net4867;
wire net509;
wire net4870;
wire net4871;
wire net8415;
wire net4872;
wire net1521;
wire net5129;
wire net9540;
wire net1932;
wire net4817;
wire net4875;
wire net5182;
wire net6699;
wire net4876;
wire net10157;
wire net4877;
wire net4879;
wire net4880;
wire net9920;
wire net4883;
wire net720;
wire net4885;
wire net4886;
wire net4887;
wire net9532;
wire net4888;
wire net7461;
wire net4889;
wire net7941;
wire net4891;
wire net8333;
wire net4892;
wire net9201;
wire net5730;
wire net6059;
wire net8431;
wire net4894;
wire net4895;
wire net4897;
wire net4092;
wire net4898;
wire net6345;
wire net4900;
wire net2433;
wire net4903;
wire net3205;
wire net4905;
wire net4906;
wire net5635;
wire net4909;
wire net6191;
wire net1675;
wire net5118;
wire net5154;
wire net6915;
wire net4912;
wire net7060;
wire net4914;
wire net7388;
wire net4916;
wire net184;
wire net4918;
wire net6687;
wire net4919;
wire net7888;
wire net4277;
wire net5485;
wire net9939;
wire net9359;
wire net7512;
wire net4920;
wire net5176;
wire net4921;
wire net9242;
wire net4923;
wire net4925;
wire net4928;
wire net8160;
wire net5847;
wire net6242;
wire net4929;
wire net2194;
wire net4932;
wire net5937;
wire net2341;
wire net4934;
wire net6550;
wire net7578;
wire net4935;
wire net4518;
wire net4936;
wire net4938;
wire net4940;
wire net8324;
wire net4941;
wire net2615;
wire net6917;
wire net4942;
wire net4943;
wire net5581;
wire net7210;
wire net4946;
wire net2961;
wire net745;
wire net4149;
wire net6738;
wire net4947;
wire net4950;
wire net4952;
wire net5111;
wire net4953;
wire net4954;
wire net299;
wire net4956;
wire net6887;
wire net4963;
wire net10450;
wire net4965;
wire net9849;
wire net6681;
wire net7099;
wire net10093;
wire net7312;
wire net4794;
wire net5444;
wire net1325;
wire net4966;
wire net353;
wire net4968;
wire net5995;
wire net4969;
wire net4974;
wire net4977;
wire net683;
wire net7247;
wire net4980;
wire net5342;
wire net4981;
wire net2281;
wire net4982;
wire net6658;
wire net6674;
wire net4983;
wire net4985;
wire net875;
wire net4986;
wire net4989;
wire net6933;
wire net5282;
wire net6486;
wire net4992;
wire net8936;
wire net4994;
wire net647;
wire net7043;
wire net4995;
wire net4997;
wire net6323;
wire net8163;
wire net6300;
wire net4115;
wire net5001;
wire net7886;
wire net5606;
wire net3018;
wire net5003;
wire net6426;
wire net2744;
wire net5006;
wire net9319;
wire net5008;
wire net5011;
wire net4013;
wire net5012;
wire net5014;
wire net4242;
wire net5015;
wire net10352;
wire net4902;
wire net5018;
wire net8566;
wire net5239;
wire net420;
wire net6304;
wire net7293;
wire net41;
wire net5020;
wire net6804;
wire net5023;
wire net3357;
wire net3674;
wire net5028;
wire net10038;
wire net2179;
wire net5029;
wire net9736;
wire net9706;
wire net5032;
wire net5033;
wire net5034;
wire net1539;
wire net5035;
wire net5039;
wire net5041;
wire net303;
wire net6180;
wire net5045;
wire net5046;
wire net5047;
wire net5050;
wire net5051;
wire net5056;
wire net4561;
wire net5063;
wire net7263;
wire net6409;
wire net8351;
wire net6540;
wire net3930;
wire net3792;
wire net7433;
wire net5226;
wire net6981;
wire net5073;
wire net5076;
wire net10502;
wire net5078;
wire net5807;
wire net6163;
wire net5079;
wire net5082;
wire net5083;
wire net7736;
wire net5793;
wire net5085;
wire net5089;
wire net9895;
wire net5094;
wire net6646;
wire net5096;
wire net7460;
wire net950;
wire net5101;
wire net5545;
wire net2598;
wire net4201;
wire net5104;
wire net5107;
wire net5109;
wire net8622;
wire net8581;
wire net5113;
wire net5234;
wire net7432;
wire net7747;
wire net548;
wire net5115;
wire net4029;
wire net5233;
wire net5120;
wire net1810;
wire net5121;
wire net5122;
wire net3287;
wire net5124;
wire net5125;
wire net7689;
wire net5127;
wire net5128;
wire net10013;
wire net6132;
wire net7279;
wire net580;
wire net5130;
wire net9837;
wire net5133;
wire net5134;
wire net10133;
wire net5136;
wire net5137;
wire net6913;
wire net1605;
wire net5138;
wire net3677;
wire net5139;
wire net1612;
wire net5141;
wire net39;
wire net5142;
wire net9498;
wire net5103;
wire net5143;
wire net5144;
wire net5145;
wire net7073;
wire net4195;
wire net5146;
wire net5149;
wire net6961;
wire net9329;
wire net820;
wire net5150;
wire net5151;
wire net5155;
wire net5160;
wire net5162;
wire net9817;
wire net2273;
wire net5163;
wire net5296;
wire net6698;
wire net5168;
wire net9539;
wire net5169;
wire net7844;
wire net814;
wire net5707;
wire net5170;
wire net5171;
wire net5174;
wire net5175;
wire net6844;
wire net6081;
wire net1111;
wire net5179;
wire net10139;
wire net5181;
wire net5185;
wire net5188;
wire net8154;
wire net5189;
wire net5196;
wire net8401;
wire net5197;
wire net8955;
wire net8670;
wire net5201;
wire net6759;
wire net5203;
wire net5204;
wire net2130;
wire net5205;
wire net5206;
wire net1166;
wire net5209;
wire net2910;
wire net6890;
wire net5212;
wire net7976;
wire net6292;
wire net5213;
wire net5219;
wire net5223;
wire net9945;
wire net6112;
wire net206;
wire net2812;
wire net363;
wire net5228;
wire net2483;
wire net6875;
wire net3136;
wire net5232;
wire net5907;
wire net7206;
wire net2467;
wire net5237;
wire net5240;
wire net6362;
wire net4959;
wire net6119;
wire net1779;
wire net5241;
wire net253;
wire net5244;
wire net5246;
wire net5249;
wire net9189;
wire net5251;
wire net1966;
wire net5252;
wire net7037;
wire net5254;
wire net4424;
wire net5256;
wire net5259;
wire net3353;
wire net4308;
wire net5260;
wire net7398;
wire net5266;
wire net10298;
wire net5270;
wire net5273;
wire net7288;
wire net6106;
wire net5275;
wire net6333;
wire net4595;
wire net5276;
wire out25;
wire net7649;
wire net5677;
wire net5280;
wire net8294;
wire net5281;
wire net5286;
wire net2837;
wire net5994;
wire net5290;
wire net1445;
wire net6386;
wire net1038;
wire net5291;
wire net6525;
wire net6164;
wire net5297;
wire net5298;
wire net8515;
wire net4473;
wire net5068;
wire net5300;
wire net5301;
wire net10213;
wire net5304;
wire net5830;
wire net5307;
wire net4878;
wire net5310;
wire net5311;
wire net2300;
wire net3794;
wire net7265;
wire net9400;
wire net5314;
wire net6536;
wire net5317;
wire net3123;
wire net5320;
wire net1979;
wire net6193;
wire net5323;
wire net3825;
wire net5324;
wire net6901;
wire net5325;
wire net5327;
wire net9094;
wire net3025;
wire net5813;
wire net5328;
wire net5331;
wire net9996;
wire net5333;
wire net5835;
wire net5334;
wire net9719;
wire net355;
wire net5336;
wire net5337;
wire net8999;
wire net8879;
wire net5338;
wire net5339;
wire net1815;
wire net5340;
wire net5627;
wire net5224;
wire net7195;
wire net5557;
wire net5773;
wire net5352;
wire net4502;
wire net5353;
wire net5356;
wire net2196;
wire net6211;
wire net5357;
wire net10427;
wire net4100;
wire net5717;
wire net6232;
wire net9572;
wire net5359;
wire net5615;
wire net5361;
wire net5364;
wire net8435;
wire net531;
wire net1764;
wire net5365;
wire net6631;
wire net5366;
wire net5370;
wire net7203;
wire net5374;
wire net5383;
wire net5385;
wire net5390;
wire net5391;
wire net6659;
wire net5393;
wire net5395;
wire net5398;
wire net4704;
wire net5402;
wire net5404;
wire net1535;
wire net5405;
wire net5408;
wire net5413;
wire net5416;
wire net5417;
wire net5418;
wire net1015;
wire net5419;
wire net26;
wire net5424;
wire net10402;
wire net5425;
wire net5426;
wire net5433;
wire net681;
wire net5435;
wire net5437;
wire net5439;
wire net10484;
wire net5775;
wire net5441;
wire net5442;
wire net10284;
wire net5445;
wire net9527;
wire net5448;
wire net5450;
wire net2925;
wire net5451;
wire net4976;
wire net5452;
wire net7283;
wire net5453;
wire net6626;
wire net104;
wire net5454;
wire net4472;
wire net5459;
wire net6216;
wire net6463;
wire net5461;
wire net5072;
wire net5462;
wire net5466;
wire net5467;
wire net5468;
wire net8491;
wire net7445;
wire net319;
wire net5535;
wire net5470;
wire net5471;
wire net6212;
wire net5472;
wire net5475;
wire net5476;
wire net5477;
wire net7316;
wire net5478;
wire net6867;
wire net6295;
wire net1049;
wire net5479;
wire net5486;
wire net5487;
wire net3020;
wire net850;
wire net1505;
wire net5489;
wire net5490;
wire net5491;
wire net9169;
wire net6140;
wire net5495;
wire net5500;
wire net5501;
wire net6617;
wire net5505;
wire net5506;
wire net9867;
wire net1156;
wire net5509;
wire net9728;
wire net5618;
wire net6800;
wire net10004;
wire net5510;
wire net5511;
wire net5513;
wire net1972;
wire net5514;
wire net9230;
wire net9179;
wire net5920;
wire net5515;
wire net5516;
wire net5517;
wire net1719;
wire net5522;
wire net2462;
wire net2059;
wire net1873;
wire net5523;
wire net5526;
wire net5527;
wire net5528;
wire net7464;
wire net5531;
wire net3896;
wire net7289;
wire net5532;
wire net6032;
wire net6407;
wire net2181;
wire net5534;
wire net5537;
wire net352;
wire net5540;
wire net4624;
wire net5541;
wire net5542;
wire net5543;
wire net5544;
wire net5547;
wire net5550;
wire net5551;
wire net3942;
wire net5552;
wire net5562;
wire net1312;
wire net5565;
wire net5566;
wire net5567;
wire net5809;
wire net7336;
wire net5942;
wire net7438;
wire net5571;
wire net111;
wire net5574;
wire net947;
wire net5575;
wire net5157;
wire net5295;
wire net5580;
wire net4210;
wire net5584;
wire net10477;
wire net5585;
wire net4779;
wire net6071;
wire net5587;
wire net5591;
wire net6742;
wire net5592;
wire net5593;
wire net9897;
wire net5595;
wire net1309;
wire net5596;
wire net10021;
wire net7835;
wire net1869;
wire net5600;
wire net5106;
wire net5504;
wire net5601;
wire net6230;
wire net5604;
wire net5605;
wire net7090;
wire net9476;
wire net5608;
wire net3506;
wire net562;
wire net267;
wire net1324;
wire net5611;
wire net4435;
wire net5616;
wire net7620;
wire net5619;
wire net3456;
wire net5620;
wire net5059;
wire net5623;
wire net5631;
wire net5636;
wire net5640;
wire net2168;
wire net1699;
wire net5641;
wire net7829;
wire net2843;
wire net119;
wire net5642;
wire net568;
wire net5643;
wire net9163;
wire net918;
wire net5644;
wire net5646;
wire net1824;
wire net3261;
wire net5650;
wire net8443;
wire net5651;
wire net5652;
wire net6884;
wire net5653;
wire net5654;
wire net5655;
wire net5657;
wire net6440;
wire net5658;
wire net8559;
wire net2166;
wire net5659;
wire net5662;
wire net6037;
wire net4365;
wire net7001;
wire net4642;
wire net5663;
wire net5665;
wire net7455;
wire net5666;
wire net5671;
wire net7532;
wire net5052;
wire net5672;
wire net32;
wire net5676;
wire net769;
wire net5679;
wire net10366;
wire net3497;
wire net3404;
wire net5684;
wire net5687;
wire net5770;
wire net5691;
wire net6623;
wire net3659;
wire net5693;
wire net5694;
wire net8848;
wire net4913;
wire net5698;
wire net6213;
wire net5804;
wire net5215;
wire net6653;
wire net5703;
wire net1872;
wire net5705;
wire net9559;
wire net2373;
wire net7174;
wire net7807;
wire net865;
wire net5706;
wire net5708;
wire net2443;
wire net5710;
wire net6819;
wire net266;
wire net5713;
wire net5714;
wire net4480;
wire net4991;
wire net5715;
wire net5716;
wire net8250;
wire net3804;
wire net6169;
wire net5718;
wire net5720;
wire net232;
wire net5721;
wire net5722;
wire net5723;
wire net5725;
wire net5726;
wire net6183;
wire net5729;
wire net9307;
wire net6842;
wire net5731;
wire net5632;
wire net5903;
wire net1128;
wire net4544;
wire net6564;
wire net5732;
wire net7348;
wire net5734;
wire net9135;
wire net5736;
wire net5737;
wire net5738;
wire net5740;
wire net8540;
wire net4623;
wire net5744;
wire net5747;
wire net6686;
wire net9334;
wire net7057;
wire net3313;
wire net5750;
wire net5751;
wire net5754;
wire net3256;
wire net5755;
wire net5757;
wire net590;
wire net5760;
wire net5761;
wire net8373;
wire net7557;
wire net5316;
wire net5762;
wire net6834;
wire net9846;
wire net5763;
wire net2607;
wire net7272;
wire net3483;
wire net2635;
wire net1995;
wire net5766;
wire net6253;
wire net5772;
wire net5777;
wire net8800;
wire net5781;
wire net7323;
wire net5783;
wire net6845;
wire net7187;
wire net5785;
wire net7885;
wire net2013;
wire net5786;
wire net4420;
wire net5787;
wire net5788;
wire net7819;
wire net5791;
wire net5796;
wire net5797;
wire net2898;
wire net5798;
wire net5915;
wire net5802;
wire net7739;
wire net5054;
wire net6790;
wire net1154;
wire net5803;
wire net5810;
wire net2860;
wire net5811;
wire net708;
wire net2739;
wire net5739;
wire net6413;
wire net10163;
wire net5812;
wire net5817;
wire net6049;
wire net5818;
wire net5819;
wire net9794;
wire net7284;
wire net2319;
wire net5821;
wire net7025;
wire net1474;
wire net5822;
wire net8561;
wire net2748;
wire net5824;
wire net5825;
wire net5826;
wire net5828;
wire net2286;
wire net5831;
wire net2862;
wire net5004;
wire net5832;
wire net5836;
wire net6822;
wire net5840;
wire net156;
wire net5842;
wire net1662;
wire net6516;
wire net5844;
wire net5805;
wire net6977;
wire net5846;
wire net3477;
wire net5850;
wire net2420;
wire net5851;
wire net764;
wire net5852;
wire net7400;
wire net10481;
wire net3223;
wire net5854;
wire net5855;
wire net4706;
wire net5856;
wire net7117;
wire net5857;
wire net5859;
wire net5860;
wire net6155;
wire net5861;
wire net5274;
wire net5862;
wire net5865;
wire net5870;
wire net5871;
wire net5872;
wire net5873;
wire net4322;
wire net5875;
wire net6695;
wire net124;
wire net4890;
wire net5880;
wire net1787;
wire net5888;
wire net8053;
wire net5153;
wire net7024;
wire net9811;
wire net1953;
wire net7454;
wire net5894;
wire net6812;
wire net5895;
wire net1880;
wire net5896;
wire net5897;
wire net1058;
wire net5898;
wire net8476;
wire net5853;
wire net5899;
wire net1377;
wire net5901;
wire net5902;
wire net3765;
wire net5904;
wire net8522;
wire net5905;
wire net5909;
wire net4873;
wire net5910;
wire net400;
wire net5911;
wire net5916;
wire net1847;
wire net5917;
wire net5918;
wire net5919;
wire net5921;
wire net5922;
wire net8697;
wire net7118;
wire net5923;
wire net5927;
wire net6279;
wire net5929;
wire net2017;
wire net5931;
wire net5932;
wire net9834;
wire net5934;
wire net3708;
wire net5935;
wire net2901;
wire net6693;
wire net5938;
wire net9697;
wire net5939;
wire net5414;
wire net305;
wire net5940;
wire net5945;
wire net7093;
wire net5949;
wire net7602;
wire net5261;
wire net5951;
wire net7389;
wire net9078;
wire net840;
wire net5954;
wire net5753;
wire net5955;
wire net6371;
wire net5956;
wire net1649;
wire net1464;
wire net5957;
wire net5958;
wire net7978;
wire net2590;
wire net5959;
wire net8883;
wire net5960;
wire net9140;
wire net3540;
wire net6471;
wire net10397;
wire net5962;
wire net1123;
wire net5964;
wire net6928;
wire net10110;
wire net1919;
wire net5969;
wire net9120;
wire net6865;
wire net5970;
wire out13;
wire net6189;
wire net9542;
wire net5971;
wire net5972;
wire net5973;
wire net2582;
wire net5975;
wire net2957;
wire net3816;
wire net5978;
wire net5979;
wire net2912;
wire net5981;
wire net6988;
wire net5982;
wire net754;
wire net5983;
wire net5985;
wire net5988;
wire net5992;
wire net9902;
wire net9815;
wire net2183;
wire net6556;
wire net5996;
wire net3213;
wire net6996;
wire net5998;
wire net6000;
wire net6005;
wire net6007;
wire net7421;
wire net2044;
wire net1752;
wire net1949;
wire net6008;
wire net6009;
wire net2470;
wire net6010;
wire net10449;
wire net6011;
wire net2851;
wire net6012;
wire net6013;
wire net6014;
wire net1229;
wire net6015;
wire net6018;
wire net2905;
wire net1392;
wire net6020;
wire net6021;
wire net8517;
wire net1825;
wire net6022;
wire net6029;
wire net6030;
wire net6031;
wire net10045;
wire net6290;
wire net5269;
wire net6033;
wire net6034;
wire net8402;
wire net6040;
wire net6041;
wire net9670;
wire net2496;
wire net2052;
wire net6042;
wire net6045;
wire net6047;
wire net6050;
wire net3334;
wire net6051;
wire net6052;
wire net6053;
wire net2611;
wire net4158;
wire net6054;
wire net1061;
wire net6055;
wire net6056;
wire net9458;
wire net6060;
wire net4488;
wire net6061;
wire net4603;
wire net6457;
wire net6512;
wire net5380;
wire net7123;
wire net5329;
wire net6062;
wire net6065;
wire net6066;
wire net6074;
wire net6075;
wire net228;
wire net5178;
wire net6076;
wire net10062;
wire net6078;
wire net6080;
wire net6082;
wire net6083;
wire net6085;
wire net6086;
wire net6143;
wire net2619;
wire net2190;
wire net6087;
wire net6090;
wire net3636;
wire net6091;
wire net4056;
wire net6093;
wire net7175;
wire net431;
wire net6098;
wire net3271;
wire net5231;
wire net6100;
wire net7826;
wire net6101;
wire net1294;
wire net6102;
wire net5409;
wire net6628;
wire net8302;
wire net1527;
wire net6158;
wire net6103;
wire net3051;
wire net6104;
wire net1041;
wire net5250;
wire net6105;
wire net7386;
wire net6108;
wire net6109;
wire net4804;
wire net6110;
wire net1263;
wire net1397;
wire net6111;
wire net6113;
wire net6399;
wire net6117;
wire net1349;
wire net6118;
wire net1352;
wire net6121;
wire net6126;
wire net6127;
wire net6129;
wire net1273;
wire net6130;
wire net1561;
wire net6133;
wire net6134;
wire net6135;
wire net4537;
wire net7213;
wire net6136;
wire net6137;
wire net6138;
wire net6139;
wire net6141;
wire net8176;
wire net6144;
wire net6146;
wire net1070;
wire net6888;
wire net10090;
wire net6154;
wire net7097;
wire net8309;
wire net6162;
wire net6902;
wire net6165;
wire net6167;
wire net7191;
wire net7981;
wire net6289;
wire net6168;
wire net6171;
wire net7299;
wire net7893;
wire net6174;
wire net7903;
wire net7443;
wire net6175;
wire net8258;
wire net6177;
wire net10537;
wire net5110;
wire net6181;
wire net6173;
wire net6182;
wire net10233;
wire net6184;
wire net6185;
wire net10035;
wire net6187;
wire net5474;
wire net1902;
wire net1540;
wire net6190;
wire net2342;
wire net6195;
wire net6196;
wire net9206;
wire net6602;
wire net1715;
wire net6199;
wire net6200;
wire net10457;
wire net6201;
wire net6206;
wire net6208;
wire net9047;
wire net6004;
wire net6209;
wire net7757;
wire net4854;
wire net6210;
wire net6215;
wire net2109;
wire net6217;
wire net3514;
wire net6219;
wire net6220;
wire net6222;
wire net3412;
wire net341;
wire net6223;
wire net6224;
wire net6227;
wire net4134;
wire net6231;
wire net6233;
wire net5016;
wire net6235;
wire net2546;
wire net6259;
wire net6236;
wire net9590;
wire net1728;
wire net6811;
wire net6238;
wire net7682;
wire net6239;
wire net6241;
wire net6243;
wire net6244;
wire net9123;
wire net1537;
wire net5667;
wire net5570;
wire net6246;
wire net7003;
wire net2035;
wire net1529;
wire net6247;
wire net6250;
wire net2158;
wire net6392;
wire net8147;
wire net6254;
wire net6257;
wire net6258;
wire net9888;
wire net5686;
wire net4911;
wire net6260;
wire net6261;
wire net9954;
wire net6262;
wire net8647;
wire net8601;
wire net1345;
wire net6263;
wire net4459;
wire net136;
wire net6265;
wire net4718;
wire net6266;
wire net8307;
wire net6269;
wire net6270;
wire net6271;
wire net6273;
wire net6274;
wire net6276;
wire net9048;
wire net6282;
wire net7846;
wire net6283;
wire net6571;
wire net6284;
wire net6285;
wire net6286;
wire net6899;
wire net6287;
wire net6291;
wire net8783;
wire net1647;
wire net6293;
wire net1807;
wire net6294;
wire net2395;
wire net1891;
wire net6301;
wire net6305;
wire net3012;
wire net6306;
wire net2124;
wire net6918;
wire net6308;
wire net1957;
wire net1096;
wire net2225;
wire net4088;
wire net6309;
wire net2762;
wire net6313;
wire net6314;
wire net9716;
wire net6406;
wire net8349;
wire net6096;
wire net6315;
wire net6317;
wire net6318;
wire net8291;
wire net6319;
wire net6321;
wire net9321;
wire net6325;
wire net2711;
wire net6326;
wire net6327;
wire net8037;
wire net595;
wire net6328;
wire net7125;
wire net6330;
wire net10128;
wire net5081;
wire net6331;
wire net6334;
wire net8180;
wire net6336;
wire net9243;
wire net6338;
wire net4307;
wire net6339;
wire net6341;
wire net8078;
wire net6468;
wire net6342;
wire net6343;
wire net6346;
wire net3583;
wire net2553;
wire net1107;
wire net6347;
wire net6348;
wire net6349;
wire net6352;
wire net6355;
wire net6359;
wire net10443;
wire net6374;
wire net6505;
wire net6364;
wire net7154;
wire net6365;
wire net9413;
wire net427;
wire net6367;
wire net8036;
wire net6369;
wire net8792;
wire net6372;
wire net6375;
wire net6377;
wire net6378;
wire net2051;
wire net6379;
wire net9460;
wire net6382;
wire net6383;
wire net10495;
wire net6384;
wire net6388;
wire net6389;
wire net169;
wire net6391;
wire net10058;
wire net6394;
wire net3131;
wire net6396;
wire net6739;
wire net8224;
wire net6397;
wire net6401;
wire net6402;
wire net6405;
wire net8962;
wire net6408;
wire net6491;
wire net6411;
wire net6753;
wire net6412;
wire net8886;
wire net1004;
wire net6415;
wire net6784;
wire net1047;
wire net6418;
wire net9655;
wire net6420;
wire net7667;
wire net2685;
wire net6903;
wire net6424;
wire net6428;
wire net7002;
wire net687;
wire net1412;
wire net7179;
wire net3742;
wire net6430;
wire net4121;
wire net6433;
wire net3472;
wire net6439;
wire net4270;
wire net6443;
wire net6444;
wire net6445;
wire net9681;
wire net6446;
wire net8246;
wire net5878;
wire net6447;
wire net3750;
wire net4391;
wire net6452;
wire net6453;
wire net6454;
wire net7039;
wire net6456;
wire net6459;
wire net6460;
wire net3385;
wire net6469;
wire net6475;
wire net1898;
wire net6477;
wire net6478;
wire net6479;
wire net1546;
wire net6480;
wire net7717;
wire net7161;
wire net4639;
wire net6487;
wire net6489;
wire net6493;
wire net1140;
wire net6494;
wire net6497;
wire net9471;
wire net6499;
wire net6501;
wire net5431;
wire net6503;
wire net5863;
wire net6535;
wire net6603;
wire net6507;
wire net6508;
wire net5733;
wire net7480;
wire net7542;
wire net6511;
wire net10083;
wire net6513;
wire net6514;
wire net9543;
wire net6515;
wire net6562;
wire net6518;
wire net2963;
wire net6519;
wire net243;
wire net6520;
wire net1390;
wire net6523;
wire net6524;
wire net7709;
wire net4741;
wire net6823;
wire net6527;
wire net6529;
wire net8122;
wire net6077;
wire net6533;
wire net10068;
wire net6538;
wire net6544;
wire net6547;
wire net6552;
wire net2348;
wire net6553;
wire net6554;
wire net6685;
wire net7393;
wire net6557;
wire net5634;
wire net6558;
wire net10010;
wire net2820;
wire net6559;
wire net6561;
wire net6563;
wire net6567;
wire net9102;
wire net1583;
wire net5546;
wire net6568;
wire net10471;
wire net6570;
wire net1102;
wire net6575;
wire net4019;
wire net6577;
wire net1138;
wire net6581;
wire net10459;
wire net10325;
wire net3324;
wire net6582;
wire net9067;
wire net6583;
wire net781;
wire net6599;
wire net6586;
wire net6587;
wire net9702;
wire net6588;
wire net6589;
wire net6202;
wire net6590;
wire net6592;
wire net7534;
wire net6593;
wire net586;
wire net4514;
wire net7391;
wire net5438;
wire net6597;
wire net6605;
wire net6608;
wire net8079;
wire net6609;
wire net6632;
wire net3359;
wire net6610;
wire net6611;
wire net8248;
wire net471;
wire net6613;
wire net6614;
wire net3614;
wire net4538;
wire net6615;
wire net6616;
wire net6620;
wire net4312;
wire net6621;
wire net6624;
wire net6627;
wire net9558;
wire net6633;
wire net6643;
wire net6648;
wire net6650;
wire net9874;
wire net6656;
wire net8490;
wire net6662;
wire net277;
wire net6665;
wire net5869;
wire net6670;
wire net6672;
wire net6675;
wire net6678;
wire net5848;
wire net6679;
wire net6683;
wire net2350;
wire net6688;
wire net4681;
wire net6690;
wire net6694;
wire net6696;
wire net6704;
wire net1337;
wire net827;
wire net6709;
wire net7734;
wire net5484;
wire net4984;
wire net6969;
wire net6710;
wire net8892;
wire net3675;
wire net5065;
wire net6711;
wire net3746;
wire net6713;
wire net10392;
wire net6716;
wire net6719;
wire net2410;
wire net6340;
wire net6722;
wire net6726;
wire net7252;
wire net6728;
wire net5521;
wire net6729;
wire net8757;
wire net6734;
wire net4582;
wire net5187;
wire net6736;
wire net547;
wire net6741;
wire net6746;
wire net6747;
wire net9501;
wire net1198;
wire net6748;
wire net6749;
wire net6750;
wire net3253;
wire net6751;
wire net6752;
wire net3190;
wire net1328;
wire net6754;
wire net10188;
wire net9763;
wire net5220;
wire net6755;
wire net6929;
wire net6756;
wire net6757;
wire net6762;
wire net7334;
wire net5318;
wire net6765;
wire net5968;
wire net6768;
wire net2340;
wire net6769;
wire net7232;
wire net6771;
wire net10373;
wire net6772;
wire net2382;
wire net109;
wire net7437;
wire net6773;
wire net1362;
wire net7146;
wire net6775;
wire net6777;
wire net6778;
wire net987;
wire net7236;
wire net6779;
wire net7050;
wire net6780;
wire net5997;
wire net6781;
wire net6794;
wire net6783;
wire net9664;
wire net165;
wire net4573;
wire net6788;
wire net6789;
wire net7062;
wire net6795;
wire net6207;
wire net6798;
wire net6801;
wire net3079;
wire net6802;
wire net7150;
wire net6803;
wire net6805;
wire net6807;
wire net6808;
wire net1659;
wire net6809;
wire net6814;
wire net6815;
wire net8700;
wire net6099;
wire net6817;
wire net6820;
wire net6825;
wire net4353;
wire net6827;
wire net1782;
wire net6828;
wire net8794;
wire net6829;
wire net1988;
wire net6830;
wire net8583;
wire net6831;
wire net9563;
wire net6833;
wire net6835;
wire net6836;
wire net6837;
wire net806;
wire net6840;
wire net2207;
wire net5795;
wire net6841;
wire net6846;
wire net6847;
wire net6848;
wire net6851;
wire net9024;
wire net6854;
wire net5569;
wire net6855;
wire net6857;
wire net8944;
wire net6859;
wire net151;
wire net6860;
wire net1905;
wire net6863;
wire net540;
wire net6869;
wire net6870;
wire net8052;
wire net1275;
wire net2315;
wire net6871;
wire net6873;
wire net5330;
wire net6874;
wire net1582;
wire net6878;
wire net6880;
wire net9593;
wire net6883;
wire net6886;
wire net6889;
wire net6891;
wire net9832;
wire net325;
wire net56;
wire net6893;
wire net6896;
wire net1794;
wire net6898;
wire net5771;
wire net6900;
wire net2148;
wire net4346;
wire net7375;
wire net6904;
wire net6906;
wire net6910;
wire net705;
wire net6912;
wire net6920;
wire net6925;
wire net10349;
wire net9718;
wire net6926;
wire net6931;
wire net5594;
wire net6935;
wire net4406;
wire net6937;
wire net6938;
wire net6939;
wire net4004;
wire net6942;
wire net1151;
wire net6943;
wire net6944;
wire net4175;
wire net6945;
wire net6947;
wire net399;
wire net6950;
wire net6952;
wire net6953;
wire net2993;
wire net6955;
wire net3863;
wire net6959;
wire net4407;
wire net6962;
wire net6963;
wire net4649;
wire net6964;
wire net2977;
wire net6966;
wire net786;
wire net7114;
wire net6967;
wire net3135;
wire net6970;
wire net2664;
wire net6972;
wire net6974;
wire net6983;
wire net10406;
wire net2682;
wire net6984;
wire net7121;
wire net6027;
wire net6985;
wire net413;
wire net6992;
wire net9842;
wire net7446;
wire net6995;
wire net7580;
wire net3987;
wire net6999;
wire net7004;
wire net8137;
wire net805;
wire net7005;
wire net1239;
wire net7007;
wire net6024;
wire net5211;
wire net7008;
wire net7010;
wire net7012;
wire net7013;
wire net7014;
wire net7017;
wire net7019;
wire net7697;
wire net7228;
wire net10528;
wire net7020;
wire net7027;
wire net7030;
wire net7032;
wire net7033;
wire net7035;
wire net7036;
wire net7038;
wire net2186;
wire net7096;
wire net7040;
wire net9560;
wire net5868;
wire net7041;
wire net7992;
wire net7045;
wire net7049;
wire net7052;
wire net7055;
wire net23;
wire net7056;
wire net7058;
wire net7063;
wire net3501;
wire net3656;
wire net1805;
wire net7064;
wire net9910;
wire net1334;
wire net7066;
wire net7068;
wire net7077;
wire net7083;
wire net4563;
wire net7086;
wire net10273;
wire net304;
wire net7087;
wire net1370;
wire net7088;
wire net5005;
wire net7089;
wire net7091;
wire net7842;
wire net7098;
wire net7325;
wire net3806;
wire net7100;
wire net7105;
wire net7106;
wire net5102;
wire net7108;
wire net9914;
wire net7110;
wire net8565;
wire net7112;
wire net3553;
wire net7113;
wire net7116;
wire net7119;
wire net7128;
wire net7129;
wire net7133;
wire net7783;
wire net2727;
wire net7134;
wire net10441;
wire net7135;
wire net7136;
wire net7138;
wire net10521;
wire net7140;
wire net7141;
wire net7143;
wire net5689;
wire net7144;
wire net7148;
wire net9487;
wire net7149;
wire net7673;
wire net6718;
wire net7152;
wire net9971;
wire net4843;
wire net7157;
wire net1624;
wire net7160;
wire net1320;
wire net7163;
wire net7851;
wire net7164;
wire net7165;
wire net1290;
wire net7167;
wire net5701;
wire net7168;
wire net7169;
wire net7496;
wire net6192;
wire net7171;
wire net1436;
wire net7172;
wire net9216;
wire net7173;
wire net7180;
wire net8535;
wire net7181;
wire net4320;
wire net7186;
wire net322;
wire net7188;
wire net7197;
wire net1176;
wire net7198;
wire net575;
wire net7199;
wire net1109;
wire net7200;
wire net307;
wire net7201;
wire net3733;
wire net7205;
wire net7207;
wire net7208;
wire net7209;
wire net7211;
wire net1708;
wire net7212;
wire net7076;
wire net7214;
wire net7215;
wire net9428;
wire net7217;
wire net7222;
wire net9456;
wire net9109;
wire net7224;
wire net7225;
wire net9835;
wire net7067;
wire net7227;
wire net7229;
wire net9915;
wire net5941;
wire net7233;
wire net9395;
wire net3022;
wire net7234;
wire net8270;
wire net4310;
wire net7238;
wire net7240;
wire net7882;
wire net7243;
wire net5293;
wire net7248;
wire net7251;
wire net7253;
wire net5892;
wire net1812;
wire net7254;
wire net6622;
wire net7255;
wire net5885;
wire net7258;
wire net7264;
wire net7780;
wire net4465;
wire net7266;
wire net7274;
wire net1875;
wire net7275;
wire net6635;
wire net7277;
wire net7280;
wire net7287;
wire out19;
wire net4456;
wire net7291;
wire net9999;
wire net7292;
wire net7297;
wire net7298;
wire net7301;
wire net2987;
wire out8;
wire net1877;
wire net7304;
wire net7305;
wire net9008;
wire net7307;
wire net7308;
wire net3865;
wire net7313;
wire net7317;
wire net9564;
wire net7318;
wire net1680;
wire net7322;
wire net7333;
wire net7337;
wire net9232;
wire net7339;
wire net7340;
wire net7341;
wire net7342;
wire net7343;
wire net7350;
wire net8364;
wire net6521;
wire net7351;
wire net7352;
wire net1430;
wire net7357;
wire net7360;
wire net7362;
wire net7434;
wire net8473;
wire net7365;
wire net7366;
wire net7367;
wire net7574;
wire net3351;
wire net7369;
wire net7371;
wire net5765;
wire net7373;
wire net9495;
wire net7376;
wire net8659;
wire net7377;
wire net7380;
wire net5343;
wire net7383;
wire net1019;
wire net7392;
wire net9546;
wire net7394;
wire net10170;
wire net61;
wire net7395;
wire net7397;
wire net7399;
wire net7401;
wire net9552;
wire net7403;
wire net1781;
wire net7404;
wire net7405;
wire net9472;
wire net7407;
wire net3778;
wire net6161;
wire net4468;
wire net3815;
wire net6116;
wire net7409;
wire net10569;
wire net7411;
wire net7412;
wire net3515;
wire net4566;
wire net7413;
wire net10557;
wire net7420;
wire net6810;
wire net7422;
wire net2063;
wire net3883;
wire net6450;
wire net7424;
wire net4047;
wire net7426;
wire net4244;
wire net7436;
wire net6495;
wire net7153;
wire net7439;
wire net7442;
wire net7447;
wire net5463;
wire net7448;
wire net7449;
wire net7451;
wire net2900;
wire net7452;
wire net7856;
wire net7453;
wire net7456;
wire net7459;
wire net4025;
wire net7468;
wire net7471;
wire net3281;
wire net7472;
wire net7473;
wire net5285;
wire net7474;
wire net7477;
wire net2173;
wire net7478;
wire net3606;
wire net7479;
wire net7482;
BUFx10_ASAP7_75t_R c26(
.A(in20),
.Y(net0)
);

BUFx12_ASAP7_75t_R c27(
.A(in17),
.Y(net1)
);

AND2x2_ASAP7_75t_R c28(
.A(net0),
.B(in11),
.Y(net2)
);

BUFx12f_ASAP7_75t_R c29(
.A(in10),
.Y(net3)
);

AND2x4_ASAP7_75t_R c30(
.A(net3),
.B(in2),
.Y(net4)
);

BUFx16f_ASAP7_75t_R c31(
.A(in8),
.Y(net5)
);

BUFx24_ASAP7_75t_R c32(
.A(in17),
.Y(net6)
);

BUFx2_ASAP7_75t_R c33(
.A(in2),
.Y(net7)
);

AND3x1_ASAP7_75t_R c34(
.A(in21),
.B(in9),
.C(net0),
.Y(net8)
);

BUFx3_ASAP7_75t_R c35(
.A(net8),
.Y(net9)
);

AND2x6_ASAP7_75t_R c36(
.A(in22),
.B(net2),
.Y(net10)
);

BUFx4_ASAP7_75t_R c37(
.A(in3),
.Y(net11)
);

AND3x2_ASAP7_75t_R c38(
.A(net9),
.B(in6),
.C(net41),
.Y(net12)
);

HAxp5_ASAP7_75t_R c39(
.A(net5),
.B(net3),
.CON(net14),
.SN(net13)
);

NAND2x1_ASAP7_75t_R c40(
.A(net40),
.B(net2),
.Y(net15)
);

AND3x4_ASAP7_75t_R c41(
.A(net7),
.B(in0),
.C(in12),
.Y(net16)
);

BUFx4f_ASAP7_75t_R c42(
.A(net10),
.Y(net17)
);

BUFx5_ASAP7_75t_R c43(
.A(in15),
.Y(net18)
);

BUFx6f_ASAP7_75t_R c44(
.A(net40),
.Y(net19)
);

BUFx8_ASAP7_75t_R c45(
.A(in6),
.Y(net20)
);

CKINVDCx10_ASAP7_75t_R c46(
.A(net18),
.Y(net21)
);

NAND2x1p5_ASAP7_75t_R c47(
.A(net19),
.B(net40),
.Y(net22)
);

CKINVDCx11_ASAP7_75t_R c48(
.A(net15),
.Y(net23)
);

CKINVDCx12_ASAP7_75t_R c49(
.A(net23),
.Y(net24)
);

CKINVDCx14_ASAP7_75t_R c50(
.A(net3),
.Y(net25)
);

CKINVDCx16_ASAP7_75t_R c51(
.A(net8),
.Y(net26)
);

NAND2x2_ASAP7_75t_R c52(
.A(in0),
.B(net2),
.Y(net27)
);

CKINVDCx20_ASAP7_75t_R c53(
.A(net24),
.Y(net28)
);

CKINVDCx5p33_ASAP7_75t_R c54(
.A(net1),
.Y(net29)
);

AO21x1_ASAP7_75t_R c55(
.A1(net24),
.A2(net28),
.B(net19),
.Y(net30)
);

CKINVDCx6p67_ASAP7_75t_R c56(
.A(net29),
.Y(net31)
);

CKINVDCx8_ASAP7_75t_R c57(
.A(net21),
.Y(net32)
);

AO21x2_ASAP7_75t_R c58(
.A1(net14),
.A2(net1),
.B(net32),
.Y(net33)
);

NAND2xp33_ASAP7_75t_R c59(
.A(net31),
.B(net30),
.Y(net34)
);

AOI21x1_ASAP7_75t_R c60(
.A1(net27),
.A2(net31),
.B(net34),
.Y(net35)
);

CKINVDCx9p33_ASAP7_75t_R c61(
.A(net12),
.Y(net36)
);

NAND2xp5_ASAP7_75t_R c62(
.A(in22),
.B(net32),
.Y(net37)
);

NAND2xp67_ASAP7_75t_R c63(
.A(net32),
.B(net35),
.Y(net38)
);

HB1xp67_ASAP7_75t_R c64(
.A(in11),
.Y(net39)
);

HB2xp67_ASAP7_75t_R c65(
.A(in1),
.Y(net40)
);

HB3xp67_ASAP7_75t_R c66(
.A(in16),
.Y(net41)
);

AOI21xp33_ASAP7_75t_R c67(
.A1(net35),
.A2(in5),
.B(net32),
.Y(net42)
);

AOI21xp5_ASAP7_75t_R c68(
.A1(net2),
.A2(net32),
.B(net3),
.Y(net43)
);

HB4xp67_ASAP7_75t_R c69(
.A(net43),
.Y(net44)
);

FAx1_ASAP7_75t_R c70(
.A(net17),
.B(net43),
.CI(net33),
.SN(net46),
.CON(net45)
);

INVx11_ASAP7_75t_R c71(
.A(net28),
.Y(net47)
);

NOR2x1_ASAP7_75t_R c72(
.A(in3),
.B(net44),
.Y(net48)
);

MAJIxp5_ASAP7_75t_R c73(
.A(net33),
.B(in18),
.C(net47),
.Y(net49)
);

NOR2x1p5_ASAP7_75t_R c74(
.A(net41),
.B(net43),
.Y(net50)
);

NOR2x2_ASAP7_75t_R c75(
.A(net46),
.B(in20),
.Y(net51)
);

MAJx2_ASAP7_75t_R c76(
.A(net39),
.B(net21),
.C(net4),
.Y(net52)
);

MAJx3_ASAP7_75t_R c77(
.A(net16),
.B(net39),
.C(net12),
.Y(net53)
);

NAND3x1_ASAP7_75t_R c78(
.A(net4),
.B(net10),
.C(net11),
.Y(net54)
);

NAND3x2_ASAP7_75t_R c79(
.B(net11),
.C(net31),
.A(net51),
.Y(net55)
);

NAND3xp33_ASAP7_75t_R c80(
.A(net29),
.B(net55),
.C(net40),
.Y(net56)
);

NOR3x1_ASAP7_75t_R c81(
.A(net56),
.B(net45),
.C(in16),
.Y(net57)
);

NOR3x2_ASAP7_75t_R c82(
.B(net26),
.C(net56),
.A(net40),
.Y(net58)
);

NOR2xp33_ASAP7_75t_R c83(
.A(net44),
.B(net31),
.Y(net59)
);

INVx13_ASAP7_75t_R c84(
.A(net9171),
.Y(net60)
);

INVx1_ASAP7_75t_R c85(
.A(net31),
.Y(net61)
);

NOR3xp33_ASAP7_75t_R c86(
.A(net25),
.B(net107),
.C(in13),
.Y(net62)
);

INVx2_ASAP7_75t_R c87(
.A(net49),
.Y(net63)
);

NOR2xp67_ASAP7_75t_R c88(
.A(net51),
.B(net106),
.Y(net64)
);

INVx3_ASAP7_75t_R c89(
.A(net9650),
.Y(net65)
);

INVx4_ASAP7_75t_R c90(
.A(in14),
.Y(net66)
);

INVx5_ASAP7_75t_R c91(
.A(net41),
.Y(net67)
);

INVx6_ASAP7_75t_R c92(
.A(in13),
.Y(net68)
);

INVx8_ASAP7_75t_R c93(
.A(net37),
.Y(net69)
);

INVxp33_ASAP7_75t_R c94(
.A(net44),
.Y(net70)
);

INVxp67_ASAP7_75t_R c95(
.A(net9171),
.Y(net71)
);

ICGx1_ASAP7_75t_R c96(
.ENA(net60),
.SE(net107),
.CLK(clk),
.GCLK(net72)
);

BUFx10_ASAP7_75t_R c97(
.A(net106),
.Y(net73)
);

BUFx12_ASAP7_75t_R c98(
.A(net37),
.Y(net74)
);

BUFx12f_ASAP7_75t_R c99(
.A(net105),
.Y(net75)
);

BUFx16f_ASAP7_75t_R c100(
.A(net73),
.Y(net76)
);

OR2x2_ASAP7_75t_R c101(
.A(in8),
.B(net25),
.Y(net77)
);

OR2x4_ASAP7_75t_R c102(
.A(net25),
.B(net41),
.Y(net78)
);

OR2x6_ASAP7_75t_R c103(
.A(net71),
.B(net75),
.Y(net79)
);

BUFx24_ASAP7_75t_R c104(
.A(net66),
.Y(net80)
);

BUFx2_ASAP7_75t_R c105(
.A(net64),
.Y(net81)
);

XNOR2x1_ASAP7_75t_R c106(
.B(net74),
.A(net75),
.Y(net82)
);

BUFx3_ASAP7_75t_R c107(
.A(net72),
.Y(net83)
);

BUFx4_ASAP7_75t_R c108(
.A(net67),
.Y(net84)
);

XNOR2x2_ASAP7_75t_R c109(
.A(net82),
.B(net70),
.Y(net85)
);

BUFx4f_ASAP7_75t_R c110(
.A(net63),
.Y(net86)
);

BUFx5_ASAP7_75t_R c111(
.A(net77),
.Y(net87)
);

XNOR2xp5_ASAP7_75t_R c112(
.A(net74),
.B(net84),
.Y(net88)
);

BUFx6f_ASAP7_75t_R c113(
.A(net57),
.Y(net89)
);

BUFx8_ASAP7_75t_R c114(
.A(in10),
.Y(net90)
);

CKINVDCx10_ASAP7_75t_R c115(
.A(net90),
.Y(net91)
);

CKINVDCx11_ASAP7_75t_R c116(
.A(net66),
.Y(net92)
);

XOR2x1_ASAP7_75t_R c117(
.A(net86),
.B(net105),
.Y(net93)
);

CKINVDCx12_ASAP7_75t_R c118(
.A(net73),
.Y(net94)
);

CKINVDCx14_ASAP7_75t_R c119(
.A(net85),
.Y(net95)
);

CKINVDCx16_ASAP7_75t_R c120(
.A(net88),
.Y(net96)
);

XOR2x2_ASAP7_75t_R c121(
.A(net63),
.B(net41),
.Y(net97)
);

CKINVDCx20_ASAP7_75t_R c122(
.A(net65),
.Y(net98)
);

CKINVDCx5p33_ASAP7_75t_R c123(
.A(net92),
.Y(net99)
);

ICGx2_ASAP7_75t_R c124(
.ENA(net83),
.SE(net38),
.CLK(clk),
.GCLK(net100)
);

XOR2xp5_ASAP7_75t_R c125(
.A(net23),
.B(net100),
.Y(net101)
);

CKINVDCx6p67_ASAP7_75t_R c126(
.A(in1),
.Y(net102)
);

AND2x2_ASAP7_75t_R c127(
.A(net71),
.B(net57),
.Y(net103)
);

DFFASRHQNx1_ASAP7_75t_R c128(
.D(net98),
.RESETN(net103),
.SETN(net92),
.CLK(clk),
.QN(net104)
);

CKINVDCx8_ASAP7_75t_R c129(
.A(net13),
.Y(net105)
);

CKINVDCx9p33_ASAP7_75t_R c130(
.A(in14),
.Y(net106)
);

HB1xp67_ASAP7_75t_R c131(
.A(net57),
.Y(net107)
);

HB2xp67_ASAP7_75t_R c132(
.A(in18),
.Y(net108)
);

HB3xp67_ASAP7_75t_R c133(
.A(net81),
.Y(net109)
);

ICGx2p67DC_ASAP7_75t_R c134(
.ENA(net84),
.SE(net86),
.CLK(clk),
.GCLK(net110)
);

HB4xp67_ASAP7_75t_R c135(
.A(net50),
.Y(net111)
);

INVx11_ASAP7_75t_R c136(
.A(net95),
.Y(net112)
);

INVx13_ASAP7_75t_R c137(
.A(net112),
.Y(net113)
);

ICGx3_ASAP7_75t_R c138(
.ENA(net86),
.SE(net89),
.CLK(clk),
.GCLK(net114)
);

AND2x4_ASAP7_75t_R c139(
.A(net85),
.B(net92),
.Y(net115)
);

OA21x2_ASAP7_75t_R c140(
.A1(net112),
.A2(net99),
.B(net84),
.Y(net116)
);

ICGx4DC_ASAP7_75t_R c141(
.ENA(net116),
.SE(net92),
.CLK(clk),
.GCLK(net117)
);

ICGx4_ASAP7_75t_R c142(
.ENA(net113),
.SE(net110),
.CLK(clk),
.GCLK(net118)
);

AND2x6_ASAP7_75t_R c143(
.A(net91),
.B(net95),
.Y(net119)
);

HAxp5_ASAP7_75t_R c144(
.A(net67),
.B(net109),
.CON(net121),
.SN(net120)
);

NAND2x1_ASAP7_75t_R c145(
.A(net118),
.B(net9650),
.Y(net122)
);

NAND2x1p5_ASAP7_75t_R c146(
.A(net106),
.B(net65),
.Y(net123)
);

SDFHx1_ASAP7_75t_R c147(
.D(net103),
.SE(net57),
.SI(net76),
.CLK(clk),
.QN(net124)
);

ICGx5_ASAP7_75t_R c148(
.ENA(net76),
.SE(net38),
.CLK(clk),
.GCLK(net125)
);

ICGx5p33DC_ASAP7_75t_R c149(
.ENA(net89),
.SE(net122),
.CLK(clk),
.GCLK(net126)
);

NAND2x2_ASAP7_75t_R c150(
.A(net125),
.B(net60),
.Y(net127)
);

NAND2xp33_ASAP7_75t_R c151(
.A(net123),
.B(net102),
.Y(net128)
);

ICGx6p67DC_ASAP7_75t_R c152(
.ENA(net82),
.SE(net116),
.CLK(clk),
.GCLK(net129)
);

NAND2xp5_ASAP7_75t_R c153(
.A(in18),
.B(net119),
.Y(net130)
);

OAI21x1_ASAP7_75t_R c154(
.A1(net128),
.A2(net117),
.B(net123),
.Y(net131)
);

NAND2xp67_ASAP7_75t_R c155(
.A(net99),
.B(net94),
.Y(net132)
);

OAI21xp33_ASAP7_75t_R c156(
.A1(net81),
.A2(net127),
.B(net131),
.Y(net133)
);

ICGx8DC_ASAP7_75t_R c157(
.ENA(net121),
.SE(net125),
.CLK(clk),
.GCLK(net134)
);

OAI21xp5_ASAP7_75t_R c158(
.A1(net110),
.A2(net124),
.B(net134),
.Y(net135)
);

A2O1A1O1Ixp25_ASAP7_75t_R c159(
.A1(net131),
.A2(net133),
.B(net132),
.C(net119),
.D(net89),
.Y(net136)
);

OR3x1_ASAP7_75t_R c160(
.A(net134),
.B(net126),
.C(net135),
.Y(net137)
);

OR3x2_ASAP7_75t_R c161(
.A(net90),
.B(net128),
.C(net119),
.Y(net138)
);

AND5x1_ASAP7_75t_R c162(
.A(net127),
.B(net83),
.C(net120),
.D(net123),
.E(net119),
.Y(net139)
);

OR3x4_ASAP7_75t_R c163(
.A(net124),
.B(net5),
.C(net74),
.Y(net140)
);

AND3x1_ASAP7_75t_R c164(
.A(net132),
.B(net104),
.C(net134),
.Y(net141)
);

AND5x2_ASAP7_75t_R c165(
.A(net104),
.B(net140),
.C(net137),
.D(net129),
.E(net119),
.Y(net142)
);

INVx1_ASAP7_75t_R c166(
.A(net78),
.Y(net143)
);

INVx2_ASAP7_75t_R c167(
.A(net50),
.Y(net144)
);

NOR2x1_ASAP7_75t_R c168(
.A(net144),
.B(net96),
.Y(net145)
);

INVx3_ASAP7_75t_R c169(
.A(net9143),
.Y(net146)
);

INVx4_ASAP7_75t_R c170(
.A(in4),
.Y(net147)
);

INVx5_ASAP7_75t_R c171(
.A(net10173),
.Y(net148)
);

INVx6_ASAP7_75t_R c172(
.A(net35),
.Y(net149)
);

INVx8_ASAP7_75t_R c173(
.A(net145),
.Y(net150)
);

NOR2x1p5_ASAP7_75t_R c174(
.A(net147),
.B(net55),
.Y(net151)
);

INVxp33_ASAP7_75t_R c175(
.A(net10174),
.Y(net152)
);

INVxp67_ASAP7_75t_R c176(
.A(net61),
.Y(net153)
);

BUFx10_ASAP7_75t_R c177(
.A(net114),
.Y(net154)
);

BUFx12_ASAP7_75t_R c178(
.A(net150),
.Y(net155)
);

BUFx12f_ASAP7_75t_R c179(
.A(net80),
.Y(net156)
);

BUFx16f_ASAP7_75t_R c180(
.A(net119),
.Y(net157)
);

BUFx24_ASAP7_75t_R c181(
.A(net10173),
.Y(net158)
);

BUFx2_ASAP7_75t_R c182(
.A(net9143),
.Y(net159)
);

BUFx3_ASAP7_75t_R c183(
.A(net158),
.Y(net160)
);

NOR2x2_ASAP7_75t_R c184(
.A(net118),
.B(net114),
.Y(net161)
);

AND3x2_ASAP7_75t_R c185(
.A(net118),
.B(net114),
.C(net87),
.Y(net162)
);

BUFx4_ASAP7_75t_R c186(
.A(net141),
.Y(net163)
);

BUFx4f_ASAP7_75t_R c187(
.A(net55),
.Y(net164)
);

NOR2xp33_ASAP7_75t_R c188(
.A(net161),
.B(net129),
.Y(net165)
);

BUFx5_ASAP7_75t_R c189(
.A(net143),
.Y(net166)
);

BUFx6f_ASAP7_75t_R c190(
.A(net159),
.Y(net167)
);

BUFx8_ASAP7_75t_R c191(
.A(net101),
.Y(net168)
);

NOR2xp67_ASAP7_75t_R c192(
.A(net140),
.B(net165),
.Y(net169)
);

CKINVDCx10_ASAP7_75t_R c193(
.A(net167),
.Y(net170)
);

CKINVDCx11_ASAP7_75t_R c194(
.A(net166),
.Y(net171)
);

CKINVDCx12_ASAP7_75t_R c195(
.A(net9232),
.Y(net172)
);

CKINVDCx14_ASAP7_75t_R c196(
.A(net170),
.Y(net173)
);

OR2x2_ASAP7_75t_R c197(
.A(net164),
.B(net55),
.Y(net174)
);

OR2x4_ASAP7_75t_R c198(
.A(net164),
.B(net152),
.Y(net175)
);

CKINVDCx16_ASAP7_75t_R c199(
.A(in4),
.Y(net176)
);

CKINVDCx20_ASAP7_75t_R c200(
.A(net114),
.Y(net177)
);

CKINVDCx5p33_ASAP7_75t_R c201(
.A(net173),
.Y(net178)
);

CKINVDCx6p67_ASAP7_75t_R c202(
.A(in21),
.Y(net179)
);

OR2x6_ASAP7_75t_R c203(
.A(net78),
.B(net162),
.Y(net180)
);

AND3x4_ASAP7_75t_R c204(
.A(net175),
.B(net144),
.C(net101),
.Y(net181)
);

CKINVDCx8_ASAP7_75t_R c205(
.A(net158),
.Y(net182)
);

AO21x1_ASAP7_75t_R c206(
.A1(net50),
.A2(net172),
.B(net10174),
.Y(net183)
);

XNOR2x1_ASAP7_75t_R c207(
.B(net179),
.A(net154),
.Y(net184)
);

XNOR2x2_ASAP7_75t_R c208(
.A(net172),
.B(net123),
.Y(net185)
);

XNOR2xp5_ASAP7_75t_R c209(
.A(net162),
.B(net87),
.Y(net186)
);

CKINVDCx9p33_ASAP7_75t_R c210(
.A(net55),
.Y(net187)
);

HB1xp67_ASAP7_75t_R c211(
.A(net9889),
.Y(net188)
);

HB2xp67_ASAP7_75t_R c212(
.A(net169),
.Y(net189)
);

XOR2x1_ASAP7_75t_R c213(
.A(net186),
.B(net153),
.Y(net190)
);

XOR2x2_ASAP7_75t_R c214(
.A(net176),
.B(net167),
.Y(net191)
);

XOR2xp5_ASAP7_75t_R c215(
.A(net141),
.B(net146),
.Y(net192)
);

HB3xp67_ASAP7_75t_R c216(
.A(net190),
.Y(net193)
);

HB4xp67_ASAP7_75t_R c217(
.A(net190),
.Y(net194)
);

AO21x2_ASAP7_75t_R c218(
.A1(net189),
.A2(net169),
.B(net179),
.Y(net195)
);

AND2x2_ASAP7_75t_R c219(
.A(net182),
.B(net164),
.Y(net196)
);

AND2x4_ASAP7_75t_R c220(
.A(net196),
.B(net119),
.Y(net197)
);

INVx11_ASAP7_75t_R c221(
.A(net150),
.Y(net198)
);

INVx13_ASAP7_75t_R c222(
.A(net9864),
.Y(net199)
);

AOI21x1_ASAP7_75t_R c223(
.A1(net194),
.A2(net167),
.B(net180),
.Y(net200)
);

INVx1_ASAP7_75t_R c224(
.A(net101),
.Y(net201)
);

ICGx1_ASAP7_75t_R c225(
.ENA(net166),
.SE(net197),
.CLK(clk),
.GCLK(net202)
);

AND2x6_ASAP7_75t_R c226(
.A(net200),
.B(net164),
.Y(net203)
);

HAxp5_ASAP7_75t_R c227(
.A(net153),
.B(net202),
.CON(net204)
);

AOI21xp33_ASAP7_75t_R c228(
.A1(net80),
.A2(net192),
.B(net197),
.Y(net205)
);

INVx2_ASAP7_75t_R c229(
.A(net195),
.Y(net206)
);

AOI21xp5_ASAP7_75t_R c230(
.A1(net171),
.A2(net118),
.B(net9712),
.Y(net207)
);

NAND2x1_ASAP7_75t_R c231(
.A(net174),
.B(net169),
.Y(net208)
);

FAx1_ASAP7_75t_R c232(
.A(net94),
.B(net111),
.CI(net161),
.SN(net210),
.CON(net209)
);

MAJIxp5_ASAP7_75t_R c233(
.A(net198),
.B(net186),
.C(net10173),
.Y(net211)
);

NAND2x1p5_ASAP7_75t_R c234(
.A(net199),
.B(net171),
.Y(net212)
);

NAND2x2_ASAP7_75t_R c235(
.A(net177),
.B(net9712),
.Y(net213)
);

INVx3_ASAP7_75t_R c236(
.A(net165),
.Y(net214)
);

INVx4_ASAP7_75t_R c237(
.A(net201),
.Y(net215)
);

NAND2xp33_ASAP7_75t_R c238(
.A(net204),
.B(net151),
.Y(net216)
);

AO222x2_ASAP7_75t_R c239(
.A1(net160),
.A2(net216),
.B1(net207),
.B2(net89),
.C1(net180),
.C2(net146),
.Y(net217)
);

SDFHx2_ASAP7_75t_R c240(
.D(net207),
.SE(net193),
.SI(net198),
.CLK(clk),
.QN(net218)
);

NAND2xp5_ASAP7_75t_R c241(
.A(net189),
.B(net10175),
.Y(net219)
);

MAJx2_ASAP7_75t_R c242(
.A(net196),
.B(net207),
.C(net10175),
.Y(net220)
);

MAJx3_ASAP7_75t_R c243(
.A(net195),
.B(net9712),
.C(net10175),
.Y(net221)
);

INVx5_ASAP7_75t_R c244(
.A(net10550),
.Y(net222)
);

NAND3x1_ASAP7_75t_R c245(
.A(net222),
.B(net200),
.C(net9712),
.Y(net223)
);

SDFHx3_ASAP7_75t_R c246(
.D(net222),
.SE(net221),
.SI(net10175),
.CLK(clk),
.QN(net224)
);

NAND3x2_ASAP7_75t_R c247(
.B(net149),
.C(net221),
.A(net10175),
.Y(net225)
);

NAND3xp33_ASAP7_75t_R c248(
.A(net163),
.B(net222),
.C(net177),
.Y(net226)
);

INVx6_ASAP7_75t_R c249(
.A(net148),
.Y(net227)
);

INVx8_ASAP7_75t_R c250(
.A(net69),
.Y(net228)
);

INVxp33_ASAP7_75t_R c251(
.A(net238),
.Y(net229)
);

INVxp67_ASAP7_75t_R c252(
.A(net173),
.Y(net230)
);

BUFx10_ASAP7_75t_R c253(
.A(net226),
.Y(net231)
);

BUFx12_ASAP7_75t_R c254(
.A(net98),
.Y(net232)
);

NAND2xp67_ASAP7_75t_R c255(
.A(net227),
.B(net161),
.Y(net233)
);

BUFx12f_ASAP7_75t_R c256(
.A(net10088),
.Y(net234)
);

BUFx16f_ASAP7_75t_R c257(
.A(net9121),
.Y(net235)
);

BUFx24_ASAP7_75t_R c258(
.A(net17),
.Y(net236)
);

BUFx2_ASAP7_75t_R c259(
.A(net75),
.Y(net237)
);

BUFx3_ASAP7_75t_R c260(
.A(net96),
.Y(net238)
);

BUFx4_ASAP7_75t_R c261(
.A(net183),
.Y(net239)
);

BUFx4f_ASAP7_75t_R c262(
.A(net26),
.Y(net240)
);

BUFx5_ASAP7_75t_R c263(
.A(net75),
.Y(net241)
);

BUFx6f_ASAP7_75t_R c264(
.A(net5),
.Y(net242)
);

BUFx8_ASAP7_75t_R c265(
.A(net213),
.Y(net243)
);

CKINVDCx10_ASAP7_75t_R c266(
.A(net236),
.Y(net244)
);

CKINVDCx11_ASAP7_75t_R c267(
.A(net234),
.Y(net245)
);

NOR2x1_ASAP7_75t_R c268(
.A(net168),
.B(net229),
.Y(net246)
);

NOR2x1p5_ASAP7_75t_R c269(
.A(net152),
.B(net183),
.Y(net247)
);

NOR2x2_ASAP7_75t_R c270(
.A(net96),
.B(net192),
.Y(net248)
);

CKINVDCx12_ASAP7_75t_R c271(
.A(net182),
.Y(net249)
);

CKINVDCx14_ASAP7_75t_R c272(
.A(net226),
.Y(net250)
);

CKINVDCx16_ASAP7_75t_R c273(
.A(net247),
.Y(net251)
);

NOR2xp33_ASAP7_75t_R c274(
.A(net251),
.B(net230),
.Y(net252)
);

CKINVDCx20_ASAP7_75t_R c275(
.A(net214),
.Y(net253)
);

CKINVDCx5p33_ASAP7_75t_R c276(
.A(net251),
.Y(net254)
);

CKINVDCx6p67_ASAP7_75t_R c277(
.A(net247),
.Y(net255)
);

CKINVDCx8_ASAP7_75t_R c278(
.A(net9121),
.Y(net256)
);

NOR3x1_ASAP7_75t_R c279(
.A(net248),
.B(net243),
.C(net256),
.Y(net257)
);

NOR3x2_ASAP7_75t_R c280(
.B(net252),
.C(net228),
.A(net255),
.Y(net258)
);

NOR2xp67_ASAP7_75t_R c281(
.A(net249),
.B(net214),
.Y(net259)
);

CKINVDCx9p33_ASAP7_75t_R c282(
.A(net238),
.Y(net260)
);

NOR3xp33_ASAP7_75t_R c283(
.A(net257),
.B(net231),
.C(net219),
.Y(net261)
);

OR2x2_ASAP7_75t_R c284(
.A(net260),
.B(net237),
.Y(net262)
);

OR2x4_ASAP7_75t_R c285(
.A(net192),
.B(net161),
.Y(net263)
);

OR2x6_ASAP7_75t_R c286(
.A(net239),
.B(net168),
.Y(net264)
);

HB1xp67_ASAP7_75t_R c287(
.A(net232),
.Y(net265)
);

HB2xp67_ASAP7_75t_R c288(
.A(net230),
.Y(net266)
);

HB3xp67_ASAP7_75t_R c289(
.A(net10415),
.Y(net267)
);

HB4xp67_ASAP7_75t_R c290(
.A(net10031),
.Y(net268)
);

INVx11_ASAP7_75t_R c291(
.A(net9828),
.Y(net269)
);

INVx13_ASAP7_75t_R c292(
.A(net9934),
.Y(net270)
);

OA21x2_ASAP7_75t_R c293(
.A1(net243),
.A2(net259),
.B(net174),
.Y(net271)
);

XNOR2x1_ASAP7_75t_R c294(
.B(net250),
.A(net137),
.Y(net272)
);

INVx1_ASAP7_75t_R c295(
.A(net161),
.Y(net273)
);

SDFHx4_ASAP7_75t_R c296(
.D(net269),
.SE(net264),
.SI(net271),
.CLK(clk),
.QN(net274)
);

AO221x1_ASAP7_75t_R c297(
.A1(net266),
.A2(net213),
.B1(net173),
.B2(net245),
.C(net270),
.Y(net275)
);

INVx2_ASAP7_75t_R c298(
.A(net273),
.Y(net276)
);

INVx3_ASAP7_75t_R c299(
.A(net275),
.Y(net277)
);

OAI21x1_ASAP7_75t_R c300(
.A1(net148),
.A2(net258),
.B(net234),
.Y(net278)
);

XNOR2x2_ASAP7_75t_R c301(
.A(net265),
.B(net229),
.Y(net279)
);

SDFLx1_ASAP7_75t_R c302(
.D(net229),
.SE(net279),
.SI(net266),
.CLK(clk),
.QN(net280)
);

XNOR2xp5_ASAP7_75t_R c303(
.A(net254),
.B(net264),
.Y(net281)
);

XOR2x1_ASAP7_75t_R c304(
.A(net235),
.B(net274),
.Y(net282)
);

INVx4_ASAP7_75t_R c305(
.A(net267),
.Y(net283)
);

INVx5_ASAP7_75t_R c306(
.A(net10507),
.Y(net284)
);

XOR2x2_ASAP7_75t_R c307(
.A(net280),
.B(net146),
.Y(net285)
);

OAI21xp33_ASAP7_75t_R c308(
.A1(net237),
.A2(net283),
.B(net256),
.Y(net286)
);

OAI21xp5_ASAP7_75t_R c309(
.A1(net286),
.A2(net285),
.B(net266),
.Y(net287)
);

XOR2xp5_ASAP7_75t_R c310(
.A(net233),
.B(net214),
.Y(net288)
);

OR3x1_ASAP7_75t_R c311(
.A(net213),
.B(net262),
.C(net69),
.Y(net289)
);

INVx6_ASAP7_75t_R c312(
.A(net10013),
.Y(net290)
);

OR3x2_ASAP7_75t_R c313(
.A(net256),
.B(net283),
.C(net10108),
.Y(net291)
);

AND2x2_ASAP7_75t_R c314(
.A(net291),
.B(net264),
.Y(net292)
);

OR3x4_ASAP7_75t_R c315(
.A(net285),
.B(net270),
.C(net9953),
.Y(net293)
);

AND2x4_ASAP7_75t_R c316(
.A(net231),
.B(net252),
.Y(net294)
);

INVx8_ASAP7_75t_R c317(
.A(net9926),
.Y(net295)
);

AND3x1_ASAP7_75t_R c318(
.A(net285),
.B(net295),
.C(net245),
.Y(net296)
);

SDFLx2_ASAP7_75t_R c319(
.D(net294),
.SE(net284),
.SI(net174),
.CLK(clk),
.QN(net297)
);

INVxp33_ASAP7_75t_R c320(
.A(net283),
.Y(net298)
);

AND2x6_ASAP7_75t_R c321(
.A(net298),
.B(net251),
.Y(net299)
);

AND3x2_ASAP7_75t_R c322(
.A(net282),
.B(net292),
.C(net250),
.Y(net300)
);

A2O1A1Ixp33_ASAP7_75t_R c323(
.A1(net234),
.A2(net283),
.B(net300),
.C(net271),
.Y(net301)
);

AO33x2_ASAP7_75t_R c324(
.A1(net296),
.A2(net300),
.A3(net259),
.B1(net245),
.B2(net10108),
.B3(net10176),
.Y(net302)
);

SDFLx3_ASAP7_75t_R c325(
.D(net219),
.SE(net271),
.SI(net9953),
.CLK(clk),
.QN(net303)
);

SDFLx4_ASAP7_75t_R c326(
.D(net258),
.SE(net285),
.SI(net291),
.CLK(clk),
.QN(net304)
);

INVxp67_ASAP7_75t_R c327(
.A(net9950),
.Y(net305)
);

HAxp5_ASAP7_75t_R c328(
.A(net292),
.B(net295),
.CON(net307),
.SN(net306)
);

AND3x4_ASAP7_75t_R c329(
.A(net307),
.B(net300),
.Y(net308)
);

AO221x2_ASAP7_75t_R c330(
.A1(net277),
.A2(net282),
.B1(net186),
.B2(net306),
.C(net9648),
.Y(net309)
);

AO32x1_ASAP7_75t_R c331(
.A1(net305),
.A2(net182),
.A3(net161),
.B1(net9648),
.B2(net10177),
.Y(net310)
);

BUFx10_ASAP7_75t_R c332(
.A(net295),
.Y(net311)
);

NAND2x1_ASAP7_75t_R c333(
.A(net129),
.B(net276),
.Y(net312)
);

BUFx12_ASAP7_75t_R c334(
.A(net154),
.Y(net313)
);

BUFx12f_ASAP7_75t_R c335(
.A(net154),
.Y(net314)
);

NAND2x1p5_ASAP7_75t_R c336(
.A(net224),
.B(net146),
.Y(net315)
);

NAND2x2_ASAP7_75t_R c337(
.A(net129),
.B(net275),
.Y(net316)
);

BUFx16f_ASAP7_75t_R c338(
.A(net180),
.Y(net317)
);

BUFx24_ASAP7_75t_R c339(
.A(net123),
.Y(net318)
);

BUFx2_ASAP7_75t_R c340(
.A(net10047),
.Y(net319)
);

BUFx3_ASAP7_75t_R c341(
.A(net10130),
.Y(net320)
);

BUFx4_ASAP7_75t_R c342(
.A(net290),
.Y(net321)
);

BUFx4f_ASAP7_75t_R c343(
.A(net275),
.Y(net322)
);

BUFx5_ASAP7_75t_R c344(
.A(net257),
.Y(net323)
);

BUFx6f_ASAP7_75t_R c345(
.A(net310),
.Y(net324)
);

BUFx8_ASAP7_75t_R c346(
.A(net274),
.Y(net325)
);

CKINVDCx10_ASAP7_75t_R c347(
.A(net10542),
.Y(net326)
);

CKINVDCx11_ASAP7_75t_R c348(
.A(net304),
.Y(net327)
);

CKINVDCx12_ASAP7_75t_R c349(
.A(net303),
.Y(net328)
);

CKINVDCx14_ASAP7_75t_R c350(
.A(net321),
.Y(net329)
);

CKINVDCx16_ASAP7_75t_R c351(
.A(net256),
.Y(net330)
);

CKINVDCx20_ASAP7_75t_R c352(
.A(net259),
.Y(net331)
);

NAND2xp33_ASAP7_75t_R c353(
.A(net274),
.B(net268),
.Y(net332)
);

CKINVDCx5p33_ASAP7_75t_R c354(
.A(net320),
.Y(net333)
);

NAND2xp5_ASAP7_75t_R c355(
.A(net333),
.B(net326),
.Y(net334)
);

CKINVDCx6p67_ASAP7_75t_R c356(
.A(net216),
.Y(net335)
);

CKINVDCx8_ASAP7_75t_R c357(
.A(net188),
.Y(net336)
);

CKINVDCx9p33_ASAP7_75t_R c358(
.A(in11),
.Y(net337)
);

NAND2xp67_ASAP7_75t_R c359(
.A(net337),
.B(net146),
.Y(net338)
);

NOR2x1_ASAP7_75t_R c360(
.A(net332),
.B(in11),
.Y(net339)
);

HB1xp67_ASAP7_75t_R c361(
.A(net334),
.Y(net340)
);

NOR2x1p5_ASAP7_75t_R c362(
.A(net303),
.B(net174),
.Y(net341)
);

NOR2x2_ASAP7_75t_R c363(
.A(net337),
.B(net325),
.Y(net342)
);

HB2xp67_ASAP7_75t_R c364(
.A(net10130),
.Y(net343)
);

NOR2xp33_ASAP7_75t_R c365(
.A(net227),
.B(net336),
.Y(net344)
);

NOR2xp67_ASAP7_75t_R c366(
.A(net329),
.B(net314),
.Y(net345)
);

HB3xp67_ASAP7_75t_R c367(
.A(net344),
.Y(net346)
);

HB4xp67_ASAP7_75t_R c368(
.A(net9239),
.Y(net347)
);

OR2x2_ASAP7_75t_R c369(
.A(net343),
.B(net316),
.Y(net348)
);

OR2x4_ASAP7_75t_R c370(
.A(net345),
.B(net259),
.Y(net349)
);

INVx11_ASAP7_75t_R c371(
.A(net320),
.Y(net350)
);

OR2x6_ASAP7_75t_R c372(
.A(net212),
.B(net339),
.Y(net351)
);

INVx13_ASAP7_75t_R c373(
.A(net268),
.Y(net352)
);

AO21x1_ASAP7_75t_R c374(
.A1(net317),
.A2(net290),
.B(net311),
.Y(net353)
);

INVx1_ASAP7_75t_R c375(
.A(net316),
.Y(net354)
);

XNOR2x1_ASAP7_75t_R c376(
.B(net328),
.A(net347),
.Y(net355)
);

XNOR2x2_ASAP7_75t_R c377(
.A(net340),
.B(net344),
.Y(net356)
);

XNOR2xp5_ASAP7_75t_R c378(
.A(net347),
.B(net344),
.Y(net357)
);

INVx2_ASAP7_75t_R c379(
.A(net9907),
.Y(net358)
);

INVx3_ASAP7_75t_R c380(
.A(net313),
.Y(net359)
);

XOR2x1_ASAP7_75t_R c381(
.A(net350),
.B(net313),
.Y(net360)
);

XOR2x2_ASAP7_75t_R c382(
.A(net346),
.B(net343),
.Y(net361)
);

XOR2xp5_ASAP7_75t_R c383(
.A(net360),
.B(net354),
.Y(net362)
);

INVx4_ASAP7_75t_R c384(
.A(net344),
.Y(net363)
);

INVx5_ASAP7_75t_R c385(
.A(net361),
.Y(net364)
);

AND2x2_ASAP7_75t_R c386(
.A(net314),
.B(net358),
.Y(net365)
);

AO21x2_ASAP7_75t_R c387(
.A1(net362),
.A2(net268),
.B(net332),
.Y(net366)
);

AND2x4_ASAP7_75t_R c388(
.A(net349),
.B(net304),
.Y(net367)
);

INVx6_ASAP7_75t_R c389(
.A(net322),
.Y(net368)
);

INVx8_ASAP7_75t_R c390(
.A(net334),
.Y(net369)
);

AND2x6_ASAP7_75t_R c391(
.A(net324),
.B(net312),
.Y(net370)
);

HAxp5_ASAP7_75t_R c392(
.A(net368),
.B(net331),
.CON(net372),
.SN(net371)
);

NAND2x1_ASAP7_75t_R c393(
.A(net336),
.B(net371),
.Y(net373)
);

NAND2x1p5_ASAP7_75t_R c394(
.A(net364),
.B(net339),
.Y(net374)
);

AOI21x1_ASAP7_75t_R c395(
.A1(net321),
.A2(net367),
.B(net180),
.Y(net375)
);

AOI21xp33_ASAP7_75t_R c396(
.A1(net360),
.A2(net369),
.B(net327),
.Y(net376)
);

NAND2x2_ASAP7_75t_R c397(
.A(net366),
.B(net352),
.Y(net377)
);

NAND2xp33_ASAP7_75t_R c398(
.A(net373),
.B(net319),
.Y(net378)
);

NAND2xp5_ASAP7_75t_R c399(
.A(net352),
.B(net376),
.Y(net379)
);

NAND2xp67_ASAP7_75t_R c400(
.A(net348),
.B(net9681),
.Y(net380)
);

AOI21xp5_ASAP7_75t_R c401(
.A1(net354),
.A2(net346),
.B(net9681),
.Y(net381)
);

DFFASRHQNx1_ASAP7_75t_R c402(
.D(net335),
.RESETN(net365),
.SETN(net345),
.CLK(clk),
.QN(net382)
);

FAx1_ASAP7_75t_R c403(
.A(net363),
.B(net370),
.CI(net374),
.SN(net383)
);

NOR2x1_ASAP7_75t_R c404(
.A(net362),
.B(net9681),
.Y(net384)
);

NOR2x1p5_ASAP7_75t_R c405(
.A(net383),
.B(net332),
.Y(net385)
);

NOR2x2_ASAP7_75t_R c406(
.A(net376),
.B(net384),
.Y(net386)
);

MAJIxp5_ASAP7_75t_R c407(
.A(net379),
.B(net314),
.C(net9681),
.Y(net387)
);

INVxp33_ASAP7_75t_R c408(
.A(net9954),
.Y(net388)
);

SDFHx1_ASAP7_75t_R c409(
.D(net369),
.SE(net384),
.SI(net388),
.CLK(clk),
.QN(net389)
);

AND4x1_ASAP7_75t_R c410(
.A(net388),
.B(net364),
.C(net389),
.D(net385),
.Y(net390)
);

AND4x2_ASAP7_75t_R c411(
.A(net357),
.B(net390),
.C(net380),
.D(net388),
.Y(net391)
);

AO211x2_ASAP7_75t_R c412(
.A1(net355),
.A2(net384),
.B(net385),
.C(net390),
.Y(net392)
);

MAJx2_ASAP7_75t_R c413(
.A(net370),
.B(net355),
.C(net9896),
.Y(net393)
);

AO22x1_ASAP7_75t_R c414(
.A1(net367),
.A2(net376),
.B1(net385),
.B2(net388),
.Y(net394)
);

INVxp67_ASAP7_75t_R c415(
.A(net293),
.Y(net395)
);

BUFx10_ASAP7_75t_R c416(
.A(net372),
.Y(net396)
);

BUFx12_ASAP7_75t_R c417(
.A(net395),
.Y(net397)
);

BUFx12f_ASAP7_75t_R c418(
.A(net9271),
.Y(net398)
);

NOR2xp33_ASAP7_75t_R c419(
.A(net361),
.B(net381),
.Y(net399)
);

MAJx3_ASAP7_75t_R c420(
.A(net385),
.B(net395),
.C(net330),
.Y(net400)
);

BUFx16f_ASAP7_75t_R c421(
.A(net397),
.Y(net401)
);

NOR2xp67_ASAP7_75t_R c422(
.A(net374),
.B(net10178),
.Y(net402)
);

BUFx24_ASAP7_75t_R c423(
.A(net401),
.Y(net403)
);

BUFx2_ASAP7_75t_R c424(
.A(net312),
.Y(net404)
);

OR2x2_ASAP7_75t_R c425(
.A(net137),
.B(net142),
.Y(net405)
);

BUFx3_ASAP7_75t_R c426(
.A(net312),
.Y(net406)
);

BUFx4_ASAP7_75t_R c427(
.A(net372),
.Y(net407)
);

OR2x4_ASAP7_75t_R c428(
.A(net406),
.B(net353),
.Y(net408)
);

AO22x2_ASAP7_75t_R c429(
.A1(net403),
.A2(net287),
.B1(net326),
.B2(net10178),
.Y(net409)
);

OR2x6_ASAP7_75t_R c430(
.A(net317),
.B(net10177),
.Y(net410)
);

BUFx4f_ASAP7_75t_R c431(
.A(net244),
.Y(net411)
);

XNOR2x1_ASAP7_75t_R c432(
.B(net393),
.A(net295),
.Y(net412)
);

BUFx5_ASAP7_75t_R c433(
.A(net411),
.Y(net413)
);

BUFx6f_ASAP7_75t_R c434(
.A(net287),
.Y(net414)
);

BUFx8_ASAP7_75t_R c435(
.A(net324),
.Y(net415)
);

CKINVDCx10_ASAP7_75t_R c436(
.A(net34),
.Y(net416)
);

CKINVDCx11_ASAP7_75t_R c437(
.A(net415),
.Y(net417)
);

CKINVDCx12_ASAP7_75t_R c438(
.A(net9090),
.Y(net418)
);

XNOR2x2_ASAP7_75t_R c439(
.A(net276),
.B(net412),
.Y(net419)
);

CKINVDCx14_ASAP7_75t_R c440(
.A(net359),
.Y(net420)
);

CKINVDCx16_ASAP7_75t_R c441(
.A(net248),
.Y(net421)
);

CKINVDCx20_ASAP7_75t_R c442(
.A(net187),
.Y(net422)
);

CKINVDCx5p33_ASAP7_75t_R c443(
.A(net418),
.Y(net423)
);

XNOR2xp5_ASAP7_75t_R c444(
.A(net157),
.B(net398),
.Y(net424)
);

XOR2x1_ASAP7_75t_R c445(
.A(net419),
.B(net415),
.Y(net425)
);

XOR2x2_ASAP7_75t_R c446(
.A(net412),
.B(net293),
.Y(net426)
);

NAND3x1_ASAP7_75t_R c447(
.A(net403),
.B(net418),
.C(net412),
.Y(net427)
);

XOR2xp5_ASAP7_75t_R c448(
.A(net416),
.B(net421),
.Y(net428)
);

CKINVDCx6p67_ASAP7_75t_R c449(
.A(net417),
.Y(net429)
);

AND2x2_ASAP7_75t_R c450(
.A(net387),
.B(net418),
.Y(net430)
);

NAND3x2_ASAP7_75t_R c451(
.B(net399),
.C(net414),
.A(net426),
.Y(net431)
);

CKINVDCx8_ASAP7_75t_R c452(
.A(net9090),
.Y(net432)
);

CKINVDCx9p33_ASAP7_75t_R c453(
.A(net9636),
.Y(net433)
);

HB1xp67_ASAP7_75t_R c454(
.A(net414),
.Y(net434)
);

HB2xp67_ASAP7_75t_R c455(
.A(net9636),
.Y(net435)
);

AND2x4_ASAP7_75t_R c456(
.A(net382),
.B(net421),
.Y(net436)
);

HB3xp67_ASAP7_75t_R c457(
.A(net416),
.Y(net437)
);

HB4xp67_ASAP7_75t_R c458(
.A(net10120),
.Y(net438)
);

INVx11_ASAP7_75t_R c459(
.A(net9269),
.Y(net439)
);

NAND3xp33_ASAP7_75t_R c460(
.A(net287),
.B(net433),
.C(net422),
.Y(net440)
);

INVx13_ASAP7_75t_R c461(
.A(net9269),
.Y(net441)
);

NOR3x1_ASAP7_75t_R c462(
.A(net310),
.B(net427),
.C(net429),
.Y(net442)
);

AND2x6_ASAP7_75t_R c463(
.A(net432),
.B(net293),
.Y(net443)
);

INVx1_ASAP7_75t_R c464(
.A(net442),
.Y(net444)
);

INVx2_ASAP7_75t_R c465(
.A(net10411),
.Y(net445)
);

NOR3x2_ASAP7_75t_R c466(
.B(net430),
.C(net331),
.A(net411),
.Y(net446)
);

HAxp5_ASAP7_75t_R c467(
.A(net415),
.B(net429),
.CON(net448),
.SN(net447)
);

NAND2x1_ASAP7_75t_R c468(
.A(net69),
.B(net409),
.Y(net449)
);

NAND2x1p5_ASAP7_75t_R c469(
.A(net399),
.B(net421),
.Y(net450)
);

NAND2x2_ASAP7_75t_R c470(
.A(net434),
.B(net439),
.Y(net451)
);

INVx3_ASAP7_75t_R c471(
.A(net438),
.Y(net452)
);

INVx4_ASAP7_75t_R c472(
.A(net430),
.Y(net453)
);

NAND2xp33_ASAP7_75t_R c473(
.A(net451),
.B(net248),
.Y(net454)
);

NOR3xp33_ASAP7_75t_R c474(
.A(net410),
.B(net434),
.C(net401),
.Y(net455)
);

OA21x2_ASAP7_75t_R c475(
.A1(net398),
.A2(net310),
.B(net435),
.Y(net456)
);

NAND2xp5_ASAP7_75t_R c476(
.A(net406),
.B(net387),
.Y(net457)
);

SDFHx2_ASAP7_75t_R c477(
.D(net437),
.SE(net417),
.SI(net382),
.CLK(clk),
.QN(net458)
);

INVx5_ASAP7_75t_R c478(
.A(net453),
.Y(net459)
);

OAI21x1_ASAP7_75t_R c479(
.A1(net459),
.A2(net451),
.B(net458),
.Y(net460)
);

OAI21xp33_ASAP7_75t_R c480(
.A1(net402),
.A2(net350),
.B(net9783),
.Y(net461)
);

NAND2xp67_ASAP7_75t_R c481(
.A(net425),
.B(net447),
.Y(net462)
);

INVx6_ASAP7_75t_R c482(
.A(net330),
.Y(net463)
);

INVx8_ASAP7_75t_R c483(
.A(net463),
.Y(net464)
);

INVxp33_ASAP7_75t_R c484(
.A(net9933),
.Y(net465)
);

NOR2x1_ASAP7_75t_R c485(
.A(net464),
.B(net10012),
.Y(net466)
);

OAI21xp5_ASAP7_75t_R c486(
.A1(net457),
.A2(net464),
.B(net9933),
.Y(net467)
);

OR3x1_ASAP7_75t_R c487(
.A(net408),
.B(net432),
.C(net459),
.Y(net468)
);

OR3x2_ASAP7_75t_R c488(
.A(net461),
.B(net406),
.C(net420),
.Y(net469)
);

OR3x4_ASAP7_75t_R c489(
.A(net433),
.B(net338),
.C(net425),
.Y(net470)
);

SDFHx3_ASAP7_75t_R c490(
.D(net456),
.SE(net426),
.SI(net437),
.CLK(clk),
.QN(net471)
);

AND3x1_ASAP7_75t_R c491(
.A(net471),
.B(net418),
.C(net10012),
.Y(net472)
);

AO32x2_ASAP7_75t_R c492(
.A1(net469),
.A2(net426),
.A3(net467),
.B1(net390),
.B2(net462),
.Y(net473)
);

NOR2x1p5_ASAP7_75t_R c493(
.A(net471),
.B(net432),
.Y(net474)
);

INVxp67_ASAP7_75t_R c494(
.A(net10481),
.Y(net475)
);

ICGx2_ASAP7_75t_R c495(
.ENA(net455),
.SE(net413),
.CLK(clk),
.GCLK(net476)
);

AND3x2_ASAP7_75t_R c496(
.A(net475),
.B(net474),
.C(net382),
.Y(net477)
);

AND3x4_ASAP7_75t_R c497(
.A(net477),
.B(net474),
.C(net467),
.Y(net478)
);

BUFx10_ASAP7_75t_R c498(
.A(net9172),
.Y(net479)
);

BUFx12_ASAP7_75t_R c499(
.A(net374),
.Y(net480)
);

NOR2x2_ASAP7_75t_R c500(
.A(net504),
.B(net10179),
.Y(net481)
);

NOR2xp33_ASAP7_75t_R c501(
.A(net59),
.B(net494),
.Y(net482)
);

BUFx12f_ASAP7_75t_R c502(
.A(net507),
.Y(net483)
);

BUFx16f_ASAP7_75t_R c503(
.A(net482),
.Y(net484)
);

NOR2xp67_ASAP7_75t_R c504(
.A(net496),
.B(net509),
.Y(net485)
);

BUFx24_ASAP7_75t_R c505(
.A(net326),
.Y(net486)
);

OR2x2_ASAP7_75t_R c506(
.A(net485),
.B(net478),
.Y(net487)
);

BUFx2_ASAP7_75t_R c507(
.A(net496),
.Y(net488)
);

OR2x4_ASAP7_75t_R c508(
.A(net505),
.B(net480),
.Y(net489)
);

OR2x6_ASAP7_75t_R c509(
.A(net489),
.B(net508),
.Y(net490)
);

BUFx3_ASAP7_75t_R c510(
.A(net9966),
.Y(net491)
);

BUFx4_ASAP7_75t_R c511(
.A(net146),
.Y(net492)
);

BUFx4f_ASAP7_75t_R c512(
.A(net494),
.Y(net493)
);

BUFx5_ASAP7_75t_R c513(
.A(net9172),
.Y(net494)
);

XNOR2x1_ASAP7_75t_R c514(
.B(net453),
.A(net245),
.Y(net495)
);

BUFx6f_ASAP7_75t_R c515(
.A(net146),
.Y(net496)
);

BUFx8_ASAP7_75t_R c516(
.A(net472),
.Y(net497)
);

CKINVDCx10_ASAP7_75t_R c517(
.A(net443),
.Y(net498)
);

CKINVDCx11_ASAP7_75t_R c518(
.A(net380),
.Y(net499)
);

CKINVDCx12_ASAP7_75t_R c519(
.A(net10177),
.Y(net500)
);

CKINVDCx14_ASAP7_75t_R c520(
.A(net495),
.Y(net501)
);

CKINVDCx16_ASAP7_75t_R c521(
.A(net446),
.Y(net502)
);

CKINVDCx20_ASAP7_75t_R c522(
.A(net380),
.Y(net503)
);

CKINVDCx5p33_ASAP7_75t_R c523(
.A(net10393),
.Y(net504)
);

XNOR2x2_ASAP7_75t_R c524(
.A(net432),
.B(net441),
.Y(net505)
);

CKINVDCx6p67_ASAP7_75t_R c525(
.A(net381),
.Y(net506)
);

CKINVDCx8_ASAP7_75t_R c526(
.A(net457),
.Y(net507)
);

CKINVDCx9p33_ASAP7_75t_R c527(
.A(net326),
.Y(net508)
);

ICGx2p67DC_ASAP7_75t_R c528(
.ENA(net341),
.SE(net501),
.CLK(clk),
.GCLK(net509)
);

HB1xp67_ASAP7_75t_R c529(
.A(net481),
.Y(net510)
);

SDFHx4_ASAP7_75t_R c530(
.D(net341),
.SE(net381),
.SI(net343),
.CLK(clk),
.QN(net511)
);

XNOR2xp5_ASAP7_75t_R c531(
.A(net507),
.B(net508),
.Y(net512)
);

XOR2x1_ASAP7_75t_R c532(
.A(net419),
.B(net34),
.Y(net513)
);

XOR2x2_ASAP7_75t_R c533(
.A(net508),
.B(net10111),
.Y(net514)
);

XOR2xp5_ASAP7_75t_R c534(
.A(net349),
.B(net498),
.Y(net515)
);

AND2x2_ASAP7_75t_R c535(
.A(net515),
.B(net493),
.Y(net516)
);

HB2xp67_ASAP7_75t_R c536(
.A(net511),
.Y(net517)
);

AO21x1_ASAP7_75t_R c537(
.A1(net492),
.A2(net339),
.B(net468),
.Y(net518)
);

AND2x4_ASAP7_75t_R c538(
.A(net514),
.B(net493),
.Y(net519)
);

HB3xp67_ASAP7_75t_R c539(
.A(net10564),
.Y(net520)
);

AO21x2_ASAP7_75t_R c540(
.A1(net470),
.A2(net423),
.B(net447),
.Y(net521)
);

AND2x6_ASAP7_75t_R c541(
.A(net480),
.B(net493),
.Y(net522)
);

HAxp5_ASAP7_75t_R c542(
.A(net374),
.B(net488),
.CON(net524),
.SN(net523)
);

NAND2x1_ASAP7_75t_R c543(
.A(net432),
.B(net9738),
.Y(net525)
);

NAND2x1p5_ASAP7_75t_R c544(
.A(net449),
.B(net511),
.Y(net526)
);

NAND2x2_ASAP7_75t_R c545(
.A(net520),
.B(net514),
.Y(net527)
);

NAND2xp33_ASAP7_75t_R c546(
.A(net465),
.B(net476),
.Y(net528)
);

HB4xp67_ASAP7_75t_R c547(
.A(net486),
.Y(net529)
);

NAND2xp5_ASAP7_75t_R c548(
.A(net523),
.B(net484),
.Y(net530)
);

NAND2xp67_ASAP7_75t_R c549(
.A(net9738),
.B(net10111),
.Y(net531)
);

NOR2x1_ASAP7_75t_R c550(
.A(net528),
.B(net520),
.Y(net532)
);

NOR2x1p5_ASAP7_75t_R c551(
.A(net493),
.B(net517),
.Y(net533)
);

NOR2x2_ASAP7_75t_R c552(
.A(net533),
.B(net530),
.Y(net534)
);

NOR2xp33_ASAP7_75t_R c553(
.A(net530),
.B(net528),
.Y(net535)
);

NOR2xp67_ASAP7_75t_R c554(
.A(net532),
.B(net512),
.Y(net536)
);

OR2x2_ASAP7_75t_R c555(
.A(net524),
.B(net531),
.Y(net537)
);

OR2x4_ASAP7_75t_R c556(
.A(net527),
.B(net412),
.Y(net538)
);

AOI221x1_ASAP7_75t_R c557(
.A1(net491),
.A2(net505),
.B1(net187),
.B2(net534),
.C(net445),
.Y(net539)
);

OR2x6_ASAP7_75t_R c558(
.A(net508),
.B(net496),
.Y(net540)
);

ICGx3_ASAP7_75t_R c559(
.ENA(net485),
.SE(net536),
.CLK(clk),
.GCLK(net541)
);

AOI222xp33_ASAP7_75t_R c560(
.A1(net504),
.A2(net514),
.B1(net492),
.B2(net496),
.C1(net534),
.C2(net541),
.Y(net542)
);

AOI21x1_ASAP7_75t_R c561(
.A1(net509),
.A2(net491),
.B(net445),
.Y(net543)
);

XNOR2x1_ASAP7_75t_R c562(
.B(net497),
.A(net533),
.Y(net544)
);

XNOR2x2_ASAP7_75t_R c563(
.A(net442),
.B(net526),
.Y(net545)
);

XNOR2xp5_ASAP7_75t_R c564(
.A(net481),
.B(net530),
.Y(net546)
);

INVx11_ASAP7_75t_R c565(
.A(net9966),
.Y(net547)
);

AOI21xp33_ASAP7_75t_R c566(
.A1(net544),
.A2(net532),
.B(net543),
.Y(net548)
);

XOR2x1_ASAP7_75t_R c567(
.A(net516),
.B(net510),
.Y(net549)
);

ICGx4DC_ASAP7_75t_R c568(
.ENA(net546),
.SE(net547),
.CLK(clk),
.GCLK(net550)
);

XOR2x2_ASAP7_75t_R c569(
.A(net540),
.B(net508),
.Y(net551)
);

INVx13_ASAP7_75t_R c570(
.A(net10139),
.Y(net552)
);

XOR2xp5_ASAP7_75t_R c571(
.A(net423),
.B(net10180),
.Y(net553)
);

AND2x2_ASAP7_75t_R c572(
.A(net513),
.B(net10181),
.Y(net554)
);

AND2x4_ASAP7_75t_R c573(
.A(net548),
.B(net553),
.Y(net555)
);

AOI21xp5_ASAP7_75t_R c574(
.A1(net555),
.A2(net10180),
.B(net10181),
.Y(net556)
);

AND2x6_ASAP7_75t_R c575(
.A(net322),
.B(net550),
.Y(net557)
);

INVx1_ASAP7_75t_R c576(
.A(net10117),
.Y(net558)
);

SDFLx1_ASAP7_75t_R c577(
.D(net478),
.SE(net546),
.SI(net558),
.CLK(clk),
.QN(net559)
);

FAx1_ASAP7_75t_R c578(
.A(net525),
.B(net465),
.CI(net555),
.SN(net561),
.CON(net560)
);

AOI321xp33_ASAP7_75t_R c579(
.A1(net552),
.A2(net472),
.A3(net560),
.B1(net558),
.B2(net534),
.C(net9948),
.Y(net562)
);

AOI33xp33_ASAP7_75t_R c580(
.A1(net479),
.A2(net554),
.A3(net559),
.B1(net493),
.B2(net558),
.B3(net10182),
.Y(net563)
);

INVx2_ASAP7_75t_R c581(
.A(net495),
.Y(net564)
);

INVx3_ASAP7_75t_R c582(
.A(net426),
.Y(net565)
);

INVx4_ASAP7_75t_R c583(
.A(net10421),
.Y(net566)
);

INVx5_ASAP7_75t_R c584(
.A(net476),
.Y(net567)
);

INVx6_ASAP7_75t_R c585(
.A(net356),
.Y(net568)
);

HAxp5_ASAP7_75t_R c586(
.A(net557),
.B(net538),
.CON(net569)
);

INVx8_ASAP7_75t_R c587(
.A(net9099),
.Y(net570)
);

NAND2x1_ASAP7_75t_R c588(
.A(net543),
.B(net427),
.Y(net571)
);

INVxp33_ASAP7_75t_R c589(
.A(net547),
.Y(net572)
);

INVxp67_ASAP7_75t_R c590(
.A(net486),
.Y(net573)
);

NAND2x1p5_ASAP7_75t_R c591(
.A(net529),
.B(net342),
.Y(net574)
);

BUFx10_ASAP7_75t_R c592(
.A(net87),
.Y(net575)
);

NAND2x2_ASAP7_75t_R c593(
.A(net488),
.B(net529),
.Y(net576)
);

BUFx12_ASAP7_75t_R c594(
.A(net79),
.Y(net577)
);

NAND2xp33_ASAP7_75t_R c595(
.A(net538),
.B(net566),
.Y(net578)
);

NAND2xp5_ASAP7_75t_R c596(
.A(net422),
.B(net559),
.Y(net579)
);

BUFx12f_ASAP7_75t_R c597(
.A(net448),
.Y(net580)
);

BUFx16f_ASAP7_75t_R c598(
.A(net342),
.Y(net581)
);

BUFx24_ASAP7_75t_R c599(
.A(net531),
.Y(net582)
);

BUFx2_ASAP7_75t_R c600(
.A(net576),
.Y(net583)
);

BUFx3_ASAP7_75t_R c601(
.A(net566),
.Y(net584)
);

BUFx4_ASAP7_75t_R c602(
.A(net9099),
.Y(net585)
);

BUFx4f_ASAP7_75t_R c603(
.A(net488),
.Y(net586)
);

BUFx5_ASAP7_75t_R c604(
.A(net572),
.Y(net587)
);

BUFx6f_ASAP7_75t_R c605(
.A(net577),
.Y(net588)
);

MAJIxp5_ASAP7_75t_R c606(
.A(net412),
.B(net578),
.C(net581),
.Y(net589)
);

NAND2xp67_ASAP7_75t_R c607(
.A(net448),
.B(net566),
.Y(net590)
);

BUFx8_ASAP7_75t_R c608(
.A(net476),
.Y(net591)
);

NOR2x1_ASAP7_75t_R c609(
.A(net583),
.B(net566),
.Y(net592)
);

CKINVDCx10_ASAP7_75t_R c610(
.A(net581),
.Y(net593)
);

CKINVDCx11_ASAP7_75t_R c611(
.A(net588),
.Y(net594)
);

CKINVDCx12_ASAP7_75t_R c612(
.A(net559),
.Y(net595)
);

CKINVDCx14_ASAP7_75t_R c613(
.A(net9228),
.Y(net596)
);

CKINVDCx16_ASAP7_75t_R c614(
.A(net593),
.Y(net597)
);

NOR2x1p5_ASAP7_75t_R c615(
.A(net583),
.B(net573),
.Y(net598)
);

NOR2x2_ASAP7_75t_R c616(
.A(net573),
.B(net553),
.Y(net599)
);

NOR2xp33_ASAP7_75t_R c617(
.A(net587),
.B(net517),
.Y(net600)
);

NOR2xp67_ASAP7_75t_R c618(
.A(net582),
.B(net587),
.Y(net601)
);

OR2x2_ASAP7_75t_R c619(
.A(net584),
.B(net601),
.Y(net602)
);

CKINVDCx20_ASAP7_75t_R c620(
.A(net519),
.Y(net603)
);

MAJx2_ASAP7_75t_R c621(
.A(net590),
.B(net594),
.C(net581),
.Y(net604)
);

CKINVDCx5p33_ASAP7_75t_R c622(
.A(net601),
.Y(net605)
);

OR2x4_ASAP7_75t_R c623(
.A(net571),
.B(net587),
.Y(net606)
);

CKINVDCx6p67_ASAP7_75t_R c624(
.A(net9251),
.Y(net607)
);

OR2x6_ASAP7_75t_R c625(
.A(net605),
.B(net342),
.Y(net608)
);

ICGx4_ASAP7_75t_R c626(
.ENA(net579),
.SE(net486),
.CLK(clk),
.GCLK(net609)
);

CKINVDCx8_ASAP7_75t_R c627(
.A(net565),
.Y(net610)
);

XNOR2x1_ASAP7_75t_R c628(
.B(net580),
.A(net574),
.Y(net611)
);

CKINVDCx9p33_ASAP7_75t_R c629(
.A(net587),
.Y(net612)
);

HB1xp67_ASAP7_75t_R c630(
.A(net609),
.Y(net613)
);

XNOR2x2_ASAP7_75t_R c631(
.A(net570),
.B(net561),
.Y(net614)
);

MAJx3_ASAP7_75t_R c632(
.A(net599),
.B(net541),
.C(net567),
.Y(net615)
);

XNOR2xp5_ASAP7_75t_R c633(
.A(net427),
.B(net582),
.Y(net616)
);

ICGx5_ASAP7_75t_R c634(
.ENA(net608),
.SE(net606),
.CLK(clk),
.GCLK(net617)
);

HB2xp67_ASAP7_75t_R c635(
.A(net575),
.Y(net618)
);

HB3xp67_ASAP7_75t_R c636(
.A(net9271),
.Y(net619)
);

NAND3x1_ASAP7_75t_R c637(
.A(net618),
.B(net573),
.C(net606),
.Y(net620)
);

HB4xp67_ASAP7_75t_R c638(
.A(net602),
.Y(net621)
);

INVx11_ASAP7_75t_R c639(
.A(net594),
.Y(net622)
);

INVx13_ASAP7_75t_R c640(
.A(net10506),
.Y(net623)
);

INVx1_ASAP7_75t_R c641(
.A(net597),
.Y(net624)
);

XOR2x1_ASAP7_75t_R c642(
.A(net603),
.B(net596),
.Y(net625)
);

XOR2x2_ASAP7_75t_R c643(
.A(net612),
.B(net608),
.Y(net626)
);

NAND3x2_ASAP7_75t_R c644(
.B(net543),
.C(net619),
.A(net612),
.Y(net627)
);

XOR2xp5_ASAP7_75t_R c645(
.A(net626),
.B(net604),
.Y(net628)
);

ICGx5p33DC_ASAP7_75t_R c646(
.ENA(net597),
.SE(net611),
.CLK(clk),
.GCLK(net629)
);

ICGx6p67DC_ASAP7_75t_R c647(
.ENA(net604),
.SE(net420),
.CLK(clk),
.GCLK(net630)
);

AND2x2_ASAP7_75t_R c648(
.A(net479),
.B(net619),
.Y(net631)
);

ICGx8DC_ASAP7_75t_R c649(
.ENA(net610),
.SE(net607),
.CLK(clk),
.GCLK(net632)
);

INVx2_ASAP7_75t_R c650(
.A(net596),
.Y(net633)
);

NAND3xp33_ASAP7_75t_R c651(
.A(net568),
.B(net565),
.C(net356),
.Y(net634)
);

SDFLx2_ASAP7_75t_R c652(
.D(net634),
.SE(net608),
.SI(net9934),
.CLK(clk),
.QN(net635)
);

INVx3_ASAP7_75t_R c653(
.A(net631),
.Y(net636)
);

NOR3x1_ASAP7_75t_R c654(
.A(net636),
.B(net632),
.C(net611),
.Y(net637)
);

INVx4_ASAP7_75t_R c655(
.A(net623),
.Y(net638)
);

AND2x4_ASAP7_75t_R c656(
.A(net621),
.B(net630),
.Y(net639)
);

NOR3x2_ASAP7_75t_R c657(
.B(net612),
.C(net636),
.A(net639),
.Y(net640)
);

NOR3xp33_ASAP7_75t_R c658(
.A(net422),
.B(net519),
.C(net608),
.Y(net641)
);

AOI221xp5_ASAP7_75t_R c659(
.A1(net187),
.A2(net634),
.B1(net575),
.B2(net574),
.C(net587),
.Y(net642)
);

OA21x2_ASAP7_75t_R c660(
.A1(net569),
.A2(net615),
.B(net543),
.Y(net643)
);

SDFLx3_ASAP7_75t_R c661(
.D(net566),
.SE(net640),
.SI(net589),
.CLK(clk),
.QN(net644)
);

OAI21x1_ASAP7_75t_R c662(
.A1(net339),
.A2(net639),
.B(net616),
.Y(net645)
);

AO31x2_ASAP7_75t_R c663(
.A1(net615),
.A2(net635),
.A3(net633),
.B(net644),
.Y(net646)
);

INVx5_ASAP7_75t_R c664(
.A(net10150),
.Y(net647)
);

INVx6_ASAP7_75t_R c665(
.A(net10182),
.Y(net648)
);

INVx8_ASAP7_75t_R c666(
.A(net591),
.Y(net649)
);

AND2x6_ASAP7_75t_R c667(
.A(net245),
.B(net629),
.Y(net650)
);

INVxp33_ASAP7_75t_R c668(
.A(net648),
.Y(net651)
);

INVxp67_ASAP7_75t_R c669(
.A(net452),
.Y(net652)
);

BUFx10_ASAP7_75t_R c670(
.A(net627),
.Y(net653)
);

BUFx12_ASAP7_75t_R c671(
.A(net10480),
.Y(net654)
);

BUFx12f_ASAP7_75t_R c672(
.A(net650),
.Y(net655)
);

BUFx16f_ASAP7_75t_R c673(
.A(net10150),
.Y(net656)
);

BUFx24_ASAP7_75t_R c674(
.A(net591),
.Y(net657)
);

BUFx2_ASAP7_75t_R c675(
.A(net9224),
.Y(net658)
);

HAxp5_ASAP7_75t_R c676(
.A(net619),
.B(net635),
.CON(net660),
.SN(net659)
);

BUFx3_ASAP7_75t_R c677(
.A(net592),
.Y(net661)
);

BUFx4_ASAP7_75t_R c678(
.A(net10017),
.Y(net662)
);

BUFx4f_ASAP7_75t_R c679(
.A(net653),
.Y(net663)
);

NAND2x1_ASAP7_75t_R c680(
.A(net636),
.B(net567),
.Y(net664)
);

BUFx5_ASAP7_75t_R c681(
.A(net618),
.Y(net665)
);

BUFx6f_ASAP7_75t_R c682(
.A(net353),
.Y(net666)
);

BUFx8_ASAP7_75t_R c683(
.A(net619),
.Y(net667)
);

CKINVDCx10_ASAP7_75t_R c684(
.A(net9273),
.Y(net668)
);

CKINVDCx11_ASAP7_75t_R c685(
.A(net631),
.Y(net669)
);

NAND2x1p5_ASAP7_75t_R c686(
.A(net592),
.B(net10017),
.Y(net670)
);

CKINVDCx12_ASAP7_75t_R c687(
.A(net670),
.Y(net671)
);

CKINVDCx14_ASAP7_75t_R c688(
.A(net648),
.Y(net672)
);

NAND2x2_ASAP7_75t_R c689(
.A(net624),
.B(net567),
.Y(net673)
);

CKINVDCx16_ASAP7_75t_R c690(
.A(net567),
.Y(net674)
);

CKINVDCx20_ASAP7_75t_R c691(
.A(net669),
.Y(net675)
);

CKINVDCx5p33_ASAP7_75t_R c692(
.A(net655),
.Y(net676)
);

CKINVDCx6p67_ASAP7_75t_R c693(
.A(net508),
.Y(net677)
);

NAND2xp33_ASAP7_75t_R c694(
.A(net644),
.B(net649),
.Y(net678)
);

CKINVDCx8_ASAP7_75t_R c695(
.A(net674),
.Y(net679)
);

CKINVDCx9p33_ASAP7_75t_R c696(
.A(net639),
.Y(net680)
);

HB1xp67_ASAP7_75t_R c697(
.A(net670),
.Y(net681)
);

HB2xp67_ASAP7_75t_R c698(
.A(net660),
.Y(net682)
);

HB3xp67_ASAP7_75t_R c699(
.A(net679),
.Y(net683)
);

NAND2xp5_ASAP7_75t_R c700(
.A(net654),
.B(net669),
.Y(net684)
);

HB4xp67_ASAP7_75t_R c701(
.A(net668),
.Y(net685)
);

INVx11_ASAP7_75t_R c702(
.A(net9273),
.Y(net686)
);

NAND2xp67_ASAP7_75t_R c703(
.A(net675),
.B(net655),
.Y(net687)
);

NOR2x1_ASAP7_75t_R c704(
.A(net684),
.B(net669),
.Y(net688)
);

INVx13_ASAP7_75t_R c705(
.A(net571),
.Y(net689)
);

INVx1_ASAP7_75t_R c706(
.A(net665),
.Y(net690)
);

NOR2x1p5_ASAP7_75t_R c707(
.A(net683),
.B(net680),
.Y(net691)
);

NOR2x2_ASAP7_75t_R c708(
.A(net690),
.B(net651),
.Y(net692)
);

AOI311xp33_ASAP7_75t_R c709(
.A1(net635),
.A2(net644),
.A3(net667),
.B(net686),
.C(net10182),
.Y(net693)
);

INVx2_ASAP7_75t_R c710(
.A(net10540),
.Y(net694)
);

NOR2xp33_ASAP7_75t_R c711(
.A(net657),
.B(net633),
.Y(net695)
);

INVx3_ASAP7_75t_R c712(
.A(net694),
.Y(net696)
);

INVx4_ASAP7_75t_R c713(
.A(net684),
.Y(net697)
);

NOR2xp67_ASAP7_75t_R c714(
.A(net663),
.B(net687),
.Y(net698)
);

OAI21xp33_ASAP7_75t_R c715(
.A1(net696),
.A2(net656),
.B(net670),
.Y(net699)
);

OR2x2_ASAP7_75t_R c716(
.A(net698),
.B(net574),
.Y(net700)
);

OR2x4_ASAP7_75t_R c717(
.A(net699),
.B(net692),
.Y(net701)
);

INVx5_ASAP7_75t_R c718(
.A(net682),
.Y(net702)
);

INVx6_ASAP7_75t_R c719(
.A(net693),
.Y(net703)
);

OR2x6_ASAP7_75t_R c720(
.A(net689),
.B(net650),
.Y(net704)
);

INVx8_ASAP7_75t_R c721(
.A(net652),
.Y(net705)
);

XNOR2x1_ASAP7_75t_R c722(
.B(net678),
.A(net700),
.Y(net706)
);

OAI21xp5_ASAP7_75t_R c723(
.A1(net420),
.A2(net685),
.B(net674),
.Y(net707)
);

OR3x1_ASAP7_75t_R c724(
.A(net342),
.B(net695),
.C(net10183),
.Y(net708)
);

INVxp33_ASAP7_75t_R c725(
.A(net676),
.Y(net709)
);

OR3x2_ASAP7_75t_R c726(
.A(net692),
.B(net600),
.C(net700),
.Y(net710)
);

ICGx1_ASAP7_75t_R c727(
.ENA(net701),
.SE(net710),
.CLK(clk),
.GCLK(net711)
);

AOI32xp33_ASAP7_75t_R c728(
.A1(net607),
.A2(net564),
.A3(net567),
.B1(net688),
.B2(net686),
.Y(net712)
);

OR3x4_ASAP7_75t_R c729(
.A(net695),
.B(net677),
.C(net661),
.Y(net713)
);

INVxp67_ASAP7_75t_R c730(
.A(net10476),
.Y(net714)
);

BUFx10_ASAP7_75t_R c731(
.A(net713),
.Y(net715)
);

XNOR2x2_ASAP7_75t_R c732(
.A(net666),
.B(net708),
.Y(net716)
);

XNOR2xp5_ASAP7_75t_R c733(
.A(net685),
.B(net714),
.Y(net717)
);

AND3x1_ASAP7_75t_R c734(
.A(net549),
.B(net651),
.C(net10184),
.Y(net718)
);

XOR2x1_ASAP7_75t_R c735(
.A(net649),
.B(net705),
.Y(net719)
);

BUFx12_ASAP7_75t_R c736(
.A(net691),
.Y(net720)
);

BUFx12f_ASAP7_75t_R c737(
.A(net719),
.Y(net721)
);

BUFx16f_ASAP7_75t_R c738(
.A(net717),
.Y(net722)
);

XOR2x2_ASAP7_75t_R c739(
.A(net707),
.B(net556),
.Y(net723)
);

AND3x2_ASAP7_75t_R c740(
.A(net708),
.B(net723),
.C(net10034),
.Y(net724)
);

BUFx24_ASAP7_75t_R c741(
.A(net723),
.Y(net725)
);

AND3x4_ASAP7_75t_R c742(
.A(net715),
.B(net690),
.C(net724),
.Y(net726)
);

AOI211x1_ASAP7_75t_R c743(
.A1(net725),
.A2(net682),
.B(net726),
.C(net693),
.Y(net727)
);

NAND5xp2_ASAP7_75t_R c744(
.A(net718),
.B(net725),
.C(net665),
.D(net633),
.E(net10184),
.Y(net728)
);

NOR5xp2_ASAP7_75t_R c745(
.A(net706),
.B(net727),
.C(net720),
.D(net726),
.E(net708),
.Y(net729)
);

XOR2xp5_ASAP7_75t_R c746(
.A(net724),
.B(net10034),
.Y(net730)
);

AND2x2_ASAP7_75t_R c747(
.A(net325),
.B(net680),
.Y(net731)
);

BUFx2_ASAP7_75t_R c748(
.A(net10376),
.Y(net732)
);

BUFx3_ASAP7_75t_R c749(
.A(net697),
.Y(net733)
);

BUFx4_ASAP7_75t_R c750(
.A(net633),
.Y(net734)
);

AND2x4_ASAP7_75t_R c751(
.A(net483),
.B(net733),
.Y(net735)
);

BUFx4f_ASAP7_75t_R c752(
.A(net720),
.Y(net736)
);

AND2x6_ASAP7_75t_R c753(
.A(net688),
.B(net10176),
.Y(net737)
);

BUFx5_ASAP7_75t_R c754(
.A(net688),
.Y(net738)
);

BUFx6f_ASAP7_75t_R c755(
.A(net600),
.Y(net739)
);

BUFx8_ASAP7_75t_R c756(
.A(net630),
.Y(net740)
);

AO21x1_ASAP7_75t_R c757(
.A1(net272),
.A2(net512),
.B(net740),
.Y(net741)
);

CKINVDCx10_ASAP7_75t_R c758(
.A(net734),
.Y(net742)
);

AO21x2_ASAP7_75t_R c759(
.A1(net724),
.A2(net617),
.B(net664),
.Y(net743)
);

CKINVDCx11_ASAP7_75t_R c760(
.A(net600),
.Y(net744)
);

CKINVDCx12_ASAP7_75t_R c761(
.A(net739),
.Y(net745)
);

CKINVDCx14_ASAP7_75t_R c762(
.A(net711),
.Y(net746)
);

HAxp5_ASAP7_75t_R c763(
.A(net72),
.B(net734),
.CON(net748),
.SN(net747)
);

NAND2x1_ASAP7_75t_R c764(
.A(net733),
.B(net686),
.Y(net749)
);

CKINVDCx16_ASAP7_75t_R c765(
.A(net595),
.Y(net750)
);

CKINVDCx20_ASAP7_75t_R c766(
.A(net750),
.Y(net751)
);

CKINVDCx5p33_ASAP7_75t_R c767(
.A(net10183),
.Y(net752)
);

CKINVDCx6p67_ASAP7_75t_R c768(
.A(net627),
.Y(net753)
);

CKINVDCx8_ASAP7_75t_R c769(
.A(net702),
.Y(net754)
);

CKINVDCx9p33_ASAP7_75t_R c770(
.A(net595),
.Y(net755)
);

HB1xp67_ASAP7_75t_R c771(
.A(net680),
.Y(net756)
);

HB2xp67_ASAP7_75t_R c772(
.A(net746),
.Y(net757)
);

NAND2x1p5_ASAP7_75t_R c773(
.A(net59),
.B(net756),
.Y(net758)
);

NAND2x2_ASAP7_75t_R c774(
.A(net744),
.B(net753),
.Y(net759)
);

HB3xp67_ASAP7_75t_R c775(
.A(net740),
.Y(net760)
);

HB4xp67_ASAP7_75t_R c776(
.A(net709),
.Y(net761)
);

INVx11_ASAP7_75t_R c777(
.A(net752),
.Y(net762)
);

NAND2xp33_ASAP7_75t_R c778(
.A(net737),
.B(net742),
.Y(net763)
);

INVx13_ASAP7_75t_R c779(
.A(net9170),
.Y(net764)
);

NAND2xp5_ASAP7_75t_R c780(
.A(net617),
.B(net755),
.Y(net765)
);

NAND2xp67_ASAP7_75t_R c781(
.A(net759),
.B(net697),
.Y(net766)
);

INVx1_ASAP7_75t_R c782(
.A(net756),
.Y(net767)
);

NOR2x1_ASAP7_75t_R c783(
.A(net761),
.B(net762),
.Y(net768)
);

INVx2_ASAP7_75t_R c784(
.A(net755),
.Y(net769)
);

AOI21x1_ASAP7_75t_R c785(
.A1(net767),
.A2(net758),
.B(net697),
.Y(net770)
);

INVx3_ASAP7_75t_R c786(
.A(net751),
.Y(net771)
);

NOR2x1p5_ASAP7_75t_R c787(
.A(net617),
.B(net710),
.Y(net772)
);

NOR2x2_ASAP7_75t_R c788(
.A(net687),
.B(net764),
.Y(net773)
);

NOR2xp33_ASAP7_75t_R c789(
.A(net766),
.B(net9657),
.Y(net774)
);

INVx4_ASAP7_75t_R c790(
.A(net753),
.Y(net775)
);

INVx5_ASAP7_75t_R c791(
.A(net771),
.Y(net776)
);

INVx6_ASAP7_75t_R c792(
.A(out0),
.Y(net777)
);

INVx8_ASAP7_75t_R c793(
.A(net765),
.Y(net778)
);

NOR2xp67_ASAP7_75t_R c794(
.A(net751),
.B(net736),
.Y(net779)
);

OR2x2_ASAP7_75t_R c795(
.A(net688),
.B(net709),
.Y(net780)
);

INVxp33_ASAP7_75t_R c796(
.A(net757),
.Y(net781)
);

INVxp67_ASAP7_75t_R c797(
.A(net767),
.Y(net782)
);

OR2x4_ASAP7_75t_R c798(
.A(net732),
.B(net755),
.Y(net783)
);

BUFx10_ASAP7_75t_R c799(
.A(net9952),
.Y(net784)
);

ICGx2_ASAP7_75t_R c800(
.ENA(net762),
.SE(net782),
.CLK(clk),
.GCLK(net785)
);

BUFx12_ASAP7_75t_R c801(
.A(net9170),
.Y(net786)
);

OR2x6_ASAP7_75t_R c802(
.A(net766),
.B(net771),
.Y(net787)
);

BUFx12f_ASAP7_75t_R c803(
.A(net731),
.Y(net788)
);

AOI211xp5_ASAP7_75t_R c804(
.A1(net774),
.A2(net783),
.B(net762),
.C(net784),
.Y(net789)
);

XNOR2x1_ASAP7_75t_R c805(
.B(net739),
.A(net780),
.Y(net790)
);

XNOR2x2_ASAP7_75t_R c806(
.A(net745),
.B(net627),
.Y(net791)
);

BUFx16f_ASAP7_75t_R c807(
.A(net9657),
.Y(net792)
);

BUFx24_ASAP7_75t_R c808(
.A(net769),
.Y(net793)
);

XNOR2xp5_ASAP7_75t_R c809(
.A(net681),
.B(net790),
.Y(net794)
);

XOR2x1_ASAP7_75t_R c810(
.A(net758),
.B(net790),
.Y(net795)
);

AOI22x1_ASAP7_75t_R c811(
.A1(net761),
.A2(net784),
.B1(net758),
.B2(net789),
.Y(net796)
);

OA221x2_ASAP7_75t_R c812(
.A1(net783),
.A2(net789),
.B1(net627),
.B2(net755),
.C(net787),
.Y(net797)
);

XOR2x2_ASAP7_75t_R c813(
.A(net744),
.B(net786),
.Y(net798)
);

BUFx2_ASAP7_75t_R c814(
.A(net10392),
.Y(net799)
);

XOR2xp5_ASAP7_75t_R c815(
.A(net658),
.B(net787),
.Y(net800)
);

AND2x2_ASAP7_75t_R c816(
.A(net768),
.B(net793),
.Y(net801)
);

AND2x4_ASAP7_75t_R c817(
.A(net801),
.B(net798),
.Y(net802)
);

ICGx2p67DC_ASAP7_75t_R c818(
.ENA(net797),
.SE(net799),
.CLK(clk),
.GCLK(net803)
);

AND2x6_ASAP7_75t_R c819(
.A(net793),
.B(net680),
.Y(net804)
);

SDFLx4_ASAP7_75t_R c820(
.D(net795),
.SE(net802),
.SI(net749),
.CLK(clk),
.QN(net805)
);

OAI221xp5_ASAP7_75t_R c821(
.A1(net802),
.A2(net781),
.B1(net767),
.B2(net789),
.C(net801),
.Y(net806)
);

AOI21xp33_ASAP7_75t_R c822(
.A1(net776),
.A2(net790),
.B(net803),
.Y(net807)
);

DFFASRHQNx1_ASAP7_75t_R c823(
.D(net806),
.RESETN(net778),
.SETN(net769),
.CLK(clk),
.QN(net808)
);

AOI21xp5_ASAP7_75t_R c824(
.A1(net808),
.A2(net633),
.B(net764),
.Y(net809)
);

OAI311xp33_ASAP7_75t_R c825(
.A1(net794),
.A2(net805),
.A3(net807),
.B1(net742),
.C1(net803),
.Y(net810)
);

AOI22xp33_ASAP7_75t_R c826(
.A1(net796),
.A2(net766),
.B1(net806),
.B2(net789),
.Y(net811)
);

HAxp5_ASAP7_75t_R c827(
.A(net800),
.B(net774),
.CON(net813),
.SN(net812)
);

NAND2x1_ASAP7_75t_R c828(
.A(net804),
.B(net781),
.Y(net814)
);

OAI32xp33_ASAP7_75t_R c829(
.A1(net814),
.A2(net807),
.A3(net812),
.B1(net789),
.B2(net738),
.Y(net815)
);

BUFx3_ASAP7_75t_R c830(
.A(net789),
.Y(net816)
);

BUFx4_ASAP7_75t_R c831(
.A(net9125),
.Y(net817)
);

BUFx4f_ASAP7_75t_R c832(
.A(net445),
.Y(net818)
);

NAND2x1p5_ASAP7_75t_R c833(
.A(net561),
.B(net531),
.Y(net819)
);

BUFx5_ASAP7_75t_R c834(
.A(net339),
.Y(net820)
);

BUFx6f_ASAP7_75t_R c835(
.A(net818),
.Y(net821)
);

BUFx8_ASAP7_75t_R c836(
.A(net818),
.Y(net822)
);

CKINVDCx10_ASAP7_75t_R c837(
.A(net820),
.Y(net823)
);

CKINVDCx11_ASAP7_75t_R c838(
.A(net819),
.Y(net824)
);

NAND2x2_ASAP7_75t_R c839(
.A(net788),
.B(net787),
.Y(net825)
);

CKINVDCx12_ASAP7_75t_R c840(
.A(net822),
.Y(net826)
);

CKINVDCx14_ASAP7_75t_R c841(
.A(net785),
.Y(net827)
);

NAND2xp33_ASAP7_75t_R c842(
.A(net827),
.B(net825),
.Y(net828)
);

CKINVDCx16_ASAP7_75t_R c843(
.A(net9666),
.Y(net829)
);

CKINVDCx20_ASAP7_75t_R c844(
.A(net9125),
.Y(net830)
);

CKINVDCx5p33_ASAP7_75t_R c845(
.A(net791),
.Y(net831)
);

NAND2xp5_ASAP7_75t_R c846(
.A(net720),
.B(net609),
.Y(net832)
);

SDFHx1_ASAP7_75t_R c847(
.D(net832),
.SE(net791),
.SI(net10185),
.CLK(clk),
.QN(net833)
);

CKINVDCx6p67_ASAP7_75t_R c848(
.A(net820),
.Y(net834)
);

CKINVDCx8_ASAP7_75t_R c849(
.A(net726),
.Y(net835)
);

SDFHx2_ASAP7_75t_R c850(
.D(net823),
.SE(net833),
.SI(net736),
.CLK(clk),
.QN(net836)
);

CKINVDCx9p33_ASAP7_75t_R c851(
.A(net754),
.Y(net837)
);

FAx1_ASAP7_75t_R c852(
.A(net833),
.B(net753),
.CI(net10185),
.SN(net839),
.CON(net838)
);

HB1xp67_ASAP7_75t_R c853(
.A(net780),
.Y(net840)
);

HB2xp67_ASAP7_75t_R c854(
.A(net837),
.Y(net841)
);

HB3xp67_ASAP7_75t_R c855(
.A(net829),
.Y(net842)
);

HB4xp67_ASAP7_75t_R c856(
.A(net826),
.Y(net843)
);

INVx11_ASAP7_75t_R c857(
.A(net742),
.Y(net844)
);

INVx13_ASAP7_75t_R c858(
.A(net788),
.Y(net845)
);

INVx1_ASAP7_75t_R c859(
.A(net819),
.Y(net846)
);

NAND2xp67_ASAP7_75t_R c860(
.A(net672),
.B(net742),
.Y(net847)
);

NOR2x1_ASAP7_75t_R c861(
.A(net697),
.B(net743),
.Y(net848)
);

NOR2x1p5_ASAP7_75t_R c862(
.A(net829),
.B(net781),
.Y(net849)
);

NOR2x2_ASAP7_75t_R c863(
.A(net844),
.B(net789),
.Y(net850)
);

NOR2xp33_ASAP7_75t_R c864(
.A(net498),
.B(net749),
.Y(net851)
);

NOR2xp67_ASAP7_75t_R c865(
.A(net849),
.B(net749),
.Y(net852)
);

INVx2_ASAP7_75t_R c866(
.A(net843),
.Y(net853)
);

INVx3_ASAP7_75t_R c867(
.A(net9265),
.Y(net854)
);

MAJIxp5_ASAP7_75t_R c868(
.A(net821),
.B(net853),
.C(net713),
.Y(net855)
);

AOI22xp5_ASAP7_75t_R c869(
.A1(net843),
.A2(net818),
.B1(net803),
.B2(net10179),
.Y(net856)
);

INVx4_ASAP7_75t_R c870(
.A(net713),
.Y(net857)
);

INVx5_ASAP7_75t_R c871(
.A(net10511),
.Y(net858)
);

OR2x2_ASAP7_75t_R c872(
.A(net842),
.B(net827),
.Y(net859)
);

INVx6_ASAP7_75t_R c873(
.A(net831),
.Y(net860)
);

INVx8_ASAP7_75t_R c874(
.A(net827),
.Y(net861)
);

OR2x4_ASAP7_75t_R c875(
.A(net853),
.B(net860),
.Y(net862)
);

INVxp33_ASAP7_75t_R c876(
.A(net9265),
.Y(net863)
);

INVxp67_ASAP7_75t_R c877(
.A(net856),
.Y(net864)
);

MAJx2_ASAP7_75t_R c878(
.A(net837),
.B(net860),
.C(net843),
.Y(net865)
);

ICGx3_ASAP7_75t_R c879(
.ENA(net850),
.SE(net863),
.CLK(clk),
.GCLK(net866)
);

MAJx3_ASAP7_75t_R c880(
.A(net534),
.B(net803),
.C(net609),
.Y(net867)
);

BUFx10_ASAP7_75t_R c881(
.A(net857),
.Y(net868)
);

BUFx12_ASAP7_75t_R c882(
.A(net858),
.Y(net869)
);

OR2x6_ASAP7_75t_R c883(
.A(net864),
.B(net851),
.Y(net870)
);

XNOR2x1_ASAP7_75t_R c884(
.B(net846),
.A(net10185),
.Y(net871)
);

XNOR2x2_ASAP7_75t_R c885(
.A(net869),
.B(net842),
.Y(net872)
);

XNOR2xp5_ASAP7_75t_R c886(
.A(net817),
.B(net780),
.Y(net873)
);

BUFx12f_ASAP7_75t_R c887(
.A(net834),
.Y(net874)
);

XOR2x1_ASAP7_75t_R c888(
.A(net841),
.B(net754),
.Y(net875)
);

BUFx16f_ASAP7_75t_R c889(
.A(net875),
.Y(net876)
);

BUFx24_ASAP7_75t_R c890(
.A(net830),
.Y(net877)
);

NAND3x1_ASAP7_75t_R c891(
.A(net840),
.B(net787),
.C(net870),
.Y(net878)
);

NAND3x2_ASAP7_75t_R c892(
.B(net789),
.C(net856),
.A(net843),
.Y(net879)
);

BUFx2_ASAP7_75t_R c893(
.A(net872),
.Y(net880)
);

BUFx3_ASAP7_75t_R c894(
.A(net9666),
.Y(net881)
);

BUFx4_ASAP7_75t_R c895(
.A(net9224),
.Y(net882)
);

BUFx4f_ASAP7_75t_R c896(
.A(net10480),
.Y(net883)
);

NAND3xp33_ASAP7_75t_R c897(
.A(net878),
.B(net860),
.C(net753),
.Y(net884)
);

XOR2x2_ASAP7_75t_R c898(
.A(net753),
.B(net851),
.Y(net885)
);

NOR3x1_ASAP7_75t_R c899(
.A(net833),
.B(net726),
.C(net9984),
.Y(net886)
);

XOR2xp5_ASAP7_75t_R c900(
.A(net877),
.B(net9984),
.Y(net887)
);

BUFx5_ASAP7_75t_R c901(
.A(net10514),
.Y(net888)
);

OA222x2_ASAP7_75t_R c902(
.A1(net882),
.A2(net884),
.B1(net853),
.B2(net860),
.C1(net849),
.C2(net837),
.Y(net889)
);

AND2x2_ASAP7_75t_R c903(
.A(net887),
.B(net885),
.Y(net890)
);

BUFx6f_ASAP7_75t_R c904(
.A(net890),
.Y(net891)
);

BUFx8_ASAP7_75t_R c905(
.A(net10087),
.Y(net892)
);

NOR3x2_ASAP7_75t_R c906(
.B(net883),
.C(net892),
.A(net859),
.Y(net893)
);

AND2x4_ASAP7_75t_R c907(
.A(net855),
.B(net781),
.Y(net894)
);

NOR3xp33_ASAP7_75t_R c908(
.A(net888),
.B(net891),
.C(net881),
.Y(net895)
);

OR5x1_ASAP7_75t_R c909(
.A(net862),
.B(net836),
.C(net893),
.D(net849),
.E(net534),
.Y(net896)
);

SDFHx3_ASAP7_75t_R c910(
.D(net877),
.SE(net892),
.SI(net850),
.CLK(clk),
.QN(net897)
);

OA21x2_ASAP7_75t_R c911(
.A1(net859),
.A2(net876),
.B(net9812),
.Y(net898)
);

AND2x6_ASAP7_75t_R c912(
.A(net898),
.B(net9791),
.Y(net899)
);

CKINVDCx10_ASAP7_75t_R c913(
.A(net36),
.Y(net900)
);

CKINVDCx11_ASAP7_75t_R c914(
.A(net9),
.Y(net901)
);

CKINVDCx12_ASAP7_75t_R c915(
.A(net52),
.Y(net902)
);

CKINVDCx14_ASAP7_75t_R c916(
.A(net27),
.Y(net903)
);

CKINVDCx16_ASAP7_75t_R c917(
.A(net49),
.Y(net904)
);

CKINVDCx20_ASAP7_75t_R c918(
.A(net6),
.Y(net905)
);

CKINVDCx5p33_ASAP7_75t_R c919(
.A(net48),
.Y(net906)
);

CKINVDCx6p67_ASAP7_75t_R c920(
.A(in23),
.Y(net907)
);

CKINVDCx8_ASAP7_75t_R c921(
.A(in5),
.Y(net908)
);

CKINVDCx9p33_ASAP7_75t_R c922(
.A(net20),
.Y(net909)
);

HB1xp67_ASAP7_75t_R c923(
.A(net6),
.Y(net910)
);

HAxp5_ASAP7_75t_R c924(
.A(in12),
.B(net52),
.CON(net912),
.SN(net911)
);

HB2xp67_ASAP7_75t_R c925(
.A(net904),
.Y(net913)
);

HB3xp67_ASAP7_75t_R c926(
.A(net9181),
.Y(net914)
);

HB4xp67_ASAP7_75t_R c927(
.A(net53),
.Y(net915)
);

INVx11_ASAP7_75t_R c928(
.A(net9181),
.Y(net916)
);

NAND2x1_ASAP7_75t_R c929(
.A(in19),
.B(net910),
.Y(net917)
);

INVx13_ASAP7_75t_R c930(
.A(net912),
.Y(net918)
);

INVx1_ASAP7_75t_R c931(
.A(in13),
.Y(net919)
);

INVx2_ASAP7_75t_R c932(
.A(net911),
.Y(net920)
);

INVx3_ASAP7_75t_R c933(
.A(net916),
.Y(net921)
);

INVx4_ASAP7_75t_R c934(
.A(in19),
.Y(net922)
);

INVx5_ASAP7_75t_R c935(
.A(net919),
.Y(net923)
);

NAND2x1p5_ASAP7_75t_R c936(
.A(net918),
.B(net920),
.Y(net924)
);

INVx6_ASAP7_75t_R c937(
.A(net916),
.Y(net925)
);

INVx8_ASAP7_75t_R c938(
.A(net925),
.Y(net926)
);

NAND2x2_ASAP7_75t_R c939(
.A(net20),
.B(net917),
.Y(net927)
);

INVxp33_ASAP7_75t_R c940(
.A(net48),
.Y(net928)
);

INVxp67_ASAP7_75t_R c941(
.A(in7),
.Y(net929)
);

BUFx10_ASAP7_75t_R c942(
.A(net909),
.Y(net930)
);

BUFx12_ASAP7_75t_R c943(
.A(net930),
.Y(net931)
);

BUFx12f_ASAP7_75t_R c944(
.A(net908),
.Y(net932)
);

BUFx16f_ASAP7_75t_R c945(
.A(net51),
.Y(net933)
);

BUFx24_ASAP7_75t_R c946(
.A(net933),
.Y(net934)
);

OAI21x1_ASAP7_75t_R c947(
.A1(net920),
.A2(net925),
.B(net932),
.Y(net935)
);

BUFx2_ASAP7_75t_R c948(
.A(net931),
.Y(net936)
);

NAND2xp33_ASAP7_75t_R c949(
.A(net53),
.B(net922),
.Y(net937)
);

BUFx3_ASAP7_75t_R c950(
.A(in9),
.Y(net938)
);

BUFx4_ASAP7_75t_R c951(
.A(net917),
.Y(net939)
);

BUFx4f_ASAP7_75t_R c952(
.A(net52),
.Y(net940)
);

BUFx5_ASAP7_75t_R c953(
.A(net938),
.Y(net941)
);

NAND2xp5_ASAP7_75t_R c954(
.A(net903),
.B(net940),
.Y(net942)
);

NAND2xp67_ASAP7_75t_R c955(
.A(net939),
.B(net942),
.Y(net943)
);

BUFx6f_ASAP7_75t_R c956(
.A(net934),
.Y(net944)
);

NOR2x1_ASAP7_75t_R c957(
.A(net935),
.B(net941),
.Y(net945)
);

NOR2x1p5_ASAP7_75t_R c958(
.A(net909),
.B(net930),
.Y(net946)
);

OAI21xp33_ASAP7_75t_R c959(
.A1(net918),
.A2(net933),
.B(net935),
.Y(net947)
);

NOR2x2_ASAP7_75t_R c960(
.A(net929),
.B(net923),
.Y(net948)
);

BUFx8_ASAP7_75t_R c961(
.A(net936),
.Y(net949)
);

OAI21xp5_ASAP7_75t_R c962(
.A1(in15),
.A2(net6),
.B(net907),
.Y(net950)
);

CKINVDCx10_ASAP7_75t_R c963(
.A(net948),
.Y(net951)
);

NOR2xp33_ASAP7_75t_R c964(
.A(net947),
.B(net6),
.Y(net952)
);

CKINVDCx11_ASAP7_75t_R c965(
.A(net937),
.Y(net953)
);

NOR2xp67_ASAP7_75t_R c966(
.A(net946),
.B(net936),
.Y(net954)
);

OR2x2_ASAP7_75t_R c967(
.A(net914),
.B(net949),
.Y(net955)
);

OR2x4_ASAP7_75t_R c968(
.A(net910),
.B(in23),
.Y(net956)
);

OR2x6_ASAP7_75t_R c969(
.A(net901),
.B(net951),
.Y(net957)
);

XNOR2x1_ASAP7_75t_R c970(
.B(net944),
.A(net953),
.Y(net958)
);

OR3x1_ASAP7_75t_R c971(
.A(net935),
.B(net914),
.C(net925),
.Y(net959)
);

XNOR2x2_ASAP7_75t_R c972(
.A(net904),
.B(net926),
.Y(net960)
);

XNOR2xp5_ASAP7_75t_R c973(
.A(net957),
.B(net948),
.Y(net961)
);

CKINVDCx12_ASAP7_75t_R c974(
.A(net926),
.Y(net962)
);

CKINVDCx14_ASAP7_75t_R c975(
.A(net956),
.Y(net963)
);

CKINVDCx16_ASAP7_75t_R c976(
.A(net961),
.Y(net964)
);

CKINVDCx20_ASAP7_75t_R c977(
.A(in9),
.Y(net965)
);

OR3x2_ASAP7_75t_R c978(
.A(net963),
.B(net964),
.C(net929),
.Y(net966)
);

XOR2x1_ASAP7_75t_R c979(
.A(net923),
.B(net935),
.Y(net967)
);

CKINVDCx5p33_ASAP7_75t_R c980(
.A(in12),
.Y(net968)
);

CKINVDCx6p67_ASAP7_75t_R c981(
.A(net953),
.Y(net969)
);

XOR2x2_ASAP7_75t_R c982(
.A(net942),
.B(net944),
.Y(net970)
);

XOR2xp5_ASAP7_75t_R c983(
.A(net969),
.B(net961),
.Y(net971)
);

AND2x2_ASAP7_75t_R c984(
.A(net970),
.B(net967),
.Y(net972)
);

OR3x4_ASAP7_75t_R c985(
.A(net940),
.B(net36),
.C(net960),
.Y(net973)
);

AND2x4_ASAP7_75t_R c986(
.A(net951),
.B(net930),
.Y(net974)
);

AND2x6_ASAP7_75t_R c987(
.A(net962),
.B(net9704),
.Y(net975)
);

OA33x2_ASAP7_75t_R c988(
.A1(net963),
.A2(net907),
.A3(net950),
.B1(net975),
.B2(net932),
.B3(net9704),
.Y(net976)
);

HAxp5_ASAP7_75t_R c989(
.A(net906),
.B(net9704),
.CON(net978),
.SN(net977)
);

OR5x2_ASAP7_75t_R c990(
.A(net971),
.B(net976),
.C(net932),
.D(net907),
.E(net9704),
.Y(net979)
);

ICGx4DC_ASAP7_75t_R c991(
.ENA(net960),
.SE(net974),
.CLK(clk),
.GCLK(net980)
);

NAND2x1_ASAP7_75t_R c992(
.A(net974),
.B(net938),
.Y(net981)
);

AOI31xp33_ASAP7_75t_R c993(
.A1(net976),
.A2(net981),
.A3(net971),
.B(net975),
.Y(net982)
);

AOI31xp67_ASAP7_75t_R c994(
.A1(net981),
.A2(net967),
.A3(net971),
.B(net925),
.Y(net983)
);

NAND4xp25_ASAP7_75t_R c995(
.A(net955),
.B(net959),
.C(net981),
.D(net925),
.Y(net984)
);

AND3x1_ASAP7_75t_R c996(
.A(net1039),
.B(net1037),
.C(net913),
.Y(net985)
);

CKINVDCx8_ASAP7_75t_R c997(
.A(net954),
.Y(net986)
);

NAND2x1p5_ASAP7_75t_R c998(
.A(net1041),
.B(net54),
.Y(net987)
);

NAND2x2_ASAP7_75t_R c999(
.A(net109),
.B(net949),
.Y(net988)
);

CKINVDCx9p33_ASAP7_75t_R c1000(
.A(net1027),
.Y(net989)
);

HB1xp67_ASAP7_75t_R c1001(
.A(net117),
.Y(net990)
);

NAND2xp33_ASAP7_75t_R c1002(
.A(net978),
.B(net1043),
.Y(net991)
);

NAND2xp5_ASAP7_75t_R c1003(
.A(net1040),
.B(net986),
.Y(net992)
);

HB2xp67_ASAP7_75t_R c1004(
.A(net9752),
.Y(net993)
);

HB3xp67_ASAP7_75t_R c1005(
.A(net1018),
.Y(net994)
);

HB4xp67_ASAP7_75t_R c1006(
.A(net989),
.Y(net995)
);

SDFHx4_ASAP7_75t_R c1007(
.D(net986),
.SE(net990),
.SI(net992),
.CLK(clk),
.QN(net996)
);

INVx11_ASAP7_75t_R c1008(
.A(net943),
.Y(net997)
);

INVx13_ASAP7_75t_R c1009(
.A(net908),
.Y(net998)
);

AND3x2_ASAP7_75t_R c1010(
.A(net993),
.B(net946),
.C(net967),
.Y(net999)
);

NAND2xp67_ASAP7_75t_R c1011(
.A(net1016),
.B(net1026),
.Y(net1000)
);

NOR2x1_ASAP7_75t_R c1012(
.A(net1025),
.B(net1034),
.Y(net1001)
);

NOR2x1p5_ASAP7_75t_R c1013(
.A(net987),
.B(net1017),
.Y(net1002)
);

NOR2x2_ASAP7_75t_R c1014(
.A(net1030),
.B(net1016),
.Y(net1003)
);

INVx1_ASAP7_75t_R c1015(
.A(net1035),
.Y(net1004)
);

INVx2_ASAP7_75t_R c1016(
.A(net1026),
.Y(net1005)
);

NOR2xp33_ASAP7_75t_R c1017(
.A(net1004),
.B(in25),
.Y(net1006)
);

INVx3_ASAP7_75t_R c1018(
.A(net9650),
.Y(net1007)
);

SDFLx1_ASAP7_75t_R c1019(
.D(net990),
.SE(net130),
.SI(net921),
.CLK(clk),
.QN(net1008)
);

OAI222xp33_ASAP7_75t_R c1020(
.A1(net1007),
.A2(net1001),
.B1(net1028),
.B2(net1022),
.C1(net932),
.C2(net913),
.Y(net1009)
);

INVx4_ASAP7_75t_R c1021(
.A(net1033),
.Y(net1010)
);

ICGx4_ASAP7_75t_R c1022(
.ENA(net1028),
.SE(net1043),
.CLK(clk),
.GCLK(net1011)
);

NOR2xp67_ASAP7_75t_R c1023(
.A(net1015),
.B(net10186),
.Y(net1012)
);

OR2x2_ASAP7_75t_R c1024(
.A(net100),
.B(net955),
.Y(net1013)
);

OR2x4_ASAP7_75t_R c1025(
.A(net977),
.B(net135),
.Y(net1014)
);

OR2x6_ASAP7_75t_R c1026(
.A(net126),
.B(net51),
.Y(net1015)
);

XNOR2x1_ASAP7_75t_R c1027(
.B(net949),
.A(net122),
.Y(net1016)
);

XNOR2x2_ASAP7_75t_R c1028(
.A(net108),
.B(net945),
.Y(net1017)
);

AND3x4_ASAP7_75t_R c1029(
.A(net54),
.B(net135),
.C(net18),
.Y(net1018)
);

SDFLx2_ASAP7_75t_R c1030(
.D(net38),
.SE(net1018),
.SI(net109),
.CLK(clk),
.QN(net1019)
);

XNOR2xp5_ASAP7_75t_R c1031(
.A(net135),
.B(net133),
.Y(net1020)
);

INVx5_ASAP7_75t_R c1032(
.A(net9105),
.Y(net1021)
);

INVx6_ASAP7_75t_R c1033(
.A(net924),
.Y(net1022)
);

ICGx5_ASAP7_75t_R c1034(
.ENA(net113),
.SE(net943),
.CLK(clk),
.GCLK(net1023)
);

XOR2x1_ASAP7_75t_R c1035(
.A(net1019),
.B(net54),
.Y(net1024)
);

INVx8_ASAP7_75t_R c1036(
.A(net64),
.Y(net1025)
);

ICGx5p33DC_ASAP7_75t_R c1037(
.ENA(net1014),
.SE(net97),
.CLK(clk),
.GCLK(net1026)
);

XOR2x2_ASAP7_75t_R c1038(
.A(net945),
.B(net68),
.Y(net1027)
);

ICGx6p67DC_ASAP7_75t_R c1039(
.ENA(net902),
.SE(net130),
.CLK(clk),
.GCLK(net1028)
);

INVxp33_ASAP7_75t_R c1040(
.A(net924),
.Y(net1029)
);

INVxp67_ASAP7_75t_R c1041(
.A(net54),
.Y(net1030)
);

BUFx10_ASAP7_75t_R c1042(
.A(net1029),
.Y(net1031)
);

BUFx12_ASAP7_75t_R c1043(
.A(net1014),
.Y(net1032)
);

BUFx12f_ASAP7_75t_R c1044(
.A(net1017),
.Y(net1033)
);

XOR2xp5_ASAP7_75t_R c1045(
.A(net77),
.B(net72),
.Y(net1034)
);

BUFx16f_ASAP7_75t_R c1046(
.A(net10407),
.Y(net1035)
);

AND2x2_ASAP7_75t_R c1047(
.A(net122),
.B(net1031),
.Y(net1036)
);

AND2x4_ASAP7_75t_R c1048(
.A(net1034),
.B(net954),
.Y(net1037)
);

BUFx24_ASAP7_75t_R c1049(
.A(net962),
.Y(net1038)
);

BUFx2_ASAP7_75t_R c1050(
.A(net68),
.Y(net1039)
);

BUFx3_ASAP7_75t_R c1051(
.A(net1031),
.Y(net1040)
);

BUFx4_ASAP7_75t_R c1052(
.A(net932),
.Y(net1041)
);

BUFx4f_ASAP7_75t_R c1053(
.A(net1030),
.Y(net1042)
);

AND2x6_ASAP7_75t_R c1054(
.A(net1036),
.B(net1017),
.Y(net1043)
);

BUFx5_ASAP7_75t_R c1055(
.A(net1037),
.Y(net1044)
);

BUFx6f_ASAP7_75t_R c1056(
.A(net133),
.Y(net1045)
);

HAxp5_ASAP7_75t_R c1057(
.A(net1001),
.B(net133),
.CON(net1046)
);

ICGx8DC_ASAP7_75t_R c1058(
.ENA(net995),
.SE(net925),
.CLK(clk),
.GCLK(net1047)
);

BUFx8_ASAP7_75t_R c1059(
.A(net9105),
.Y(net1048)
);

AO21x1_ASAP7_75t_R c1060(
.A1(net1010),
.A2(net968),
.B(net1047),
.Y(net1049)
);

NAND2x1_ASAP7_75t_R c1061(
.A(net1019),
.B(net1012),
.Y(net1050)
);

NAND4xp75_ASAP7_75t_R c1062(
.A(net1011),
.B(net993),
.C(net1035),
.D(net1022),
.Y(net1051)
);

NAND2x1p5_ASAP7_75t_R c1063(
.A(net1006),
.B(net932),
.Y(net1052)
);

NAND2x2_ASAP7_75t_R c1064(
.A(net122),
.B(net9752),
.Y(net1053)
);

ICGx1_ASAP7_75t_R c1065(
.ENA(net97),
.SE(net1050),
.CLK(clk),
.GCLK(net1054)
);

NAND2xp33_ASAP7_75t_R c1066(
.A(net1047),
.B(net9744),
.Y(net1055)
);

NAND2xp5_ASAP7_75t_R c1067(
.A(net1054),
.B(net996),
.Y(net1056)
);

NOR4xp25_ASAP7_75t_R c1068(
.A(net1013),
.B(net987),
.C(net1022),
.D(net1047),
.Y(net1057)
);

NAND2xp67_ASAP7_75t_R c1069(
.A(net1047),
.B(net1057),
.Y(net1058)
);

NOR2x1_ASAP7_75t_R c1070(
.A(net1057),
.B(net1048),
.Y(net1059)
);

A2O1A1O1Ixp25_ASAP7_75t_R c1071(
.A1(net1050),
.A2(net1035),
.B(net924),
.C(net994),
.D(net1057),
.Y(net1060)
);

CKINVDCx10_ASAP7_75t_R c1072(
.A(net9864),
.Y(net1061)
);

NOR4xp75_ASAP7_75t_R c1073(
.A(net1056),
.B(net1060),
.C(net1047),
.D(net1057),
.Y(net1062)
);

NOR2x1p5_ASAP7_75t_R c1074(
.A(net130),
.B(net1061),
.Y(net1063)
);

NOR2x2_ASAP7_75t_R c1075(
.A(net1061),
.B(net1003),
.Y(net1064)
);

OAI321xp33_ASAP7_75t_R c1076(
.A1(net992),
.A2(net1054),
.A3(net1012),
.B1(net1051),
.B2(net1057),
.C(net10186),
.Y(net1065)
);

O2A1O1Ixp33_ASAP7_75t_R c1077(
.A1(net1045),
.A2(net1064),
.B(net1038),
.C(net10188),
.Y(net1066)
);

OAI33xp33_ASAP7_75t_R c1078(
.A1(net943),
.A2(net1057),
.A3(net1038),
.B1(net9752),
.B2(net10188),
.B3(net10189),
.Y(net1067)
);

CKINVDCx11_ASAP7_75t_R c1079(
.A(net9200),
.Y(net1068)
);

CKINVDCx12_ASAP7_75t_R c1080(
.A(net9185),
.Y(net1069)
);

CKINVDCx14_ASAP7_75t_R c1081(
.A(net147),
.Y(net1070)
);

CKINVDCx16_ASAP7_75t_R c1082(
.A(net178),
.Y(net1071)
);

CKINVDCx20_ASAP7_75t_R c1083(
.A(net9185),
.Y(net1072)
);

CKINVDCx5p33_ASAP7_75t_R c1084(
.A(net1055),
.Y(net1073)
);

NOR2xp33_ASAP7_75t_R c1085(
.A(in25),
.B(net61),
.Y(net1074)
);

CKINVDCx6p67_ASAP7_75t_R c1086(
.A(net185),
.Y(net1075)
);

CKINVDCx8_ASAP7_75t_R c1087(
.A(net91),
.Y(net1076)
);

NOR2xp67_ASAP7_75t_R c1088(
.A(net1047),
.B(net1074),
.Y(net1077)
);

CKINVDCx9p33_ASAP7_75t_R c1089(
.A(net1005),
.Y(net1078)
);

HB1xp67_ASAP7_75t_R c1090(
.A(net981),
.Y(net1079)
);

HB2xp67_ASAP7_75t_R c1091(
.A(net1036),
.Y(net1080)
);

HB3xp67_ASAP7_75t_R c1092(
.A(net170),
.Y(net1081)
);

AO21x2_ASAP7_75t_R c1093(
.A1(net1081),
.A2(net946),
.B(net1071),
.Y(net1082)
);

HB4xp67_ASAP7_75t_R c1094(
.A(net1021),
.Y(net1083)
);

INVx11_ASAP7_75t_R c1095(
.A(net9200),
.Y(net1084)
);

INVx13_ASAP7_75t_R c1096(
.A(net1000),
.Y(net1085)
);

INVx1_ASAP7_75t_R c1097(
.A(net921),
.Y(net1086)
);

INVx2_ASAP7_75t_R c1098(
.A(net215),
.Y(net1087)
);

INVx3_ASAP7_75t_R c1099(
.A(net1002),
.Y(net1088)
);

INVx4_ASAP7_75t_R c1100(
.A(net210),
.Y(net1089)
);

INVx5_ASAP7_75t_R c1101(
.A(net1072),
.Y(net1090)
);

INVx6_ASAP7_75t_R c1102(
.A(net1070),
.Y(net1091)
);

INVx8_ASAP7_75t_R c1103(
.A(net10496),
.Y(net1092)
);

OR2x2_ASAP7_75t_R c1104(
.A(net1075),
.B(net10188),
.Y(net1093)
);

INVxp33_ASAP7_75t_R c1105(
.A(net9221),
.Y(net1094)
);

INVxp67_ASAP7_75t_R c1106(
.A(net9828),
.Y(net1095)
);

BUFx10_ASAP7_75t_R c1107(
.A(net9291),
.Y(net1096)
);

OR2x4_ASAP7_75t_R c1108(
.A(net1084),
.B(net1093),
.Y(net1097)
);

BUFx12_ASAP7_75t_R c1109(
.A(net946),
.Y(net1098)
);

SDFLx3_ASAP7_75t_R c1110(
.D(net220),
.SE(net191),
.SI(net902),
.CLK(clk),
.QN(net1099)
);

OR2x6_ASAP7_75t_R c1111(
.A(net111),
.B(net1021),
.Y(net1100)
);

XNOR2x1_ASAP7_75t_R c1112(
.B(net1097),
.A(net1085),
.Y(net1101)
);

AOI21x1_ASAP7_75t_R c1113(
.A1(net1000),
.A2(net1093),
.B(net10188),
.Y(net1102)
);

BUFx12f_ASAP7_75t_R c1114(
.A(net193),
.Y(net1103)
);

XNOR2x2_ASAP7_75t_R c1115(
.A(net1074),
.B(net1096),
.Y(net1104)
);

BUFx16f_ASAP7_75t_R c1116(
.A(net9825),
.Y(net1105)
);

BUFx24_ASAP7_75t_R c1117(
.A(net156),
.Y(net1106)
);

SDFLx4_ASAP7_75t_R c1118(
.D(net1106),
.SE(net1101),
.SI(net1085),
.CLK(clk),
.QN(net1107)
);

XNOR2xp5_ASAP7_75t_R c1119(
.A(net1039),
.B(net1085),
.Y(net1108)
);

XOR2x1_ASAP7_75t_R c1120(
.A(net151),
.B(net1081),
.Y(net1109)
);

AOI21xp33_ASAP7_75t_R c1121(
.A1(net108),
.A2(net1107),
.B(net1051),
.Y(net1110)
);

BUFx2_ASAP7_75t_R c1122(
.A(net156),
.Y(net1111)
);

XOR2x2_ASAP7_75t_R c1123(
.A(net185),
.B(net91),
.Y(net1112)
);

ICGx2_ASAP7_75t_R c1124(
.ENA(net218),
.SE(net1108),
.CLK(clk),
.GCLK(net1113)
);

XOR2xp5_ASAP7_75t_R c1125(
.A(net1070),
.B(net1075),
.Y(net1114)
);

BUFx3_ASAP7_75t_R c1126(
.A(net111),
.Y(net1115)
);

AND2x2_ASAP7_75t_R c1127(
.A(net70),
.B(net1107),
.Y(net1116)
);

AND2x4_ASAP7_75t_R c1128(
.A(net1103),
.B(net1110),
.Y(net1117)
);

BUFx4_ASAP7_75t_R c1129(
.A(net1115),
.Y(net1118)
);

AOI21xp5_ASAP7_75t_R c1130(
.A1(net1044),
.A2(net965),
.B(net10188),
.Y(net1119)
);

FAx1_ASAP7_75t_R c1131(
.A(net1098),
.B(net1112),
.CI(net1083),
.SN(net1120)
);

AND2x6_ASAP7_75t_R c1132(
.A(net184),
.B(net210),
.Y(net1121)
);

BUFx4f_ASAP7_75t_R c1133(
.A(net9953),
.Y(net1122)
);

HAxp5_ASAP7_75t_R c1134(
.A(net1095),
.B(net218),
.CON(net1124),
.SN(net1123)
);

NAND2x1_ASAP7_75t_R c1135(
.A(net1124),
.B(net1112),
.Y(net1125)
);

NAND2x1p5_ASAP7_75t_R c1136(
.A(net191),
.B(net1051),
.Y(net1126)
);

BUFx5_ASAP7_75t_R c1137(
.A(net1091),
.Y(net1127)
);

MAJIxp5_ASAP7_75t_R c1138(
.A(net1079),
.B(net1127),
.C(net88),
.Y(net1128)
);

NAND2x2_ASAP7_75t_R c1139(
.A(net61),
.B(net1104),
.Y(net1129)
);

NAND2xp33_ASAP7_75t_R c1140(
.A(net1094),
.B(net1121),
.Y(net1130)
);

MAJx2_ASAP7_75t_R c1141(
.A(net1073),
.B(net1078),
.C(net981),
.Y(net1131)
);

NAND2xp5_ASAP7_75t_R c1142(
.A(net1071),
.B(net1129),
.Y(net1132)
);

MAJx3_ASAP7_75t_R c1143(
.A(net1084),
.B(net1121),
.C(net108),
.Y(net1133)
);

DFFASRHQNx1_ASAP7_75t_R c1144(
.D(net1117),
.RESETN(net1127),
.SETN(net1128),
.CLK(clk),
.QN(net1134)
);

NAND3x1_ASAP7_75t_R c1145(
.A(net1133),
.B(net1123),
.C(net1132),
.Y(net1135)
);

NAND2xp67_ASAP7_75t_R c1146(
.A(net1129),
.B(net1122),
.Y(net1136)
);

BUFx6f_ASAP7_75t_R c1147(
.A(net1118),
.Y(net1137)
);

NAND3x2_ASAP7_75t_R c1148(
.B(net172),
.C(net1093),
.A(net1128),
.Y(net1138)
);

NOR2x1_ASAP7_75t_R c1149(
.A(net1104),
.B(net1092),
.Y(net1139)
);

NAND3xp33_ASAP7_75t_R c1150(
.A(net1137),
.B(net215),
.C(net1139),
.Y(net1140)
);

AND5x1_ASAP7_75t_R c1151(
.A(net1119),
.B(net1130),
.C(net1128),
.D(net913),
.E(net1140),
.Y(net1141)
);

NOR3x1_ASAP7_75t_R c1152(
.A(net1128),
.B(net1086),
.C(net1113),
.Y(net1142)
);

NOR3x2_ASAP7_75t_R c1153(
.B(net1130),
.C(net1140),
.A(net1079),
.Y(net1143)
);

NOR3xp33_ASAP7_75t_R c1154(
.A(net1113),
.B(net1140),
.C(net9992),
.Y(net1144)
);

NOR2x1p5_ASAP7_75t_R c1155(
.A(net186),
.B(net9992),
.Y(net1145)
);

NOR2x2_ASAP7_75t_R c1156(
.A(net1139),
.B(net1138),
.Y(net1146)
);

ICGx2p67DC_ASAP7_75t_R c1157(
.ENA(net1146),
.SE(net184),
.CLK(clk),
.GCLK(net1147)
);

SDFHx1_ASAP7_75t_R c1158(
.D(net1145),
.SE(net1140),
.SI(net1146),
.CLK(clk),
.QN(net1148)
);

OA21x2_ASAP7_75t_R c1159(
.A1(net1096),
.A2(net1137),
.B(net1073),
.Y(net1149)
);

OAI21x1_ASAP7_75t_R c1160(
.A1(net1116),
.A2(net1142),
.B(net1136),
.Y(net1150)
);

AO222x2_ASAP7_75t_R c1161(
.A1(net907),
.A2(net1150),
.B1(net1140),
.B2(net1047),
.C1(net1021),
.C2(net9746),
.Y(net1151)
);

BUFx8_ASAP7_75t_R c1162(
.A(net9238),
.Y(net1152)
);

CKINVDCx10_ASAP7_75t_R c1163(
.A(net253),
.Y(net1153)
);

CKINVDCx11_ASAP7_75t_R c1164(
.A(net241),
.Y(net1154)
);

CKINVDCx12_ASAP7_75t_R c1165(
.A(net1086),
.Y(net1155)
);

CKINVDCx14_ASAP7_75t_R c1166(
.A(net965),
.Y(net1156)
);

CKINVDCx16_ASAP7_75t_R c1167(
.A(net9969),
.Y(net1157)
);

CKINVDCx20_ASAP7_75t_R c1168(
.A(net9969),
.Y(net1158)
);

CKINVDCx5p33_ASAP7_75t_R c1169(
.A(net1155),
.Y(net1159)
);

CKINVDCx6p67_ASAP7_75t_R c1170(
.A(net1159),
.Y(net1160)
);

CKINVDCx8_ASAP7_75t_R c1171(
.A(net10095),
.Y(net1161)
);

CKINVDCx9p33_ASAP7_75t_R c1172(
.A(net1142),
.Y(net1162)
);

NOR2xp33_ASAP7_75t_R c1173(
.A(net202),
.B(net1132),
.Y(net1163)
);

HB1xp67_ASAP7_75t_R c1174(
.A(net253),
.Y(net1164)
);

HB2xp67_ASAP7_75t_R c1175(
.A(net10427),
.Y(net1165)
);

HB3xp67_ASAP7_75t_R c1176(
.A(net997),
.Y(net1166)
);

HB4xp67_ASAP7_75t_R c1177(
.A(net10522),
.Y(net1167)
);

NOR2xp67_ASAP7_75t_R c1178(
.A(net1051),
.B(net1038),
.Y(net1168)
);

OR2x2_ASAP7_75t_R c1179(
.A(net1162),
.B(net1140),
.Y(net1169)
);

OR2x4_ASAP7_75t_R c1180(
.A(net1112),
.B(net228),
.Y(net1170)
);

OR2x6_ASAP7_75t_R c1181(
.A(net997),
.B(net1153),
.Y(net1171)
);

INVx11_ASAP7_75t_R c1182(
.A(net1099),
.Y(net1172)
);

INVx13_ASAP7_75t_R c1183(
.A(net10427),
.Y(net1173)
);

INVx1_ASAP7_75t_R c1184(
.A(net242),
.Y(net1174)
);

INVx2_ASAP7_75t_R c1185(
.A(net9650),
.Y(net1175)
);

OAI21xp33_ASAP7_75t_R c1186(
.A1(net1133),
.A2(net1101),
.B(net1171),
.Y(net1176)
);

INVx3_ASAP7_75t_R c1187(
.A(net1077),
.Y(net1177)
);

INVx4_ASAP7_75t_R c1188(
.A(net1165),
.Y(net1178)
);

XNOR2x1_ASAP7_75t_R c1189(
.B(net1100),
.A(net1157),
.Y(net1179)
);

OAI21xp5_ASAP7_75t_R c1190(
.A1(net186),
.A2(net1023),
.B(net1069),
.Y(net1180)
);

XNOR2x2_ASAP7_75t_R c1191(
.A(net307),
.B(net1156),
.Y(net1181)
);

INVx5_ASAP7_75t_R c1192(
.A(net1175),
.Y(net1182)
);

INVx6_ASAP7_75t_R c1193(
.A(net1175),
.Y(net1183)
);

INVx8_ASAP7_75t_R c1194(
.A(net1174),
.Y(net1184)
);

XNOR2xp5_ASAP7_75t_R c1195(
.A(net1023),
.B(net59),
.Y(net1185)
);

XOR2x1_ASAP7_75t_R c1196(
.A(net1158),
.B(net1167),
.Y(net1186)
);

XOR2x2_ASAP7_75t_R c1197(
.A(net1177),
.B(net1186),
.Y(net1187)
);

INVxp33_ASAP7_75t_R c1198(
.A(net1082),
.Y(net1188)
);

INVxp67_ASAP7_75t_R c1199(
.A(net1081),
.Y(net1189)
);

XOR2xp5_ASAP7_75t_R c1200(
.A(net1152),
.B(net9993),
.Y(net1190)
);

AND2x2_ASAP7_75t_R c1201(
.A(net1127),
.B(net1186),
.Y(net1191)
);

BUFx10_ASAP7_75t_R c1202(
.A(net1188),
.Y(net1192)
);

ICGx3_ASAP7_75t_R c1203(
.ENA(net1101),
.SE(net299),
.CLK(clk),
.GCLK(net1193)
);

BUFx12_ASAP7_75t_R c1204(
.A(net9221),
.Y(net1194)
);

BUFx12f_ASAP7_75t_R c1205(
.A(net1193),
.Y(net1195)
);

BUFx16f_ASAP7_75t_R c1206(
.A(net1166),
.Y(net1196)
);

AND2x4_ASAP7_75t_R c1207(
.A(net902),
.B(net1186),
.Y(net1197)
);

OR3x1_ASAP7_75t_R c1208(
.A(net1192),
.B(net1171),
.C(net1173),
.Y(net1198)
);

OR3x2_ASAP7_75t_R c1209(
.A(net228),
.B(net1198),
.C(net1153),
.Y(net1199)
);

BUFx24_ASAP7_75t_R c1210(
.A(net1189),
.Y(net1200)
);

AND2x6_ASAP7_75t_R c1211(
.A(net1185),
.B(net1158),
.Y(net1201)
);

BUFx2_ASAP7_75t_R c1212(
.A(net1178),
.Y(net1202)
);

O2A1O1Ixp5_ASAP7_75t_R c1213(
.A1(net1121),
.A2(net297),
.B(net47),
.C(net1038),
.Y(net1203)
);

HAxp5_ASAP7_75t_R c1214(
.A(net1068),
.B(net1189),
.CON(net1204)
);

NAND2x1_ASAP7_75t_R c1215(
.A(net1191),
.B(net1197),
.Y(net1205)
);

BUFx3_ASAP7_75t_R c1216(
.A(net10006),
.Y(net1206)
);

NAND2x1p5_ASAP7_75t_R c1217(
.A(net1186),
.B(net1200),
.Y(net1207)
);

BUFx4_ASAP7_75t_R c1218(
.A(net1203),
.Y(net1208)
);

NAND2x2_ASAP7_75t_R c1219(
.A(net1162),
.B(net1191),
.Y(net1209)
);

NAND2xp33_ASAP7_75t_R c1220(
.A(net1180),
.B(net1177),
.Y(net1210)
);

NAND2xp5_ASAP7_75t_R c1221(
.A(net1200),
.B(net1186),
.Y(net1211)
);

BUFx4f_ASAP7_75t_R c1222(
.A(net10430),
.Y(net1212)
);

NAND2xp67_ASAP7_75t_R c1223(
.A(net1174),
.B(net1197),
.Y(net1213)
);

NOR2x1_ASAP7_75t_R c1224(
.A(net1187),
.B(net1188),
.Y(net1214)
);

OR3x4_ASAP7_75t_R c1225(
.A(net1087),
.B(net297),
.C(net1214),
.Y(net1215)
);

AND3x1_ASAP7_75t_R c1226(
.A(net297),
.B(net1207),
.C(net1185),
.Y(net1216)
);

NOR2x1p5_ASAP7_75t_R c1227(
.A(net1154),
.B(net1178),
.Y(net1217)
);

NOR2x2_ASAP7_75t_R c1228(
.A(net1210),
.B(net965),
.Y(net1218)
);

NOR2xp33_ASAP7_75t_R c1229(
.A(net1216),
.B(net9652),
.Y(net1219)
);

NOR2xp67_ASAP7_75t_R c1230(
.A(net1215),
.B(net1171),
.Y(net1220)
);

OR2x2_ASAP7_75t_R c1231(
.A(net18),
.B(net1187),
.Y(net1221)
);

AND3x2_ASAP7_75t_R c1232(
.A(net1206),
.B(net1219),
.C(net1211),
.Y(net1222)
);

OR2x4_ASAP7_75t_R c1233(
.A(net240),
.B(net1189),
.Y(net1223)
);

AND3x4_ASAP7_75t_R c1234(
.A(net1218),
.B(net1193),
.C(net1167),
.Y(net1224)
);

SDFHx2_ASAP7_75t_R c1235(
.D(net1198),
.SE(net1174),
.SI(net1162),
.CLK(clk),
.QN(net1225)
);

AO21x1_ASAP7_75t_R c1236(
.A1(net1223),
.A2(net1210),
.B(net1224),
.Y(net1226)
);

AO21x2_ASAP7_75t_R c1237(
.A1(net1182),
.A2(net1085),
.B(net10006),
.Y(net1227)
);

AOI21x1_ASAP7_75t_R c1238(
.A1(net1207),
.A2(net1201),
.B(net1175),
.Y(net1228)
);

AO33x2_ASAP7_75t_R c1239(
.A1(net1206),
.A2(net1051),
.A3(net1160),
.B1(net1190),
.B2(net245),
.B3(net10108),
.Y(net1229)
);

OA211x2_ASAP7_75t_R c1240(
.A1(net1201),
.A2(net1210),
.B(net1112),
.C(net1155),
.Y(net1230)
);

OA22x2_ASAP7_75t_R c1241(
.A1(net1228),
.A2(net1198),
.B1(net1224),
.B2(net1193),
.Y(net1231)
);

AOI222xp33_ASAP7_75t_R c1242(
.A1(net288),
.A2(net1202),
.B1(net240),
.B2(net1193),
.C1(net1155),
.C2(net245),
.Y(net1232)
);

OR2x6_ASAP7_75t_R c1243(
.A(net1213),
.B(net1230),
.Y(net1233)
);

XNOR2x1_ASAP7_75t_R c1244(
.B(net1216),
.A(net1223),
.Y(net1234)
);

BUFx5_ASAP7_75t_R c1245(
.A(net9963),
.Y(net1235)
);

BUFx6f_ASAP7_75t_R c1246(
.A(net319),
.Y(net1236)
);

BUFx8_ASAP7_75t_R c1247(
.A(net1125),
.Y(net1237)
);

CKINVDCx10_ASAP7_75t_R c1248(
.A(net9652),
.Y(net1238)
);

XNOR2x2_ASAP7_75t_R c1249(
.A(net290),
.B(net1109),
.Y(net1239)
);

CKINVDCx11_ASAP7_75t_R c1250(
.A(net1171),
.Y(net1240)
);

CKINVDCx12_ASAP7_75t_R c1251(
.A(net1069),
.Y(net1241)
);

CKINVDCx14_ASAP7_75t_R c1252(
.A(net10126),
.Y(net1242)
);

XNOR2xp5_ASAP7_75t_R c1253(
.A(net1238),
.B(net9828),
.Y(net1243)
);

CKINVDCx16_ASAP7_75t_R c1254(
.A(net9131),
.Y(net1244)
);

CKINVDCx20_ASAP7_75t_R c1255(
.A(net9963),
.Y(net1245)
);

CKINVDCx5p33_ASAP7_75t_R c1256(
.A(net1240),
.Y(net1246)
);

XOR2x1_ASAP7_75t_R c1257(
.A(net174),
.B(net389),
.Y(net1247)
);

CKINVDCx6p67_ASAP7_75t_R c1258(
.A(net9131),
.Y(net1248)
);

CKINVDCx8_ASAP7_75t_R c1259(
.A(net1244),
.Y(net1249)
);

CKINVDCx9p33_ASAP7_75t_R c1260(
.A(net1200),
.Y(net1250)
);

XOR2x2_ASAP7_75t_R c1261(
.A(net47),
.B(net1219),
.Y(net1251)
);

ICGx4DC_ASAP7_75t_R c1262(
.ENA(net384),
.SE(net1138),
.CLK(clk),
.GCLK(net1252)
);

AOI21xp33_ASAP7_75t_R c1263(
.A1(net1202),
.A2(net1160),
.B(net9896),
.Y(net1253)
);

HB1xp67_ASAP7_75t_R c1264(
.A(net1085),
.Y(net1254)
);

HB2xp67_ASAP7_75t_R c1265(
.A(net304),
.Y(net1255)
);

HB3xp67_ASAP7_75t_R c1266(
.A(net1242),
.Y(net1256)
);

HB4xp67_ASAP7_75t_R c1267(
.A(net1086),
.Y(net1257)
);

INVx11_ASAP7_75t_R c1268(
.A(net1241),
.Y(net1258)
);

AND5x2_ASAP7_75t_R c1269(
.A(net216),
.B(net1257),
.C(net1155),
.D(net1038),
.E(net1190),
.Y(net1259)
);

INVx13_ASAP7_75t_R c1270(
.A(net256),
.Y(net1260)
);

INVx1_ASAP7_75t_R c1271(
.A(net1202),
.Y(net1261)
);

XOR2xp5_ASAP7_75t_R c1272(
.A(net1152),
.B(net1167),
.Y(net1262)
);

INVx2_ASAP7_75t_R c1273(
.A(net1105),
.Y(net1263)
);

INVx3_ASAP7_75t_R c1274(
.A(net1109),
.Y(net1264)
);

INVx4_ASAP7_75t_R c1275(
.A(net9261),
.Y(net1265)
);

AND2x2_ASAP7_75t_R c1276(
.A(net1160),
.B(net9993),
.Y(net1266)
);

INVx5_ASAP7_75t_R c1277(
.A(net370),
.Y(net1267)
);

INVx6_ASAP7_75t_R c1278(
.A(net1126),
.Y(net1268)
);

INVx8_ASAP7_75t_R c1279(
.A(net1249),
.Y(net1269)
);

INVxp33_ASAP7_75t_R c1280(
.A(net1262),
.Y(net1270)
);

OA31x2_ASAP7_75t_R c1281(
.A1(net1236),
.A2(net1227),
.A3(net1244),
.B1(net389),
.Y(net1271)
);

INVxp67_ASAP7_75t_R c1282(
.A(net1263),
.Y(net1272)
);

BUFx10_ASAP7_75t_R c1283(
.A(net1270),
.Y(net1273)
);

AND2x4_ASAP7_75t_R c1284(
.A(net276),
.B(net10191),
.Y(net1274)
);

BUFx12_ASAP7_75t_R c1285(
.A(net1243),
.Y(net1275)
);

AOI21xp5_ASAP7_75t_R c1286(
.A1(net1268),
.A2(net1171),
.B(net1257),
.Y(net1276)
);

BUFx12f_ASAP7_75t_R c1287(
.A(net1260),
.Y(net1277)
);

BUFx16f_ASAP7_75t_R c1288(
.A(net9946),
.Y(net1278)
);

BUFx24_ASAP7_75t_R c1289(
.A(net9248),
.Y(net1279)
);

BUFx2_ASAP7_75t_R c1290(
.A(net10006),
.Y(net1280)
);

OAI211xp5_ASAP7_75t_R c1291(
.A1(net311),
.A2(net1257),
.B(net1238),
.C(net9828),
.Y(net1281)
);

AND2x6_ASAP7_75t_R c1292(
.A(net1274),
.B(net1280),
.Y(net1282)
);

BUFx3_ASAP7_75t_R c1293(
.A(net10095),
.Y(net1283)
);

BUFx4_ASAP7_75t_R c1294(
.A(net1261),
.Y(net1284)
);

BUFx4f_ASAP7_75t_R c1295(
.A(net1284),
.Y(net1285)
);

HAxp5_ASAP7_75t_R c1296(
.A(net1246),
.B(net1168),
.CON(net1286)
);

BUFx5_ASAP7_75t_R c1297(
.A(net9261),
.Y(net1287)
);

NAND2x1_ASAP7_75t_R c1298(
.A(net1269),
.B(net1270),
.Y(net1288)
);

NAND2x1p5_ASAP7_75t_R c1299(
.A(net1288),
.B(net1263),
.Y(net1289)
);

BUFx6f_ASAP7_75t_R c1300(
.A(net9889),
.Y(net1290)
);

NAND2x2_ASAP7_75t_R c1301(
.A(net318),
.B(net1282),
.Y(net1291)
);

BUFx8_ASAP7_75t_R c1302(
.A(net375),
.Y(net1292)
);

FAx1_ASAP7_75t_R c1303(
.A(net358),
.B(net1263),
.CI(net9946),
.SN(net1294),
.CON(net1293)
);

NAND2xp33_ASAP7_75t_R c1304(
.A(net1113),
.B(net1288),
.Y(net1295)
);

NAND2xp5_ASAP7_75t_R c1305(
.A(net1237),
.B(net1290),
.Y(net1296)
);

NAND2xp67_ASAP7_75t_R c1306(
.A(net1291),
.B(net1155),
.Y(net1297)
);

NOR2x1_ASAP7_75t_R c1307(
.A(net1255),
.B(net1279),
.Y(net1298)
);

CKINVDCx10_ASAP7_75t_R c1308(
.A(net1296),
.Y(net1299)
);

OAI22x1_ASAP7_75t_R c1309(
.A1(net1253),
.A2(net389),
.B1(net394),
.B2(net1190),
.Y(net1300)
);

CKINVDCx11_ASAP7_75t_R c1310(
.A(net1281),
.Y(net1301)
);

CKINVDCx12_ASAP7_75t_R c1311(
.A(net10038),
.Y(net1302)
);

NOR2x1p5_ASAP7_75t_R c1312(
.A(net351),
.B(net1125),
.Y(net1303)
);

NOR2x2_ASAP7_75t_R c1313(
.A(net1161),
.B(net1290),
.Y(net1304)
);

MAJIxp5_ASAP7_75t_R c1314(
.A(net1302),
.B(net1298),
.C(net958),
.Y(net1305)
);

NOR2xp33_ASAP7_75t_R c1315(
.A(net1285),
.B(net1252),
.Y(net1306)
);

CKINVDCx14_ASAP7_75t_R c1316(
.A(net9954),
.Y(net1307)
);

OAI22xp33_ASAP7_75t_R c1317(
.A1(net1306),
.A2(net1263),
.B1(net1282),
.B2(net9832),
.Y(net1308)
);

MAJx2_ASAP7_75t_R c1318(
.A(net1265),
.B(net1249),
.C(net1269),
.Y(net1309)
);

OAI22xp5_ASAP7_75t_R c1319(
.A1(net1208),
.A2(net1155),
.B1(net331),
.B2(net1290),
.Y(net1310)
);

NOR2xp67_ASAP7_75t_R c1320(
.A(net10051),
.B(net10191),
.Y(net1311)
);

MAJx3_ASAP7_75t_R c1321(
.A(net1307),
.B(net1308),
.C(net10051),
.Y(net1312)
);

OR2x2_ASAP7_75t_R c1322(
.A(net1301),
.B(net1312),
.Y(net1313)
);

NAND3x1_ASAP7_75t_R c1323(
.A(net1225),
.B(net1269),
.C(net9832),
.Y(net1314)
);

AO221x1_ASAP7_75t_R c1324(
.A1(net1297),
.A2(net1298),
.B1(net1290),
.B2(net1313),
.C(net1292),
.Y(net1315)
);

SDFHx3_ASAP7_75t_R c1325(
.D(net1164),
.SE(net1208),
.SI(net1259),
.CLK(clk),
.QN(net1316)
);

OR2x4_ASAP7_75t_R c1326(
.A(net1309),
.B(net1293),
.Y(net1317)
);

NAND3x2_ASAP7_75t_R c1327(
.B(net1315),
.C(net1316),
.A(net1317),
.Y(net1318)
);

CKINVDCx16_ASAP7_75t_R c1328(
.A(net9239),
.Y(net1319)
);

CKINVDCx20_ASAP7_75t_R c1329(
.A(net1311),
.Y(net1320)
);

OR2x6_ASAP7_75t_R c1330(
.A(net295),
.B(net402),
.Y(net1321)
);

CKINVDCx5p33_ASAP7_75t_R c1331(
.A(net10035),
.Y(net1322)
);

XNOR2x1_ASAP7_75t_R c1332(
.B(net1225),
.A(net1219),
.Y(net1323)
);

CKINVDCx6p67_ASAP7_75t_R c1333(
.A(net1097),
.Y(net1324)
);

XNOR2x2_ASAP7_75t_R c1334(
.A(net157),
.B(net1292),
.Y(net1325)
);

SDFHx4_ASAP7_75t_R c1335(
.D(net293),
.SE(net1168),
.SI(net1254),
.CLK(clk),
.QN(net1326)
);

XNOR2xp5_ASAP7_75t_R c1336(
.A(net145),
.B(net429),
.Y(net1327)
);

CKINVDCx8_ASAP7_75t_R c1337(
.A(net421),
.Y(net1328)
);

XOR2x1_ASAP7_75t_R c1338(
.A(net402),
.B(net10177),
.Y(net1329)
);

XOR2x2_ASAP7_75t_R c1339(
.A(net1327),
.B(net1257),
.Y(net1330)
);

CKINVDCx9p33_ASAP7_75t_R c1340(
.A(net477),
.Y(net1331)
);

XOR2xp5_ASAP7_75t_R c1341(
.A(net1170),
.B(net1316),
.Y(net1332)
);

OAI31xp33_ASAP7_75t_R c1342(
.A1(net410),
.A2(net1332),
.A3(net1275),
.B(net1312),
.Y(net1333)
);

HB1xp67_ASAP7_75t_R c1343(
.A(net1219),
.Y(net1334)
);

NAND3xp33_ASAP7_75t_R c1344(
.A(net1235),
.B(net428),
.C(net10192),
.Y(net1335)
);

HB2xp67_ASAP7_75t_R c1345(
.A(net418),
.Y(net1336)
);

HB3xp67_ASAP7_75t_R c1346(
.A(net435),
.Y(net1337)
);

AND2x2_ASAP7_75t_R c1347(
.A(net1180),
.B(net1279),
.Y(net1338)
);

AND2x4_ASAP7_75t_R c1348(
.A(net1217),
.B(net458),
.Y(net1339)
);

HB4xp67_ASAP7_75t_R c1349(
.A(net331),
.Y(net1340)
);

ICGx4_ASAP7_75t_R c1350(
.ENA(net1254),
.SE(net462),
.CLK(clk),
.GCLK(net1341)
);

INVx11_ASAP7_75t_R c1351(
.A(net10570),
.Y(net1342)
);

INVx13_ASAP7_75t_R c1352(
.A(net1245),
.Y(net1343)
);

INVx1_ASAP7_75t_R c1353(
.A(net10045),
.Y(net1344)
);

INVx2_ASAP7_75t_R c1354(
.A(net1332),
.Y(net1345)
);

AND2x6_ASAP7_75t_R c1355(
.A(net1225),
.B(net9904),
.Y(net1346)
);

INVx3_ASAP7_75t_R c1356(
.A(net1343),
.Y(net1347)
);

INVx4_ASAP7_75t_R c1357(
.A(net1283),
.Y(net1348)
);

INVx5_ASAP7_75t_R c1358(
.A(net393),
.Y(net1349)
);

HAxp5_ASAP7_75t_R c1359(
.A(net409),
.B(net1339),
.CON(net1351),
.SN(net1350)
);

INVx6_ASAP7_75t_R c1360(
.A(net1329),
.Y(net1352)
);

NAND2x1_ASAP7_75t_R c1361(
.A(net1252),
.B(net1303),
.Y(net1353)
);

NAND2x1p5_ASAP7_75t_R c1362(
.A(net439),
.B(net1348),
.Y(net1354)
);

NAND2x2_ASAP7_75t_R c1363(
.A(net466),
.B(net1350),
.Y(net1355)
);

NAND2xp33_ASAP7_75t_R c1364(
.A(net413),
.B(net10192),
.Y(net1356)
);

INVx8_ASAP7_75t_R c1365(
.A(net9933),
.Y(net1357)
);

INVxp33_ASAP7_75t_R c1366(
.A(net272),
.Y(net1358)
);

INVxp67_ASAP7_75t_R c1367(
.A(net1357),
.Y(net1359)
);

OAI31xp67_ASAP7_75t_R c1368(
.A1(net1359),
.A2(net1337),
.A3(net441),
.B(net1038),
.Y(net1360)
);

NOR3x1_ASAP7_75t_R c1369(
.A(net1319),
.B(net1331),
.C(net1341),
.Y(net1361)
);

BUFx10_ASAP7_75t_R c1370(
.A(net10071),
.Y(net1362)
);

NAND2xp5_ASAP7_75t_R c1371(
.A(net458),
.B(net1344),
.Y(net1363)
);

NAND2xp67_ASAP7_75t_R c1372(
.A(net1279),
.B(net421),
.Y(net1364)
);

BUFx12_ASAP7_75t_R c1373(
.A(net1295),
.Y(net1365)
);

BUFx12f_ASAP7_75t_R c1374(
.A(net1361),
.Y(net1366)
);

NOR2x1_ASAP7_75t_R c1375(
.A(net1324),
.B(net10192),
.Y(net1367)
);

NOR3x2_ASAP7_75t_R c1376(
.B(net1322),
.C(net1242),
.A(net1338),
.Y(net1368)
);

NOR2x1p5_ASAP7_75t_R c1377(
.A(net1353),
.B(net413),
.Y(net1369)
);

NOR2x2_ASAP7_75t_R c1378(
.A(net1366),
.B(net410),
.Y(net1370)
);

BUFx16f_ASAP7_75t_R c1379(
.A(net1242),
.Y(net1371)
);

BUFx24_ASAP7_75t_R c1380(
.A(net10045),
.Y(net1372)
);

BUFx2_ASAP7_75t_R c1381(
.A(net1333),
.Y(net1373)
);

BUFx3_ASAP7_75t_R c1382(
.A(net1362),
.Y(net1374)
);

AO221x2_ASAP7_75t_R c1383(
.A1(net1334),
.A2(net1343),
.B1(net1357),
.B2(net1168),
.C(net1348),
.Y(net1375)
);

NOR3xp33_ASAP7_75t_R c1384(
.A(net1316),
.B(net1345),
.C(net10193),
.Y(net1376)
);

OR4x1_ASAP7_75t_R c1385(
.A(net1376),
.B(net1346),
.C(net1365),
.D(net1336),
.Y(net1377)
);

SDFLx1_ASAP7_75t_R c1386(
.D(net1361),
.SE(net436),
.SI(net9832),
.CLK(clk),
.QN(net1378)
);

BUFx4_ASAP7_75t_R c1387(
.A(net10499),
.Y(net1379)
);

NOR2xp33_ASAP7_75t_R c1388(
.A(net1344),
.B(net1341),
.Y(net1380)
);

BUFx4f_ASAP7_75t_R c1389(
.A(net10390),
.Y(net1381)
);

BUFx5_ASAP7_75t_R c1390(
.A(net10409),
.Y(net1382)
);

NOR2xp67_ASAP7_75t_R c1391(
.A(net1382),
.B(net1365),
.Y(net1383)
);

OR2x2_ASAP7_75t_R c1392(
.A(net1380),
.B(net1292),
.Y(net1384)
);

OA21x2_ASAP7_75t_R c1393(
.A1(net1354),
.A2(net1312),
.B(net1378),
.Y(net1385)
);

OR2x4_ASAP7_75t_R c1394(
.A(net1379),
.B(net10065),
.Y(net1386)
);

OR2x6_ASAP7_75t_R c1395(
.A(net1372),
.B(net466),
.Y(net1387)
);

XNOR2x1_ASAP7_75t_R c1396(
.B(net1385),
.A(net1225),
.Y(net1388)
);

XNOR2x2_ASAP7_75t_R c1397(
.A(net1387),
.B(net1313),
.Y(net1389)
);

XNOR2xp5_ASAP7_75t_R c1398(
.A(net1370),
.B(net1344),
.Y(net1390)
);

XOR2x1_ASAP7_75t_R c1399(
.A(net1374),
.B(net1368),
.Y(net1391)
);

OAI21x1_ASAP7_75t_R c1400(
.A1(net1311),
.A2(net10065),
.B(net10193),
.Y(net1392)
);

BUFx6f_ASAP7_75t_R c1401(
.A(net10035),
.Y(net1393)
);

AO32x1_ASAP7_75t_R c1402(
.A1(net1392),
.A2(net1364),
.A3(net1347),
.B1(net331),
.B2(net1324),
.Y(net1394)
);

AO32x2_ASAP7_75t_R c1403(
.A1(net1384),
.A2(net1379),
.A3(net1304),
.B1(net1348),
.B2(net1365),
.Y(net1395)
);

OR4x2_ASAP7_75t_R c1404(
.A(net1275),
.B(net1388),
.C(net1376),
.D(net1338),
.Y(net1396)
);

A2O1A1Ixp33_ASAP7_75t_R c1405(
.A1(net1356),
.A2(net1391),
.B(net1257),
.C(net10194),
.Y(net1397)
);

BUFx8_ASAP7_75t_R c1406(
.A(net10111),
.Y(net1398)
);

AND4x1_ASAP7_75t_R c1407(
.A(net1391),
.B(net1386),
.C(net1355),
.D(net9985),
.Y(net1399)
);

OAI21xp33_ASAP7_75t_R c1408(
.A1(net1304),
.A2(net1398),
.B(net1380),
.Y(net1400)
);

OAI21xp5_ASAP7_75t_R c1409(
.A1(net1400),
.A2(net270),
.B(net1392),
.Y(net1401)
);

AOI321xp33_ASAP7_75t_R c1410(
.A1(net1321),
.A2(net1400),
.A3(net1155),
.B1(net1348),
.B2(net9985),
.C(net10195),
.Y(net1402)
);

CKINVDCx10_ASAP7_75t_R c1411(
.A(net9281),
.Y(net1403)
);

CKINVDCx11_ASAP7_75t_R c1412(
.A(net9144),
.Y(net1404)
);

XOR2x2_ASAP7_75t_R c1413(
.A(net526),
.B(net1336),
.Y(net1405)
);

XOR2xp5_ASAP7_75t_R c1414(
.A(net381),
.B(net1340),
.Y(net1406)
);

OR3x1_ASAP7_75t_R c1415(
.A(net551),
.B(net537),
.C(net1250),
.Y(net1407)
);

CKINVDCx12_ASAP7_75t_R c1416(
.A(net9285),
.Y(net1408)
);

AND2x2_ASAP7_75t_R c1417(
.A(net1373),
.B(net9783),
.Y(net1409)
);

AND2x4_ASAP7_75t_R c1418(
.A(net1341),
.B(net1303),
.Y(net1410)
);

CKINVDCx14_ASAP7_75t_R c1419(
.A(net10139),
.Y(net1411)
);

CKINVDCx16_ASAP7_75t_R c1420(
.A(net1349),
.Y(net1412)
);

CKINVDCx20_ASAP7_75t_R c1421(
.A(net10193),
.Y(net1413)
);

AND2x6_ASAP7_75t_R c1422(
.A(net550),
.B(net444),
.Y(net1414)
);

CKINVDCx5p33_ASAP7_75t_R c1423(
.A(net1342),
.Y(net1415)
);

AND4x2_ASAP7_75t_R c1424(
.A(net506),
.B(net500),
.C(net356),
.D(net1348),
.Y(net1416)
);

OR3x2_ASAP7_75t_R c1425(
.A(net502),
.B(net484),
.C(net1386),
.Y(net1417)
);

CKINVDCx6p67_ASAP7_75t_R c1426(
.A(net10131),
.Y(net1418)
);

CKINVDCx8_ASAP7_75t_R c1427(
.A(net522),
.Y(net1419)
);

CKINVDCx9p33_ASAP7_75t_R c1428(
.A(net1345),
.Y(net1420)
);

HB1xp67_ASAP7_75t_R c1429(
.A(net10131),
.Y(net1421)
);

HB2xp67_ASAP7_75t_R c1430(
.A(net244),
.Y(net1422)
);

HB3xp67_ASAP7_75t_R c1431(
.A(net10165),
.Y(net1423)
);

HB4xp67_ASAP7_75t_R c1432(
.A(net9248),
.Y(net1424)
);

HAxp5_ASAP7_75t_R c1433(
.A(net1421),
.B(net445),
.CON(net1426),
.SN(net1425)
);

INVx11_ASAP7_75t_R c1434(
.A(net9251),
.Y(net1427)
);

NAND2x1_ASAP7_75t_R c1435(
.A(net1156),
.B(net1235),
.Y(net1428)
);

INVx13_ASAP7_75t_R c1436(
.A(net1427),
.Y(net1429)
);

SDFLx2_ASAP7_75t_R c1437(
.D(net1410),
.SE(net1425),
.SI(net10101),
.CLK(clk),
.QN(net1430)
);

INVx1_ASAP7_75t_R c1438(
.A(net515),
.Y(net1431)
);

INVx2_ASAP7_75t_R c1439(
.A(net1423),
.Y(net1432)
);

INVx3_ASAP7_75t_R c1440(
.A(net10139),
.Y(net1433)
);

NAND2x1p5_ASAP7_75t_R c1441(
.A(net1419),
.B(net244),
.Y(net1434)
);

INVx4_ASAP7_75t_R c1442(
.A(net489),
.Y(net1435)
);

INVx5_ASAP7_75t_R c1443(
.A(net1383),
.Y(net1436)
);

NAND2x2_ASAP7_75t_R c1444(
.A(net1411),
.B(net1421),
.Y(net1437)
);

NAND2xp33_ASAP7_75t_R c1445(
.A(net343),
.B(net1430),
.Y(net1438)
);

INVx6_ASAP7_75t_R c1446(
.A(net10131),
.Y(net1439)
);

OR3x4_ASAP7_75t_R c1447(
.A(net1435),
.B(net1415),
.C(net502),
.Y(net1440)
);

INVx8_ASAP7_75t_R c1448(
.A(net9281),
.Y(net1441)
);

AND3x1_ASAP7_75t_R c1449(
.A(net1406),
.B(net1436),
.C(net512),
.Y(net1442)
);

INVxp33_ASAP7_75t_R c1450(
.A(net10082),
.Y(net1443)
);

AO211x2_ASAP7_75t_R c1451(
.A1(net1235),
.A2(net1373),
.B(net9964),
.C(net10193),
.Y(net1444)
);

NAND2xp5_ASAP7_75t_R c1452(
.A(net1404),
.B(net558),
.Y(net1445)
);

NAND2xp67_ASAP7_75t_R c1453(
.A(net1422),
.B(net10194),
.Y(net1446)
);

INVxp67_ASAP7_75t_R c1454(
.A(net1386),
.Y(net1447)
);

ICGx5_ASAP7_75t_R c1455(
.ENA(net1436),
.SE(net501),
.CLK(clk),
.GCLK(net1448)
);

AND3x2_ASAP7_75t_R c1456(
.A(net1438),
.B(net1423),
.C(net1412),
.Y(net1449)
);

NOR2x1_ASAP7_75t_R c1457(
.A(net1257),
.B(net1448),
.Y(net1450)
);

BUFx10_ASAP7_75t_R c1458(
.A(net1346),
.Y(net1451)
);

NOR2x1p5_ASAP7_75t_R c1459(
.A(net426),
.B(net1446),
.Y(net1452)
);

BUFx12_ASAP7_75t_R c1460(
.A(net10101),
.Y(net1453)
);

BUFx12f_ASAP7_75t_R c1461(
.A(net1418),
.Y(net1454)
);

NOR2x2_ASAP7_75t_R c1462(
.A(net1428),
.B(net498),
.Y(net1455)
);

NOR2xp33_ASAP7_75t_R c1463(
.A(net1441),
.B(net429),
.Y(net1456)
);

BUFx16f_ASAP7_75t_R c1464(
.A(net1303),
.Y(net1457)
);

NOR2xp67_ASAP7_75t_R c1465(
.A(net1451),
.B(net558),
.Y(net1458)
);

OR2x2_ASAP7_75t_R c1466(
.A(net484),
.B(net560),
.Y(net1459)
);

BUFx24_ASAP7_75t_R c1467(
.A(net9144),
.Y(net1460)
);

BUFx2_ASAP7_75t_R c1468(
.A(net429),
.Y(net1461)
);

OR2x4_ASAP7_75t_R c1469(
.A(net1429),
.B(net1421),
.Y(net1462)
);

AOI33xp33_ASAP7_75t_R c1470(
.A1(net537),
.A2(net1435),
.A3(net1462),
.B1(net517),
.B2(net1449),
.B3(net534),
.Y(net1463)
);

AND3x4_ASAP7_75t_R c1471(
.A(net1431),
.B(net558),
.C(net1326),
.Y(net1464)
);

OR2x6_ASAP7_75t_R c1472(
.A(net1448),
.B(net1389),
.Y(net1465)
);

AO21x1_ASAP7_75t_R c1473(
.A1(net1147),
.A2(net551),
.B(net245),
.Y(net1466)
);

AO21x2_ASAP7_75t_R c1474(
.A1(net1445),
.A2(net537),
.B(net10194),
.Y(net1467)
);

XNOR2x1_ASAP7_75t_R c1475(
.B(net1426),
.A(net1449),
.Y(net1468)
);

AOI21x1_ASAP7_75t_R c1476(
.A1(net501),
.A2(net1456),
.B(net1460),
.Y(net1469)
);

XNOR2x2_ASAP7_75t_R c1477(
.A(net1468),
.B(net1449),
.Y(net1470)
);

AOI21xp33_ASAP7_75t_R c1478(
.A1(net1430),
.A2(net506),
.B(net1460),
.Y(net1471)
);

XNOR2xp5_ASAP7_75t_R c1479(
.A(net1443),
.B(net10082),
.Y(net1472)
);

XOR2x1_ASAP7_75t_R c1480(
.A(net1433),
.B(net1439),
.Y(net1473)
);

XOR2x2_ASAP7_75t_R c1481(
.A(net1452),
.B(net1458),
.Y(net1474)
);

SDFLx3_ASAP7_75t_R c1482(
.D(net1449),
.SE(net1346),
.SI(net1474),
.CLK(clk),
.QN(net1475)
);

AOI21xp5_ASAP7_75t_R c1483(
.A1(net1448),
.A2(net1475),
.B(net10126),
.Y(net1476)
);

OA222x2_ASAP7_75t_R c1484(
.A1(net1413),
.A2(net1464),
.B1(net1451),
.B2(net1160),
.C1(net1446),
.C2(net558),
.Y(net1477)
);

SDFLx4_ASAP7_75t_R c1485(
.D(net1323),
.SE(net1430),
.SI(net1474),
.CLK(clk),
.QN(net1478)
);

DFFASRHQNx1_ASAP7_75t_R c1486(
.D(net1478),
.RESETN(net1474),
.SETN(net9964),
.CLK(clk),
.QN(net1479)
);

SDFHx1_ASAP7_75t_R c1487(
.D(net1456),
.SE(net1423),
.SI(net1474),
.CLK(clk),
.QN(net1480)
);

AO22x1_ASAP7_75t_R c1488(
.A1(net1460),
.A2(net1445),
.B1(net1466),
.B2(net1449),
.Y(net1481)
);

OA33x2_ASAP7_75t_R c1489(
.A1(net1326),
.A2(net1439),
.A3(net1454),
.B1(net1474),
.B2(net558),
.B3(net534),
.Y(net1482)
);

FAx1_ASAP7_75t_R c1490(
.A(net1466),
.B(net1480),
.CI(net9956),
.SN(net1484),
.CON(net1483)
);

SDFHx2_ASAP7_75t_R c1491(
.D(net1453),
.SE(net1474),
.SI(net1483),
.CLK(clk),
.QN(net1485)
);

MAJIxp5_ASAP7_75t_R c1492(
.A(net1485),
.B(net1473),
.C(net9956),
.Y(net1486)
);

MAJx2_ASAP7_75t_R c1493(
.A(net1477),
.B(net1481),
.C(net10082),
.Y(net1487)
);

XOR2xp5_ASAP7_75t_R c1494(
.A(net1011),
.B(net613),
.Y(net1488)
);

BUFx3_ASAP7_75t_R c1495(
.A(net10152),
.Y(net1489)
);

BUFx4_ASAP7_75t_R c1496(
.A(net9264),
.Y(net1490)
);

AO22x2_ASAP7_75t_R c1497(
.A1(net553),
.A2(net626),
.B1(net483),
.B2(net629),
.Y(net1491)
);

BUFx4f_ASAP7_75t_R c1498(
.A(net1486),
.Y(net1492)
);

BUFx5_ASAP7_75t_R c1499(
.A(net586),
.Y(net1493)
);

BUFx6f_ASAP7_75t_R c1500(
.A(net632),
.Y(net1494)
);

BUFx8_ASAP7_75t_R c1501(
.A(net638),
.Y(net1495)
);

CKINVDCx10_ASAP7_75t_R c1502(
.A(net646),
.Y(net1496)
);

CKINVDCx11_ASAP7_75t_R c1503(
.A(net558),
.Y(net1497)
);

AND2x2_ASAP7_75t_R c1504(
.A(net598),
.B(net10177),
.Y(net1498)
);

CKINVDCx12_ASAP7_75t_R c1505(
.A(net1493),
.Y(net1499)
);

CKINVDCx14_ASAP7_75t_R c1506(
.A(net541),
.Y(net1500)
);

CKINVDCx16_ASAP7_75t_R c1507(
.A(net1495),
.Y(net1501)
);

MAJx3_ASAP7_75t_R c1508(
.A(net1493),
.B(net613),
.C(net1497),
.Y(net1502)
);

AND2x4_ASAP7_75t_R c1509(
.A(net625),
.B(net327),
.Y(net1503)
);

AND2x6_ASAP7_75t_R c1510(
.A(net578),
.B(net1479),
.Y(net1504)
);

CKINVDCx20_ASAP7_75t_R c1511(
.A(net10152),
.Y(net1505)
);

CKINVDCx5p33_ASAP7_75t_R c1512(
.A(net1484),
.Y(net1506)
);

CKINVDCx6p67_ASAP7_75t_R c1513(
.A(net9955),
.Y(net1507)
);

CKINVDCx8_ASAP7_75t_R c1514(
.A(net9955),
.Y(net1508)
);

CKINVDCx9p33_ASAP7_75t_R c1515(
.A(net10107),
.Y(net1509)
);

ICGx5p33DC_ASAP7_75t_R c1516(
.ENA(net1491),
.SE(net441),
.CLK(clk),
.GCLK(net1510)
);

HB1xp67_ASAP7_75t_R c1517(
.A(net1495),
.Y(net1511)
);

NAND3x1_ASAP7_75t_R c1518(
.A(net1502),
.B(net1510),
.C(net1488),
.Y(net1512)
);

HAxp5_ASAP7_75t_R c1519(
.A(net1266),
.B(net1493),
.CON(net1514),
.SN(net1513)
);

HB2xp67_ASAP7_75t_R c1520(
.A(net10126),
.Y(net1515)
);

NAND2x1_ASAP7_75t_R c1521(
.A(net614),
.B(net441),
.Y(net1516)
);

HB3xp67_ASAP7_75t_R c1522(
.A(net1472),
.Y(net1517)
);

HB4xp67_ASAP7_75t_R c1523(
.A(net1479),
.Y(net1518)
);

ICGx6p67DC_ASAP7_75t_R c1524(
.ENA(net1504),
.SE(net1510),
.CLK(clk),
.GCLK(net1519)
);

INVx11_ASAP7_75t_R c1525(
.A(net613),
.Y(net1520)
);

INVx13_ASAP7_75t_R c1526(
.A(net1475),
.Y(net1521)
);

INVx1_ASAP7_75t_R c1527(
.A(net9264),
.Y(net1522)
);

NAND2x1p5_ASAP7_75t_R c1528(
.A(net1498),
.B(net1382),
.Y(net1523)
);

NAND2x2_ASAP7_75t_R c1529(
.A(net1488),
.B(net585),
.Y(net1524)
);

NAND2xp33_ASAP7_75t_R c1530(
.A(net640),
.B(net1312),
.Y(net1525)
);

NAND2xp5_ASAP7_75t_R c1531(
.A(net1489),
.B(net1522),
.Y(net1526)
);

INVx2_ASAP7_75t_R c1532(
.A(net1516),
.Y(net1527)
);

INVx3_ASAP7_75t_R c1533(
.A(net1512),
.Y(net1528)
);

INVx4_ASAP7_75t_R c1534(
.A(net605),
.Y(net1529)
);

INVx5_ASAP7_75t_R c1535(
.A(net356),
.Y(net1530)
);

NAND2xp67_ASAP7_75t_R c1536(
.A(net1527),
.B(net1461),
.Y(net1531)
);

NOR2x1_ASAP7_75t_R c1537(
.A(net616),
.B(net1266),
.Y(net1532)
);

NOR2x1p5_ASAP7_75t_R c1538(
.A(net1506),
.B(net1454),
.Y(net1533)
);

INVx6_ASAP7_75t_R c1539(
.A(net10466),
.Y(net1534)
);

NOR2x2_ASAP7_75t_R c1540(
.A(net1505),
.B(net1531),
.Y(net1535)
);

NOR2xp33_ASAP7_75t_R c1541(
.A(net1461),
.B(net1506),
.Y(net1536)
);

NOR2xp67_ASAP7_75t_R c1542(
.A(net1525),
.B(net1528),
.Y(net1537)
);

OR2x2_ASAP7_75t_R c1543(
.A(net1497),
.B(net1530),
.Y(net1538)
);

INVx8_ASAP7_75t_R c1544(
.A(net10490),
.Y(net1539)
);

AO31x2_ASAP7_75t_R c1545(
.A1(net1520),
.A2(net1530),
.A3(net640),
.B(net1526),
.Y(net1540)
);

OR2x4_ASAP7_75t_R c1546(
.A(net1507),
.B(net1532),
.Y(net1541)
);

AOI221x1_ASAP7_75t_R c1547(
.A1(net1363),
.A2(net1536),
.B1(net1518),
.B2(net445),
.C(net606),
.Y(net1542)
);

INVxp33_ASAP7_75t_R c1548(
.A(net1529),
.Y(net1543)
);

OR2x6_ASAP7_75t_R c1549(
.A(net1415),
.B(net1479),
.Y(net1544)
);

XNOR2x1_ASAP7_75t_R c1550(
.B(net1524),
.A(net1493),
.Y(net1545)
);

INVxp67_ASAP7_75t_R c1551(
.A(net1533),
.Y(net1546)
);

XNOR2x2_ASAP7_75t_R c1552(
.A(net1523),
.B(net1363),
.Y(net1547)
);

XNOR2xp5_ASAP7_75t_R c1553(
.A(net441),
.B(net1521),
.Y(net1548)
);

BUFx10_ASAP7_75t_R c1554(
.A(net1503),
.Y(net1549)
);

XOR2x1_ASAP7_75t_R c1555(
.A(net1494),
.B(net9927),
.Y(net1550)
);

XOR2x2_ASAP7_75t_R c1556(
.A(net585),
.B(net1518),
.Y(net1551)
);

XOR2xp5_ASAP7_75t_R c1557(
.A(net1518),
.B(net1538),
.Y(net1552)
);

NAND3x2_ASAP7_75t_R c1558(
.B(net1519),
.C(net1550),
.A(net462),
.Y(net1553)
);

AND2x2_ASAP7_75t_R c1559(
.A(net1538),
.B(net1524),
.Y(net1554)
);

AOI211x1_ASAP7_75t_R c1560(
.A1(net1544),
.A2(net1477),
.B(net606),
.C(net1526),
.Y(net1555)
);

NAND3xp33_ASAP7_75t_R c1561(
.A(net1549),
.B(net1523),
.C(net1527),
.Y(net1556)
);

BUFx12_ASAP7_75t_R c1562(
.A(net10385),
.Y(net1557)
);

NOR3x1_ASAP7_75t_R c1563(
.A(net1547),
.B(net1551),
.C(net1519),
.Y(net1558)
);

AND2x4_ASAP7_75t_R c1564(
.A(net1539),
.B(net1363),
.Y(net1559)
);

AND2x6_ASAP7_75t_R c1565(
.A(net1550),
.B(net1556),
.Y(net1560)
);

BUFx12f_ASAP7_75t_R c1566(
.A(net1552),
.Y(net1561)
);

AOI211xp5_ASAP7_75t_R c1567(
.A1(net1528),
.A2(net1554),
.B(net1556),
.C(net1561),
.Y(net1562)
);

AOI221xp5_ASAP7_75t_R c1568(
.A1(net1494),
.A2(net1502),
.B1(net1011),
.B2(net1513),
.C(net1531),
.Y(net1563)
);

HAxp5_ASAP7_75t_R c1569(
.A(net1557),
.B(net9747),
.CON(net1565),
.SN(net1564)
);

AOI22x1_ASAP7_75t_R c1570(
.A1(net1556),
.A2(net1517),
.B1(net1561),
.B2(net10199),
.Y(net1566)
);

NAND2x1_ASAP7_75t_R c1571(
.A(net1547),
.B(net9747),
.Y(net1567)
);

NOR3x2_ASAP7_75t_R c1572(
.B(net556),
.C(net1564),
.A(net9927),
.Y(net1568)
);

NOR3xp33_ASAP7_75t_R c1573(
.A(net1500),
.B(net1568),
.C(net1526),
.Y(net1569)
);

AOI22xp33_ASAP7_75t_R c1574(
.A1(net1543),
.A2(net1565),
.B1(net1511),
.B2(net1526),
.Y(net1570)
);

NAND2x1p5_ASAP7_75t_R c1575(
.A(net1554),
.B(net10199),
.Y(net1571)
);

OA21x2_ASAP7_75t_R c1576(
.A1(net1517),
.A2(net1432),
.B(net1569),
.Y(net1572)
);

BUFx16f_ASAP7_75t_R c1577(
.A(net557),
.Y(net1573)
);

BUFx24_ASAP7_75t_R c1578(
.A(net633),
.Y(net1574)
);

OAI21x1_ASAP7_75t_R c1579(
.A1(net327),
.A2(net1312),
.B(net1505),
.Y(net1575)
);

BUFx2_ASAP7_75t_R c1580(
.A(net662),
.Y(net1576)
);

BUFx3_ASAP7_75t_R c1581(
.A(net676),
.Y(net1577)
);

BUFx4_ASAP7_75t_R c1582(
.A(net630),
.Y(net1578)
);

BUFx4f_ASAP7_75t_R c1583(
.A(net1160),
.Y(net1579)
);

BUFx5_ASAP7_75t_R c1584(
.A(net1579),
.Y(net1580)
);

NAND2x2_ASAP7_75t_R c1585(
.A(net654),
.B(net677),
.Y(net1581)
);

AOI22xp5_ASAP7_75t_R c1586(
.A1(net338),
.A2(net1579),
.B1(net693),
.B2(net1526),
.Y(net1582)
);

BUFx6f_ASAP7_75t_R c1587(
.A(net1581),
.Y(net1583)
);

BUFx8_ASAP7_75t_R c1588(
.A(net10199),
.Y(net1584)
);

CKINVDCx10_ASAP7_75t_R c1589(
.A(net705),
.Y(net1585)
);

CKINVDCx11_ASAP7_75t_R c1590(
.A(net572),
.Y(net1586)
);

CKINVDCx12_ASAP7_75t_R c1591(
.A(net1439),
.Y(net1587)
);

NAND2xp33_ASAP7_75t_R c1592(
.A(net1573),
.B(net1570),
.Y(net1588)
);

CKINVDCx14_ASAP7_75t_R c1593(
.A(net639),
.Y(net1589)
);

CKINVDCx16_ASAP7_75t_R c1594(
.A(net1505),
.Y(net1590)
);

NAND2xp5_ASAP7_75t_R c1595(
.A(net1590),
.B(net1568),
.Y(net1591)
);

CKINVDCx20_ASAP7_75t_R c1596(
.A(net1501),
.Y(net1592)
);

CKINVDCx5p33_ASAP7_75t_R c1597(
.A(net10056),
.Y(net1593)
);

CKINVDCx6p67_ASAP7_75t_R c1598(
.A(net1514),
.Y(net1594)
);

CKINVDCx8_ASAP7_75t_R c1599(
.A(net510),
.Y(net1595)
);

CKINVDCx9p33_ASAP7_75t_R c1600(
.A(net1574),
.Y(net1596)
);

HB1xp67_ASAP7_75t_R c1601(
.A(net700),
.Y(net1597)
);

HB2xp67_ASAP7_75t_R c1602(
.A(net10056),
.Y(net1598)
);

HB3xp67_ASAP7_75t_R c1603(
.A(net1496),
.Y(net1599)
);

HB4xp67_ASAP7_75t_R c1604(
.A(net682),
.Y(net1600)
);

NAND2xp67_ASAP7_75t_R c1605(
.A(net574),
.B(net700),
.Y(net1601)
);

OAI21xp33_ASAP7_75t_R c1606(
.A1(net705),
.A2(net664),
.B(net9927),
.Y(net1602)
);

INVx11_ASAP7_75t_R c1607(
.A(net1601),
.Y(net1603)
);

NOR2x1_ASAP7_75t_R c1608(
.A(net1575),
.B(net1600),
.Y(net1604)
);

INVx13_ASAP7_75t_R c1609(
.A(net1573),
.Y(net1605)
);

INVx1_ASAP7_75t_R c1610(
.A(net1597),
.Y(net1606)
);

NOR2x1p5_ASAP7_75t_R c1611(
.A(net1551),
.B(net1576),
.Y(net1607)
);

NOR2x2_ASAP7_75t_R c1612(
.A(net1539),
.B(net1580),
.Y(net1608)
);

NOR2xp33_ASAP7_75t_R c1613(
.A(net1492),
.B(net724),
.Y(net1609)
);

INVx2_ASAP7_75t_R c1614(
.A(net1579),
.Y(net1610)
);

INVx3_ASAP7_75t_R c1615(
.A(net517),
.Y(net1611)
);

NOR2xp67_ASAP7_75t_R c1616(
.A(net1530),
.B(net1564),
.Y(net1612)
);

INVx4_ASAP7_75t_R c1617(
.A(net10373),
.Y(net1613)
);

OR2x2_ASAP7_75t_R c1618(
.A(net1584),
.B(net498),
.Y(net1614)
);

OR2x4_ASAP7_75t_R c1619(
.A(net1596),
.B(net1597),
.Y(net1615)
);

INVx5_ASAP7_75t_R c1620(
.A(net10124),
.Y(net1616)
);

INVx6_ASAP7_75t_R c1621(
.A(net10100),
.Y(net1617)
);

INVx8_ASAP7_75t_R c1622(
.A(net708),
.Y(net1618)
);

INVxp33_ASAP7_75t_R c1623(
.A(net1589),
.Y(net1619)
);

INVxp67_ASAP7_75t_R c1624(
.A(net10376),
.Y(net1620)
);

ICGx8DC_ASAP7_75t_R c1625(
.ENA(net1603),
.SE(net1606),
.CLK(clk),
.GCLK(net1621)
);

BUFx10_ASAP7_75t_R c1626(
.A(net1577),
.Y(net1622)
);

OR2x6_ASAP7_75t_R c1627(
.A(net1607),
.B(net1608),
.Y(net1623)
);

OAI21xp5_ASAP7_75t_R c1628(
.A1(net1586),
.A2(net1606),
.B(net727),
.Y(net1624)
);

OR3x1_ASAP7_75t_R c1629(
.A(net1594),
.B(net1611),
.C(net1622),
.Y(net1625)
);

XNOR2x1_ASAP7_75t_R c1630(
.B(net703),
.A(net1611),
.Y(net1626)
);

XNOR2x2_ASAP7_75t_R c1631(
.A(net721),
.B(net1625),
.Y(net1627)
);

ICGx1_ASAP7_75t_R c1632(
.ENA(net1619),
.SE(net1606),
.CLK(clk),
.GCLK(net1628)
);

XNOR2xp5_ASAP7_75t_R c1633(
.A(net1590),
.B(net1576),
.Y(net1629)
);

BUFx12_ASAP7_75t_R c1634(
.A(net10525),
.Y(net1630)
);

XOR2x1_ASAP7_75t_R c1635(
.A(net1515),
.B(net1575),
.Y(net1631)
);

AOI31xp33_ASAP7_75t_R c1636(
.A1(net1613),
.A2(net1196),
.A3(net671),
.B(net633),
.Y(net1632)
);

XOR2x2_ASAP7_75t_R c1637(
.A(net629),
.B(net1530),
.Y(net1633)
);

ICGx2_ASAP7_75t_R c1638(
.ENA(net1632),
.SE(net1594),
.CLK(clk),
.GCLK(net1634)
);

XOR2xp5_ASAP7_75t_R c1639(
.A(net1609),
.B(net10184),
.Y(net1635)
);

OR3x2_ASAP7_75t_R c1640(
.A(net1599),
.B(net1355),
.C(net722),
.Y(net1636)
);

BUFx12f_ASAP7_75t_R c1641(
.A(net10572),
.Y(net1637)
);

AND2x2_ASAP7_75t_R c1642(
.A(net1580),
.B(net1634),
.Y(net1638)
);

BUFx16f_ASAP7_75t_R c1643(
.A(net10378),
.Y(net1639)
);

AOI31xp67_ASAP7_75t_R c1644(
.A1(net1578),
.A2(net1637),
.A3(net1622),
.B(net667),
.Y(net1640)
);

AND2x4_ASAP7_75t_R c1645(
.A(net1608),
.B(net1510),
.Y(net1641)
);

AND2x6_ASAP7_75t_R c1646(
.A(net1637),
.B(net10078),
.Y(net1642)
);

BUFx24_ASAP7_75t_R c1647(
.A(net1593),
.Y(net1643)
);

HAxp5_ASAP7_75t_R c1648(
.A(net1601),
.B(net1625),
.CON(net1644)
);

OR3x4_ASAP7_75t_R c1649(
.A(net1641),
.B(net1630),
.C(net1643),
.Y(net1645)
);

NAND2x1_ASAP7_75t_R c1650(
.A(net1642),
.B(net1618),
.Y(net1646)
);

AND3x1_ASAP7_75t_R c1651(
.A(net1633),
.B(net1638),
.C(net629),
.Y(net1647)
);

AND3x2_ASAP7_75t_R c1652(
.A(net1582),
.B(net517),
.C(net1641),
.Y(net1648)
);

AND3x4_ASAP7_75t_R c1653(
.A(net661),
.B(net1642),
.C(net1509),
.Y(net1649)
);

NAND2x1p5_ASAP7_75t_R c1654(
.A(net1639),
.B(net1575),
.Y(net1650)
);

NAND2x2_ASAP7_75t_R c1655(
.A(net1649),
.B(net1539),
.Y(net1651)
);

NAND2xp33_ASAP7_75t_R c1656(
.A(net1643),
.B(net651),
.Y(net1652)
);

ICGx2p67DC_ASAP7_75t_R c1657(
.ENA(net1648),
.SE(net1630),
.CLK(clk),
.GCLK(net1653)
);

OAI222xp33_ASAP7_75t_R c1658(
.A1(net1647),
.A2(net1601),
.B1(net1653),
.B2(net1350),
.C1(net686),
.C2(net1561),
.Y(net1654)
);

NAND4xp25_ASAP7_75t_R c1659(
.A(net556),
.B(net1651),
.C(net1597),
.D(net1625),
.Y(net1655)
);

AO21x1_ASAP7_75t_R c1660(
.A1(net771),
.A2(net798),
.B(net1611),
.Y(net1656)
);

BUFx2_ASAP7_75t_R c1661(
.A(net1448),
.Y(net1657)
);

NAND2xp5_ASAP7_75t_R c1662(
.A(net781),
.B(net10139),
.Y(net1658)
);

NAND2xp67_ASAP7_75t_R c1663(
.A(net1548),
.B(net808),
.Y(net1659)
);

AO21x2_ASAP7_75t_R c1664(
.A1(net1640),
.A2(net738),
.B(net10183),
.Y(net1660)
);

BUFx3_ASAP7_75t_R c1665(
.A(net1595),
.Y(net1661)
);

NOR2x1_ASAP7_75t_R c1666(
.A(net1450),
.B(net1351),
.Y(net1662)
);

NOR2x1p5_ASAP7_75t_R c1667(
.A(net649),
.B(net743),
.Y(net1663)
);

BUFx4_ASAP7_75t_R c1668(
.A(net9941),
.Y(net1664)
);

BUFx4f_ASAP7_75t_R c1669(
.A(net1565),
.Y(net1665)
);

BUFx5_ASAP7_75t_R c1670(
.A(net1510),
.Y(net1666)
);

BUFx6f_ASAP7_75t_R c1671(
.A(net1665),
.Y(net1667)
);

BUFx8_ASAP7_75t_R c1672(
.A(net9104),
.Y(net1668)
);

NOR2x2_ASAP7_75t_R c1673(
.A(net807),
.B(net1522),
.Y(net1669)
);

AOI311xp33_ASAP7_75t_R c1674(
.A1(net714),
.A2(net598),
.A3(net1448),
.B(net1526),
.C(net1664),
.Y(net1670)
);

CKINVDCx10_ASAP7_75t_R c1675(
.A(net1509),
.Y(net1671)
);

SDFHx3_ASAP7_75t_R c1676(
.D(net813),
.SE(net1628),
.SI(net778),
.CLK(clk),
.QN(net1672)
);

NOR2xp33_ASAP7_75t_R c1677(
.A(net1668),
.B(net1572),
.Y(net1673)
);

CKINVDCx11_ASAP7_75t_R c1678(
.A(net1619),
.Y(net1674)
);

CKINVDCx12_ASAP7_75t_R c1679(
.A(net1674),
.Y(net1675)
);

CKINVDCx14_ASAP7_75t_R c1680(
.A(net10097),
.Y(net1676)
);

CKINVDCx16_ASAP7_75t_R c1681(
.A(net9246),
.Y(net1677)
);

CKINVDCx20_ASAP7_75t_R c1682(
.A(net760),
.Y(net1678)
);

NAND4xp75_ASAP7_75t_R c1683(
.A(net1676),
.B(net1677),
.C(net735),
.D(net798),
.Y(net1679)
);

SDFHx4_ASAP7_75t_R c1684(
.D(net735),
.SE(net1677),
.SI(net711),
.CLK(clk),
.QN(net1680)
);

NOR2xp67_ASAP7_75t_R c1685(
.A(net1666),
.B(net1638),
.Y(net1681)
);

CKINVDCx5p33_ASAP7_75t_R c1686(
.A(net734),
.Y(net1682)
);

CKINVDCx6p67_ASAP7_75t_R c1687(
.A(net773),
.Y(net1683)
);

AOI21x1_ASAP7_75t_R c1688(
.A1(net808),
.A2(net1672),
.B(net10197),
.Y(net1684)
);

OR2x2_ASAP7_75t_R c1689(
.A(net1683),
.B(net1652),
.Y(net1685)
);

OR2x4_ASAP7_75t_R c1690(
.A(net1646),
.B(net790),
.Y(net1686)
);

OR2x6_ASAP7_75t_R c1691(
.A(net1661),
.B(net798),
.Y(net1687)
);

CKINVDCx8_ASAP7_75t_R c1692(
.A(net1660),
.Y(net1688)
);

XNOR2x1_ASAP7_75t_R c1693(
.B(net1622),
.A(net1675),
.Y(net1689)
);

CKINVDCx9p33_ASAP7_75t_R c1694(
.A(net778),
.Y(net1690)
);

HB1xp67_ASAP7_75t_R c1695(
.A(net9246),
.Y(net1691)
);

HB2xp67_ASAP7_75t_R c1696(
.A(net1667),
.Y(net1692)
);

XNOR2x2_ASAP7_75t_R c1697(
.A(net1688),
.B(net1685),
.Y(net1693)
);

HB3xp67_ASAP7_75t_R c1698(
.A(net764),
.Y(net1694)
);

HB4xp67_ASAP7_75t_R c1699(
.A(net1669),
.Y(net1695)
);

INVx11_ASAP7_75t_R c1700(
.A(net1677),
.Y(net1696)
);

INVx13_ASAP7_75t_R c1701(
.A(net1691),
.Y(net1697)
);

INVx1_ASAP7_75t_R c1702(
.A(net9270),
.Y(net1698)
);

OAI321xp33_ASAP7_75t_R c1703(
.A1(net1623),
.A2(net760),
.A3(net1677),
.B1(net1671),
.B2(net1637),
.C(net1664),
.Y(net1699)
);

INVx2_ASAP7_75t_R c1704(
.A(net9270),
.Y(net1700)
);

INVx3_ASAP7_75t_R c1705(
.A(net9250),
.Y(net1701)
);

XNOR2xp5_ASAP7_75t_R c1706(
.A(net1628),
.B(net1595),
.Y(net1702)
);

AOI32xp33_ASAP7_75t_R c1707(
.A1(net1698),
.A2(net1702),
.A3(net1160),
.B1(net1664),
.B2(net9683),
.Y(net1703)
);

INVx4_ASAP7_75t_R c1708(
.A(net9957),
.Y(net1704)
);

INVx5_ASAP7_75t_R c1709(
.A(net1696),
.Y(net1705)
);

INVx6_ASAP7_75t_R c1710(
.A(net1690),
.Y(net1706)
);

XOR2x1_ASAP7_75t_R c1711(
.A(net1704),
.B(net660),
.Y(net1707)
);

XOR2x2_ASAP7_75t_R c1712(
.A(net1681),
.B(net1680),
.Y(net1708)
);

INVx8_ASAP7_75t_R c1713(
.A(net1670),
.Y(net1709)
);

INVxp33_ASAP7_75t_R c1714(
.A(net786),
.Y(net1710)
);

XOR2xp5_ASAP7_75t_R c1715(
.A(net1574),
.B(net1707),
.Y(net1711)
);

AOI21xp33_ASAP7_75t_R c1716(
.A1(net1698),
.A2(net630),
.B(net10184),
.Y(net1712)
);

NOR4xp25_ASAP7_75t_R c1717(
.A(net1684),
.B(net1670),
.C(net1612),
.D(net1664),
.Y(net1713)
);

INVxp67_ASAP7_75t_R c1718(
.A(net1705),
.Y(net1714)
);

AOI21xp5_ASAP7_75t_R c1719(
.A1(net1686),
.A2(net1432),
.B(net9683),
.Y(net1715)
);

BUFx10_ASAP7_75t_R c1720(
.A(net1630),
.Y(net1716)
);

AND2x2_ASAP7_75t_R c1721(
.A(net1716),
.B(net1707),
.Y(net1717)
);

BUFx12_ASAP7_75t_R c1722(
.A(net1701),
.Y(net1718)
);

AND2x4_ASAP7_75t_R c1723(
.A(net1686),
.B(net10197),
.Y(net1719)
);

AND2x6_ASAP7_75t_R c1724(
.A(net1707),
.B(net1704),
.Y(net1720)
);

BUFx12f_ASAP7_75t_R c1725(
.A(net1656),
.Y(net1721)
);

FAx1_ASAP7_75t_R c1726(
.A(net1657),
.B(net1704),
.CI(net10179),
.SN(net1723),
.CON(net1722)
);

MAJIxp5_ASAP7_75t_R c1727(
.A(net1692),
.B(net1721),
.C(net747),
.Y(net1724)
);

HAxp5_ASAP7_75t_R c1728(
.A(net1715),
.B(net1682),
.CON(net1726),
.SN(net1725)
);

BUFx16f_ASAP7_75t_R c1729(
.A(net9250),
.Y(net1727)
);

NAND2x1_ASAP7_75t_R c1730(
.A(net1702),
.B(net1722),
.Y(net1728)
);

NAND2x1p5_ASAP7_75t_R c1731(
.A(net1713),
.B(net1710),
.Y(net1729)
);

NAND2x2_ASAP7_75t_R c1732(
.A(net1711),
.B(net1548),
.Y(net1730)
);

BUFx24_ASAP7_75t_R c1733(
.A(net9104),
.Y(net1731)
);

MAJx2_ASAP7_75t_R c1734(
.A(net1728),
.B(net1623),
.C(net1709),
.Y(net1732)
);

NAND2xp33_ASAP7_75t_R c1735(
.A(net1714),
.B(net1697),
.Y(net1733)
);

MAJx3_ASAP7_75t_R c1736(
.A(net1687),
.B(net1733),
.C(net1706),
.Y(net1734)
);

NAND2xp5_ASAP7_75t_R c1737(
.A(net1733),
.B(net1704),
.Y(net1735)
);

NAND3x1_ASAP7_75t_R c1738(
.A(net1522),
.B(net1658),
.C(net630),
.Y(net1736)
);

NAND2xp67_ASAP7_75t_R c1739(
.A(net763),
.B(net1724),
.Y(net1737)
);

NAND3x2_ASAP7_75t_R c1740(
.B(net1723),
.C(net1737),
.A(net1707),
.Y(net1738)
);

NAND3xp33_ASAP7_75t_R c1741(
.A(net1731),
.B(net1732),
.C(net1737),
.Y(net1739)
);

BUFx2_ASAP7_75t_R c1742(
.A(net10022),
.Y(net1740)
);

BUFx3_ASAP7_75t_R c1743(
.A(net1717),
.Y(net1741)
);

BUFx4_ASAP7_75t_R c1744(
.A(net1703),
.Y(net1742)
);

NOR2x1_ASAP7_75t_R c1745(
.A(net1706),
.B(net1561),
.Y(net1743)
);

BUFx4f_ASAP7_75t_R c1746(
.A(net1734),
.Y(net1744)
);

BUFx5_ASAP7_75t_R c1747(
.A(net1351),
.Y(net1745)
);

NOR2x1p5_ASAP7_75t_R c1748(
.A(net1675),
.B(net898),
.Y(net1746)
);

BUFx6f_ASAP7_75t_R c1749(
.A(net10528),
.Y(net1747)
);

BUFx8_ASAP7_75t_R c1750(
.A(net1723),
.Y(net1748)
);

ICGx3_ASAP7_75t_R c1751(
.ENA(net899),
.SE(net861),
.CLK(clk),
.GCLK(net1749)
);

NOR2x2_ASAP7_75t_R c1752(
.A(net1749),
.B(net1682),
.Y(net1750)
);

NOR2xp33_ASAP7_75t_R c1753(
.A(net1745),
.B(net1706),
.Y(net1751)
);

NOR2xp67_ASAP7_75t_R c1754(
.A(net781),
.B(net847),
.Y(net1752)
);

OR2x2_ASAP7_75t_R c1755(
.A(net1752),
.B(net865),
.Y(net1753)
);

CKINVDCx10_ASAP7_75t_R c1756(
.A(net9089),
.Y(net1754)
);

CKINVDCx11_ASAP7_75t_R c1757(
.A(net852),
.Y(net1755)
);

OR2x4_ASAP7_75t_R c1758(
.A(net1747),
.B(net784),
.Y(net1756)
);

CKINVDCx12_ASAP7_75t_R c1759(
.A(net809),
.Y(net1757)
);

OR2x6_ASAP7_75t_R c1760(
.A(net851),
.B(net1754),
.Y(net1758)
);

XNOR2x1_ASAP7_75t_R c1761(
.B(net785),
.A(net866),
.Y(net1759)
);

CKINVDCx14_ASAP7_75t_R c1762(
.A(net822),
.Y(net1760)
);

XNOR2x2_ASAP7_75t_R c1763(
.A(net1754),
.B(net1521),
.Y(net1761)
);

NOR4xp75_ASAP7_75t_R c1764(
.A(net1742),
.B(net899),
.C(net824),
.D(net849),
.Y(net1762)
);

XNOR2xp5_ASAP7_75t_R c1765(
.A(net865),
.B(net1637),
.Y(net1763)
);

CKINVDCx16_ASAP7_75t_R c1766(
.A(net1761),
.Y(net1764)
);

XOR2x1_ASAP7_75t_R c1767(
.A(net845),
.B(net1744),
.Y(net1765)
);

XOR2x2_ASAP7_75t_R c1768(
.A(net874),
.B(net1743),
.Y(net1766)
);

CKINVDCx20_ASAP7_75t_R c1769(
.A(net9888),
.Y(net1767)
);

XOR2xp5_ASAP7_75t_R c1770(
.A(net1682),
.B(net10201),
.Y(net1768)
);

NOR3x1_ASAP7_75t_R c1771(
.A(net672),
.B(net859),
.C(net1744),
.Y(net1769)
);

O2A1O1Ixp33_ASAP7_75t_R c1772(
.A1(net886),
.A2(net1753),
.B(net865),
.C(net1744),
.Y(net1770)
);

AND2x2_ASAP7_75t_R c1773(
.A(net1659),
.B(net1759),
.Y(net1771)
);

AND2x4_ASAP7_75t_R c1774(
.A(net846),
.B(net1749),
.Y(net1772)
);

AND2x6_ASAP7_75t_R c1775(
.A(net894),
.B(net1757),
.Y(net1773)
);

CKINVDCx5p33_ASAP7_75t_R c1776(
.A(net847),
.Y(net1774)
);

CKINVDCx6p67_ASAP7_75t_R c1777(
.A(net1638),
.Y(net1775)
);

HAxp5_ASAP7_75t_R c1778(
.A(net1758),
.B(net10201),
.CON(net1776)
);

NAND2x1_ASAP7_75t_R c1779(
.A(net874),
.B(net10202),
.Y(net1777)
);

NOR3x2_ASAP7_75t_R c1780(
.B(net1250),
.C(net1717),
.A(net749),
.Y(net1778)
);

CKINVDCx8_ASAP7_75t_R c1781(
.A(net1768),
.Y(net1779)
);

NAND2x1p5_ASAP7_75t_R c1782(
.A(net854),
.B(net893),
.Y(net1780)
);

CKINVDCx9p33_ASAP7_75t_R c1783(
.A(net9089),
.Y(net1781)
);

NAND2x2_ASAP7_75t_R c1784(
.A(net1637),
.B(net1764),
.Y(net1782)
);

NOR3xp33_ASAP7_75t_R c1785(
.A(net1764),
.B(net1749),
.C(net822),
.Y(net1783)
);

NAND2xp33_ASAP7_75t_R c1786(
.A(net1783),
.B(net1756),
.Y(net1784)
);

NAND2xp5_ASAP7_75t_R c1787(
.A(net1772),
.B(net809),
.Y(net1785)
);

OA21x2_ASAP7_75t_R c1788(
.A1(net1773),
.A2(net1760),
.B(net1767),
.Y(net1786)
);

NAND2xp67_ASAP7_75t_R c1789(
.A(net1778),
.B(net1756),
.Y(net1787)
);

NOR2x1_ASAP7_75t_R c1790(
.A(net664),
.B(net1749),
.Y(net1788)
);

NOR2x1p5_ASAP7_75t_R c1791(
.A(net849),
.B(net9957),
.Y(net1789)
);

NOR2x2_ASAP7_75t_R c1792(
.A(net1766),
.B(net810),
.Y(net1790)
);

NOR2xp33_ASAP7_75t_R c1793(
.A(net861),
.B(net9888),
.Y(net1791)
);

NOR2xp67_ASAP7_75t_R c1794(
.A(net1779),
.B(net1767),
.Y(net1792)
);

OR2x2_ASAP7_75t_R c1795(
.A(net1678),
.B(net1675),
.Y(net1793)
);

OAI21x1_ASAP7_75t_R c1796(
.A1(net870),
.A2(net898),
.B(net1774),
.Y(net1794)
);

OR2x4_ASAP7_75t_R c1797(
.A(net1741),
.B(net787),
.Y(net1795)
);

OR2x6_ASAP7_75t_R c1798(
.A(net1761),
.B(net9957),
.Y(net1796)
);

XNOR2x1_ASAP7_75t_R c1799(
.B(net730),
.A(net1760),
.Y(net1797)
);

HB1xp67_ASAP7_75t_R c1800(
.A(net10408),
.Y(net1798)
);

OAI33xp33_ASAP7_75t_R c1801(
.A1(net1763),
.A2(net897),
.A3(net836),
.B1(net824),
.B2(net1744),
.B3(net9920),
.Y(net1799)
);

XNOR2x2_ASAP7_75t_R c1802(
.A(net1792),
.B(net1761),
.Y(net1800)
);

OAI21xp33_ASAP7_75t_R c1803(
.A1(net1771),
.A2(net1450),
.B(net1785),
.Y(net1801)
);

ICGx4DC_ASAP7_75t_R c1804(
.ENA(net1767),
.SE(net1675),
.CLK(clk),
.GCLK(net1802)
);

SDFLx1_ASAP7_75t_R c1805(
.D(net898),
.SE(net1797),
.SI(net10201),
.CLK(clk),
.QN(net1803)
);

OAI21xp5_ASAP7_75t_R c1806(
.A1(net1795),
.A2(net1783),
.B(net886),
.Y(net1804)
);

XNOR2xp5_ASAP7_75t_R c1807(
.A(net1450),
.B(net1789),
.Y(net1805)
);

OR3x1_ASAP7_75t_R c1808(
.A(net1800),
.B(net1734),
.C(net1802),
.Y(net1806)
);

SDFLx2_ASAP7_75t_R c1809(
.D(net1806),
.SE(net866),
.SI(net1797),
.CLK(clk),
.QN(net1807)
);

OR3x2_ASAP7_75t_R c1810(
.A(net894),
.B(net1805),
.C(net9791),
.Y(net1808)
);

NAND5xp2_ASAP7_75t_R c1811(
.A(net1776),
.B(net1744),
.C(net1805),
.D(net873),
.E(net836),
.Y(net1809)
);

OR3x4_ASAP7_75t_R c1812(
.A(net1796),
.B(net1807),
.C(net10062),
.Y(net1810)
);

AND3x1_ASAP7_75t_R c1813(
.A(net1808),
.B(net1803),
.C(net1798),
.Y(net1811)
);

XOR2x1_ASAP7_75t_R c1814(
.A(net1808),
.B(net9922),
.Y(net1812)
);

O2A1O1Ixp5_ASAP7_75t_R c1815(
.A1(net1810),
.A2(net1756),
.B(net1803),
.C(net836),
.Y(net1813)
);

XOR2x2_ASAP7_75t_R c1816(
.A(net1789),
.B(net1678),
.Y(net1814)
);

XOR2xp5_ASAP7_75t_R c1817(
.A(net1814),
.B(net1764),
.Y(net1815)
);

OA211x2_ASAP7_75t_R c1818(
.A1(net1813),
.A2(net1752),
.B(net1787),
.C(net10202),
.Y(net1816)
);

AND2x2_ASAP7_75t_R c1819(
.A(net1755),
.B(net10203),
.Y(net1817)
);

NOR5xp2_ASAP7_75t_R c1820(
.A(net1743),
.B(net854),
.C(net1802),
.D(net1749),
.E(net836),
.Y(net1818)
);

AND2x4_ASAP7_75t_R c1821(
.A(net826),
.B(net1785),
.Y(net1819)
);

AND2x6_ASAP7_75t_R c1822(
.A(net1818),
.B(net9812),
.Y(net1820)
);

OA22x2_ASAP7_75t_R c1823(
.A1(net1805),
.A2(net1816),
.B1(net1798),
.B2(net1759),
.Y(net1821)
);

SDFLx3_ASAP7_75t_R c1824(
.D(net1821),
.SE(net1818),
.SI(net10062),
.CLK(clk),
.QN(net1822)
);

SDFLx4_ASAP7_75t_R c1825(
.D(net1753),
.SE(net1822),
.SI(net9782),
.CLK(clk),
.QN(net1823)
);

HB2xp67_ASAP7_75t_R c1826(
.A(net915),
.Y(net1824)
);

HB3xp67_ASAP7_75t_R c1827(
.A(net1824),
.Y(net1825)
);

HB4xp67_ASAP7_75t_R c1828(
.A(net16),
.Y(net1826)
);

INVx11_ASAP7_75t_R c1829(
.A(net1826),
.Y(net1827)
);

INVx13_ASAP7_75t_R c1830(
.A(net58),
.Y(net1828)
);

INVx1_ASAP7_75t_R c1831(
.A(net9190),
.Y(net1829)
);

ICGx4_ASAP7_75t_R c1832(
.ENA(net901),
.SE(net913),
.CLK(clk),
.GCLK(net1830)
);

INVx2_ASAP7_75t_R c1833(
.A(net7),
.Y(net1831)
);

INVx3_ASAP7_75t_R c1834(
.A(net1825),
.Y(net1832)
);

INVx4_ASAP7_75t_R c1835(
.A(net1831),
.Y(net1833)
);

INVx5_ASAP7_75t_R c1836(
.A(net984),
.Y(net1834)
);

INVx6_ASAP7_75t_R c1837(
.A(net9190),
.Y(net1835)
);

INVx8_ASAP7_75t_R c1838(
.A(net952),
.Y(net1836)
);

INVxp33_ASAP7_75t_R c1839(
.A(net966),
.Y(net1837)
);

HAxp5_ASAP7_75t_R c1840(
.A(net968),
.B(net1837),
.CON(net1839),
.SN(net1838)
);

INVxp67_ASAP7_75t_R c1841(
.A(net1835),
.Y(net1840)
);

NAND2x1_ASAP7_75t_R c1842(
.A(net937),
.B(net1838),
.Y(net1841)
);

BUFx10_ASAP7_75t_R c1843(
.A(net1830),
.Y(net1842)
);

NAND2x1p5_ASAP7_75t_R c1844(
.A(net927),
.B(net1825),
.Y(net1843)
);

AND3x2_ASAP7_75t_R c1845(
.A(net1835),
.B(net7),
.C(net9649),
.Y(net1844)
);

BUFx12_ASAP7_75t_R c1846(
.A(net9244),
.Y(net1845)
);

NAND2x2_ASAP7_75t_R c1847(
.A(net966),
.B(net1831),
.Y(net1846)
);

BUFx12f_ASAP7_75t_R c1848(
.A(net905),
.Y(net1847)
);

BUFx16f_ASAP7_75t_R c1849(
.A(net58),
.Y(net1848)
);

AND3x4_ASAP7_75t_R c1850(
.A(net915),
.B(net1842),
.C(net955),
.Y(net1849)
);

BUFx24_ASAP7_75t_R c1851(
.A(net1840),
.Y(net1850)
);

NAND2xp33_ASAP7_75t_R c1852(
.A(net939),
.B(net1834),
.Y(net1851)
);

NAND2xp5_ASAP7_75t_R c1853(
.A(net928),
.B(net1837),
.Y(net1852)
);

NAND2xp67_ASAP7_75t_R c1854(
.A(net984),
.B(net1834),
.Y(net1853)
);

BUFx2_ASAP7_75t_R c1855(
.A(net22),
.Y(net1854)
);

AO21x1_ASAP7_75t_R c1856(
.A1(net1848),
.A2(net1846),
.B(net913),
.Y(net1855)
);

AO21x2_ASAP7_75t_R c1857(
.A1(net1837),
.A2(net971),
.B(net30),
.Y(net1856)
);

ICGx5_ASAP7_75t_R c1858(
.ENA(net1853),
.SE(net1830),
.CLK(clk),
.GCLK(net1857)
);

NOR2x1_ASAP7_75t_R c1859(
.A(net1834),
.B(net1857),
.Y(net1858)
);

BUFx3_ASAP7_75t_R c1860(
.A(net9316),
.Y(net1859)
);

DFFASRHQNx1_ASAP7_75t_R c1861(
.D(net1836),
.RESETN(net1828),
.SETN(net979),
.CLK(clk),
.QN(net1860)
);

BUFx4_ASAP7_75t_R c1862(
.A(net1860),
.Y(net1861)
);

NOR2x1p5_ASAP7_75t_R c1863(
.A(net1852),
.B(net9649),
.Y(net1862)
);

ICGx5p33DC_ASAP7_75t_R c1864(
.ENA(net1851),
.SE(net1859),
.CLK(clk),
.GCLK(net1863)
);

ICGx6p67DC_ASAP7_75t_R c1865(
.ENA(net1825),
.SE(net1858),
.CLK(clk),
.GCLK(net1864)
);

BUFx4f_ASAP7_75t_R c1866(
.A(net9316),
.Y(net1865)
);

NOR2x2_ASAP7_75t_R c1867(
.A(net1854),
.B(net1859),
.Y(net1866)
);

BUFx5_ASAP7_75t_R c1868(
.A(net1843),
.Y(net1867)
);

BUFx6f_ASAP7_75t_R c1869(
.A(net952),
.Y(net1868)
);

NOR2xp33_ASAP7_75t_R c1870(
.A(net1849),
.B(net907),
.Y(net1869)
);

BUFx8_ASAP7_75t_R c1871(
.A(net1850),
.Y(net1870)
);

NOR2xp67_ASAP7_75t_R c1872(
.A(net1829),
.B(net905),
.Y(net1871)
);

OR2x2_ASAP7_75t_R c1873(
.A(net1846),
.B(net966),
.Y(net1872)
);

CKINVDCx10_ASAP7_75t_R c1874(
.A(net1824),
.Y(net1873)
);

ICGx8DC_ASAP7_75t_R c1875(
.ENA(net1853),
.SE(net975),
.CLK(clk),
.GCLK(net1874)
);

OR2x4_ASAP7_75t_R c1876(
.A(net1863),
.B(net1871),
.Y(net1875)
);

OR2x6_ASAP7_75t_R c1877(
.A(net1871),
.B(net1840),
.Y(net1876)
);

AOI21x1_ASAP7_75t_R c1878(
.A1(net941),
.A2(net1871),
.B(net1837),
.Y(net1877)
);

CKINVDCx11_ASAP7_75t_R c1879(
.A(net9232),
.Y(net1878)
);

ICGx1_ASAP7_75t_R c1880(
.ENA(net1873),
.SE(net1877),
.CLK(clk),
.GCLK(net1879)
);

AOI21xp33_ASAP7_75t_R c1881(
.A1(net1859),
.A2(net1840),
.B(net970),
.Y(net1880)
);

CKINVDCx12_ASAP7_75t_R c1882(
.A(net1876),
.Y(net1881)
);

ICGx2_ASAP7_75t_R c1883(
.ENA(net1868),
.SE(net1857),
.CLK(clk),
.GCLK(net1882)
);

ICGx2p67DC_ASAP7_75t_R c1884(
.ENA(net1836),
.SE(net1882),
.CLK(clk),
.GCLK(net1883)
);

XNOR2x1_ASAP7_75t_R c1885(
.B(net1881),
.A(net1849),
.Y(net1884)
);

CKINVDCx14_ASAP7_75t_R c1886(
.A(net1876),
.Y(net1885)
);

CKINVDCx16_ASAP7_75t_R c1887(
.A(net1878),
.Y(net1886)
);

XNOR2x2_ASAP7_75t_R c1888(
.A(net1830),
.B(net1859),
.Y(net1887)
);

XNOR2xp5_ASAP7_75t_R c1889(
.A(net1847),
.B(net1850),
.Y(net1888)
);

XOR2x1_ASAP7_75t_R c1890(
.A(net1887),
.B(net1884),
.Y(net1889)
);

AOI21xp5_ASAP7_75t_R c1891(
.A1(net1888),
.A2(net1881),
.B(net971),
.Y(net1890)
);

ICGx3_ASAP7_75t_R c1892(
.ENA(net971),
.SE(net1872),
.CLK(clk),
.GCLK(net1891)
);

ICGx4DC_ASAP7_75t_R c1893(
.ENA(net1872),
.SE(net1865),
.CLK(clk),
.GCLK(net1892)
);

XOR2x2_ASAP7_75t_R c1894(
.A(net1892),
.B(net1874),
.Y(net1893)
);

OA221x2_ASAP7_75t_R c1895(
.A1(net931),
.A2(net1890),
.B1(net58),
.B2(net1869),
.C(net47),
.Y(net1894)
);

FAx1_ASAP7_75t_R c1896(
.A(net1870),
.B(net1860),
.CI(net9756),
.SN(net1896),
.CON(net1895)
);

SDFHx1_ASAP7_75t_R c1897(
.D(net1885),
.SE(net1858),
.SI(net1895),
.CLK(clk),
.QN(net1897)
);

XOR2xp5_ASAP7_75t_R c1898(
.A(net22),
.B(net1885),
.Y(net1898)
);

SDFHx2_ASAP7_75t_R c1899(
.D(net1874),
.SE(net1897),
.SI(net1853),
.CLK(clk),
.QN(net1899)
);

MAJIxp5_ASAP7_75t_R c1900(
.A(net1899),
.B(net1875),
.C(net9849),
.Y(net1900)
);

ICGx4_ASAP7_75t_R c1901(
.ENA(net1828),
.SE(net1868),
.CLK(clk),
.GCLK(net1901)
);

SDFHx3_ASAP7_75t_R c1902(
.D(net1899),
.SE(net1889),
.SI(net1898),
.CLK(clk),
.QN(net1902)
);

AND2x2_ASAP7_75t_R c1903(
.A(net1889),
.B(net1902),
.Y(net1903)
);

SDFHx4_ASAP7_75t_R c1904(
.D(net1863),
.SE(net1887),
.SI(net1890),
.CLK(clk),
.QN(net1904)
);

AND2x4_ASAP7_75t_R c1905(
.A(net1865),
.B(net9748),
.Y(net1905)
);

AO222x2_ASAP7_75t_R c1906(
.A1(in25),
.A2(net1887),
.B1(net1902),
.B2(net913),
.C1(net925),
.C2(net1833),
.Y(net1906)
);

MAJx2_ASAP7_75t_R c1907(
.A(net1870),
.B(net1882),
.C(net1905),
.Y(net1907)
);

OA31x2_ASAP7_75t_R c1908(
.A1(net1902),
.A2(net1900),
.A3(net1907),
.B1(net1856),
.Y(net1908)
);

CKINVDCx20_ASAP7_75t_R c1909(
.A(net1053),
.Y(net1909)
);

AND2x6_ASAP7_75t_R c1910(
.A(net47),
.B(net59),
.Y(net1910)
);

CKINVDCx5p33_ASAP7_75t_R c1911(
.A(net1871),
.Y(net1911)
);

HAxp5_ASAP7_75t_R c1912(
.A(net1905),
.B(net1008),
.CON(net1913),
.SN(net1912)
);

CKINVDCx6p67_ASAP7_75t_R c1913(
.A(net102),
.Y(net1914)
);

CKINVDCx8_ASAP7_75t_R c1914(
.A(net1911),
.Y(net1915)
);

CKINVDCx9p33_ASAP7_75t_R c1915(
.A(net115),
.Y(net1916)
);

NAND2x1_ASAP7_75t_R c1916(
.A(net1913),
.B(net10186),
.Y(net1917)
);

HB1xp67_ASAP7_75t_R c1917(
.A(net9197),
.Y(net1918)
);

NAND2x1p5_ASAP7_75t_R c1918(
.A(net925),
.B(net1905),
.Y(net1919)
);

HB2xp67_ASAP7_75t_R c1919(
.A(net9133),
.Y(net1920)
);

NAND2x2_ASAP7_75t_R c1920(
.A(net1920),
.B(net1064),
.Y(net1921)
);

HB3xp67_ASAP7_75t_R c1921(
.A(net9133),
.Y(net1922)
);

HB4xp67_ASAP7_75t_R c1922(
.A(net1866),
.Y(net1923)
);

INVx11_ASAP7_75t_R c1923(
.A(net1901),
.Y(net1924)
);

INVx13_ASAP7_75t_R c1924(
.A(net1914),
.Y(net1925)
);

INVx1_ASAP7_75t_R c1925(
.A(net1907),
.Y(net1926)
);

SDFLx1_ASAP7_75t_R c1926(
.D(net102),
.SE(net1043),
.SI(net1917),
.CLK(clk),
.QN(net1927)
);

INVx2_ASAP7_75t_R c1927(
.A(net9212),
.Y(net1928)
);

NAND2xp33_ASAP7_75t_R c1928(
.A(net1893),
.B(net1924),
.Y(net1929)
);

NAND2xp5_ASAP7_75t_R c1929(
.A(net1043),
.B(net1866),
.Y(net1930)
);

INVx3_ASAP7_75t_R c1930(
.A(net9213),
.Y(net1931)
);

INVx4_ASAP7_75t_R c1931(
.A(net9213),
.Y(net1932)
);

NAND2xp67_ASAP7_75t_R c1932(
.A(net1913),
.B(net955),
.Y(net1933)
);

NOR2x1_ASAP7_75t_R c1933(
.A(net1042),
.B(net47),
.Y(net1934)
);

INVx5_ASAP7_75t_R c1934(
.A(net1882),
.Y(net1935)
);

NOR2x1p5_ASAP7_75t_R c1935(
.A(net1916),
.B(net1901),
.Y(net1936)
);

INVx6_ASAP7_75t_R c1936(
.A(net955),
.Y(net1937)
);

ICGx5_ASAP7_75t_R c1937(
.ENA(net1042),
.SE(net1936),
.CLK(clk),
.GCLK(net1938)
);

INVx8_ASAP7_75t_R c1938(
.A(net10498),
.Y(net1939)
);

INVxp33_ASAP7_75t_R c1939(
.A(net1923),
.Y(net1940)
);

INVxp67_ASAP7_75t_R c1940(
.A(net10407),
.Y(net1941)
);

MAJx3_ASAP7_75t_R c1941(
.A(net1937),
.B(net1940),
.C(net999),
.Y(net1942)
);

NAND3x1_ASAP7_75t_R c1942(
.A(net1910),
.B(net1929),
.C(net1898),
.Y(net1943)
);

BUFx10_ASAP7_75t_R c1943(
.A(net1918),
.Y(net1944)
);

BUFx12_ASAP7_75t_R c1944(
.A(net1917),
.Y(net1945)
);

NOR2x2_ASAP7_75t_R c1945(
.A(net1837),
.B(net88),
.Y(net1946)
);

SDFLx2_ASAP7_75t_R c1946(
.D(net1924),
.SE(net1852),
.SI(net9748),
.CLK(clk),
.QN(net1947)
);

BUFx12f_ASAP7_75t_R c1947(
.A(net1934),
.Y(net1948)
);

BUFx16f_ASAP7_75t_R c1948(
.A(net1942),
.Y(net1949)
);

BUFx24_ASAP7_75t_R c1949(
.A(net1064),
.Y(net1950)
);

NOR2xp33_ASAP7_75t_R c1950(
.A(net1932),
.B(net1914),
.Y(net1951)
);

NAND3x2_ASAP7_75t_R c1951(
.B(net949),
.C(net1911),
.A(net1893),
.Y(net1952)
);

BUFx2_ASAP7_75t_R c1952(
.A(net1933),
.Y(net1953)
);

BUFx3_ASAP7_75t_R c1953(
.A(net1934),
.Y(net1954)
);

BUFx4_ASAP7_75t_R c1954(
.A(net967),
.Y(net1955)
);

BUFx4f_ASAP7_75t_R c1955(
.A(net10436),
.Y(net1956)
);

BUFx5_ASAP7_75t_R c1956(
.A(net1929),
.Y(net1957)
);

NOR2xp67_ASAP7_75t_R c1957(
.A(net1957),
.B(net9849),
.Y(net1958)
);

BUFx6f_ASAP7_75t_R c1958(
.A(net1832),
.Y(net1959)
);

ICGx5p33DC_ASAP7_75t_R c1959(
.ENA(net1951),
.SE(net983),
.CLK(clk),
.GCLK(net1960)
);

BUFx8_ASAP7_75t_R c1960(
.A(net999),
.Y(net1961)
);

NAND3xp33_ASAP7_75t_R c1961(
.A(net1956),
.B(net1042),
.C(net1882),
.Y(net1962)
);

ICGx6p67DC_ASAP7_75t_R c1962(
.ENA(net1940),
.SE(net1856),
.CLK(clk),
.GCLK(net1963)
);

OR2x2_ASAP7_75t_R c1963(
.A(net1915),
.B(net1924),
.Y(net1964)
);

OR2x4_ASAP7_75t_R c1964(
.A(net1959),
.B(net1961),
.Y(net1965)
);

CKINVDCx10_ASAP7_75t_R c1965(
.A(net1937),
.Y(net1966)
);

OR2x6_ASAP7_75t_R c1966(
.A(net1924),
.B(net1960),
.Y(net1967)
);

XNOR2x1_ASAP7_75t_R c1967(
.B(net1053),
.A(net1927),
.Y(net1968)
);

XNOR2x2_ASAP7_75t_R c1968(
.A(net1960),
.B(net1943),
.Y(net1969)
);

XNOR2xp5_ASAP7_75t_R c1969(
.A(net1955),
.B(net1963),
.Y(net1970)
);

CKINVDCx11_ASAP7_75t_R c1970(
.A(net1943),
.Y(net1971)
);

CKINVDCx12_ASAP7_75t_R c1971(
.A(net9864),
.Y(net1972)
);

ICGx8DC_ASAP7_75t_R c1972(
.ENA(net1969),
.SE(net1909),
.CLK(clk),
.GCLK(net1973)
);

XOR2x1_ASAP7_75t_R c1973(
.A(net1909),
.B(net1963),
.Y(net1974)
);

NOR3x1_ASAP7_75t_R c1974(
.A(net1946),
.B(net1973),
.C(net1968),
.Y(net1975)
);

XOR2x2_ASAP7_75t_R c1975(
.A(net1964),
.B(net1966),
.Y(net1976)
);

XOR2xp5_ASAP7_75t_R c1976(
.A(net1968),
.B(net1963),
.Y(net1977)
);

ICGx1_ASAP7_75t_R c1977(
.ENA(net1950),
.SE(net1962),
.CLK(clk),
.GCLK(net1978)
);

NOR3x2_ASAP7_75t_R c1978(
.B(net1935),
.C(net1974),
.A(net925),
.Y(net1979)
);

NOR3xp33_ASAP7_75t_R c1979(
.A(net1925),
.B(net1960),
.C(net1896),
.Y(net1980)
);

AND2x2_ASAP7_75t_R c1980(
.A(net1973),
.B(net9889),
.Y(net1981)
);

AO33x2_ASAP7_75t_R c1981(
.A1(net1979),
.A2(net1972),
.A3(net1912),
.B1(net1844),
.B2(net994),
.B3(net1915),
.Y(net1982)
);

AND2x4_ASAP7_75t_R c1982(
.A(net1928),
.B(net1978),
.Y(net1983)
);

OA21x2_ASAP7_75t_R c1983(
.A1(net1977),
.A2(net1982),
.B(net1962),
.Y(net1984)
);

OAI21x1_ASAP7_75t_R c1984(
.A1(net998),
.A2(net1982),
.B(net1960),
.Y(net1985)
);

OAI21xp33_ASAP7_75t_R c1985(
.A1(net119),
.A2(net1978),
.B(net1980),
.Y(net1986)
);

AND2x6_ASAP7_75t_R c1986(
.A(net1985),
.B(net10187),
.Y(net1987)
);

HAxp5_ASAP7_75t_R c1987(
.A(net1967),
.B(net1980),
.CON(net1989),
.SN(net1988)
);

NAND2x1_ASAP7_75t_R c1988(
.A(net1958),
.B(net1987),
.Y(net1990)
);

OAI21xp5_ASAP7_75t_R c1989(
.A1(net1910),
.A2(net1989),
.B(net1980),
.Y(net1991)
);

OR3x1_ASAP7_75t_R c1990(
.A(net1949),
.B(net1991),
.C(net10186),
.Y(net1992)
);

OR3x2_ASAP7_75t_R c1991(
.A(net1991),
.B(net1978),
.C(net9702),
.Y(net1993)
);

CKINVDCx14_ASAP7_75t_R c1992(
.A(net2073),
.Y(net1994)
);

CKINVDCx16_ASAP7_75t_R c1993(
.A(net1905),
.Y(net1995)
);

CKINVDCx20_ASAP7_75t_R c1994(
.A(net1090),
.Y(net1996)
);

CKINVDCx5p33_ASAP7_75t_R c1995(
.A(net2078),
.Y(net1997)
);

ICGx2_ASAP7_75t_R c1996(
.ENA(net2068),
.SE(net1092),
.CLK(clk),
.GCLK(net1998)
);

CKINVDCx6p67_ASAP7_75t_R c1997(
.A(net1107),
.Y(net1999)
);

CKINVDCx8_ASAP7_75t_R c1998(
.A(net10565),
.Y(net2000)
);

NAND2x1p5_ASAP7_75t_R c1999(
.A(net1998),
.B(net9821),
.Y(net2001)
);

CKINVDCx9p33_ASAP7_75t_R c2000(
.A(net1134),
.Y(net2002)
);

OR3x4_ASAP7_75t_R c2001(
.A(net2002),
.B(net1995),
.C(net1869),
.Y(net2003)
);

NAND2x2_ASAP7_75t_R c2002(
.A(net2000),
.B(net2060),
.Y(net2004)
);

NAND2xp33_ASAP7_75t_R c2003(
.A(net2003),
.B(net202),
.Y(net2005)
);

HB1xp67_ASAP7_75t_R c2004(
.A(net9103),
.Y(net2006)
);

HB2xp67_ASAP7_75t_R c2005(
.A(net9103),
.Y(net2007)
);

OAI221xp5_ASAP7_75t_R c2006(
.A1(net1076),
.A2(net1108),
.B1(net1999),
.B2(net2052),
.C(net180),
.Y(net2008)
);

NAND2xp5_ASAP7_75t_R c2007(
.A(net2078),
.B(net2073),
.Y(net2009)
);

HB3xp67_ASAP7_75t_R c2008(
.A(net1994),
.Y(net2010)
);

HB4xp67_ASAP7_75t_R c2009(
.A(net9212),
.Y(net2011)
);

NAND2xp67_ASAP7_75t_R c2010(
.A(net2004),
.B(net2011),
.Y(net2012)
);

OAI311xp33_ASAP7_75t_R c2011(
.A1(net2010),
.A2(net115),
.A3(net224),
.B1(net1051),
.C1(net2052),
.Y(net2013)
);

NOR2x1_ASAP7_75t_R c2012(
.A(net2007),
.B(net1898),
.Y(net2014)
);

AND3x1_ASAP7_75t_R c2013(
.A(net1995),
.B(net1089),
.C(net1861),
.Y(net2015)
);

NOR2x1p5_ASAP7_75t_R c2014(
.A(net2009),
.B(net2001),
.Y(net2016)
);

NOR2x2_ASAP7_75t_R c2015(
.A(net2057),
.B(net2011),
.Y(net2017)
);

AND3x2_ASAP7_75t_R c2016(
.A(net1983),
.B(net2009),
.C(net1111),
.Y(net2018)
);

INVx11_ASAP7_75t_R c2017(
.A(net10453),
.Y(net2019)
);

NOR2xp33_ASAP7_75t_R c2018(
.A(net2064),
.B(net1895),
.Y(net2020)
);

AND3x4_ASAP7_75t_R c2019(
.A(net2016),
.B(net2004),
.C(net1052),
.Y(net2021)
);

NOR2xp67_ASAP7_75t_R c2020(
.A(net2011),
.B(net2078),
.Y(net2022)
);

OR2x2_ASAP7_75t_R c2021(
.A(net1122),
.B(net2002),
.Y(net2023)
);

OR2x4_ASAP7_75t_R c2022(
.A(net2020),
.B(net2065),
.Y(net2024)
);

INVx13_ASAP7_75t_R c2023(
.A(net2012),
.Y(net2025)
);

INVx1_ASAP7_75t_R c2024(
.A(net2025),
.Y(net2026)
);

OR2x6_ASAP7_75t_R c2025(
.A(net2013),
.B(net2019),
.Y(net2027)
);

AO21x1_ASAP7_75t_R c2026(
.A1(net2015),
.A2(net2020),
.B(net9950),
.Y(net2028)
);

XNOR2x1_ASAP7_75t_R c2027(
.B(net1953),
.A(net1131),
.Y(net2029)
);

AO21x2_ASAP7_75t_R c2028(
.A1(net1092),
.A2(net2020),
.B(net2065),
.Y(net2030)
);

INVx2_ASAP7_75t_R c2029(
.A(net2023),
.Y(net2031)
);

INVx3_ASAP7_75t_R c2030(
.A(net1998),
.Y(net2032)
);

XNOR2x2_ASAP7_75t_R c2031(
.A(net2074),
.B(net2004),
.Y(net2033)
);

INVx4_ASAP7_75t_R c2032(
.A(net10415),
.Y(net2034)
);

AOI21x1_ASAP7_75t_R c2033(
.A1(net2015),
.A2(net2012),
.B(net1005),
.Y(net2035)
);

INVx5_ASAP7_75t_R c2034(
.A(net9267),
.Y(net2036)
);

SDFLx3_ASAP7_75t_R c2035(
.D(net2029),
.SE(net2031),
.SI(net1122),
.CLK(clk),
.QN(net2037)
);

AOI21xp33_ASAP7_75t_R c2036(
.A1(net2001),
.A2(net2033),
.B(net2071),
.Y(net2038)
);

OAI211xp5_ASAP7_75t_R c2037(
.A1(net1083),
.A2(net2037),
.B(net2021),
.C(net2071),
.Y(net2039)
);

XNOR2xp5_ASAP7_75t_R c2038(
.A(net2024),
.B(net2037),
.Y(net2040)
);

AOI21xp5_ASAP7_75t_R c2039(
.A1(net2030),
.A2(net1998),
.B(net1938),
.Y(net2041)
);

XOR2x1_ASAP7_75t_R c2040(
.A(net202),
.B(net2033),
.Y(net2042)
);

FAx1_ASAP7_75t_R c2041(
.A(net1052),
.B(net1994),
.CI(net10126),
.SN(net2044),
.CON(net2043)
);

MAJIxp5_ASAP7_75t_R c2042(
.A(net2022),
.B(net59),
.C(net10064),
.Y(net2045)
);

MAJx2_ASAP7_75t_R c2043(
.A(net2028),
.B(net2043),
.C(net10064),
.Y(net2046)
);

OAI32xp33_ASAP7_75t_R c2044(
.A1(net2006),
.A2(net2035),
.A3(net1867),
.B1(net1135),
.B2(net1057),
.Y(net2047)
);

OAI22x1_ASAP7_75t_R c2045(
.A1(net2032),
.A2(net2070),
.B1(net2045),
.B2(net10205),
.Y(net2048)
);

XOR2x2_ASAP7_75t_R c2046(
.A(net2026),
.B(net10205),
.Y(net2049)
);

OR5x1_ASAP7_75t_R c2047(
.A(net2013),
.B(net1148),
.C(net2049),
.D(net119),
.E(net10205),
.Y(net2050)
);

OR5x2_ASAP7_75t_R c2048(
.A(net2021),
.B(net1147),
.C(net2049),
.D(net1915),
.E(net10205),
.Y(net2051)
);

INVx6_ASAP7_75t_R c2049(
.A(net1098),
.Y(net2052)
);

MAJx3_ASAP7_75t_R c2050(
.A(net1990),
.B(net1114),
.C(net1827),
.Y(net2053)
);

INVx8_ASAP7_75t_R c2051(
.A(net9315),
.Y(net2054)
);

XOR2xp5_ASAP7_75t_R c2052(
.A(net1075),
.B(net202),
.Y(net2055)
);

INVxp33_ASAP7_75t_R c2053(
.A(net9291),
.Y(net2056)
);

INVxp67_ASAP7_75t_R c2054(
.A(net1148),
.Y(net2057)
);

BUFx10_ASAP7_75t_R c2055(
.A(net10136),
.Y(net2058)
);

NAND3x1_ASAP7_75t_R c2056(
.A(net1108),
.B(net1149),
.C(net1092),
.Y(net2059)
);

BUFx12_ASAP7_75t_R c2057(
.A(net1106),
.Y(net2060)
);

A2O1A1O1Ixp25_ASAP7_75t_R c2058(
.A1(net201),
.A2(net1869),
.B(net1972),
.C(net1107),
.D(net2060),
.Y(net2061)
);

BUFx12f_ASAP7_75t_R c2059(
.A(net2060),
.Y(net2062)
);

AND2x2_ASAP7_75t_R c2060(
.A(net1057),
.B(net1076),
.Y(net2063)
);

AND2x4_ASAP7_75t_R c2061(
.A(net1022),
.B(net2060),
.Y(net2064)
);

AND2x6_ASAP7_75t_R c2062(
.A(net1136),
.B(net2052),
.Y(net2065)
);

NAND3x2_ASAP7_75t_R c2063(
.B(net88),
.C(net1134),
.A(net2062),
.Y(net2066)
);

HAxp5_ASAP7_75t_R c2064(
.A(net2065),
.B(net1957),
.CON(net2068),
.SN(net2067)
);

BUFx16f_ASAP7_75t_R c2065(
.A(net2066),
.Y(net2069)
);

NAND2x1_ASAP7_75t_R c2066(
.A(net2066),
.B(net1090),
.Y(net2070)
);

NAND2x1p5_ASAP7_75t_R c2067(
.A(net2056),
.B(net1896),
.Y(net2071)
);

NAND2x2_ASAP7_75t_R c2068(
.A(net1110),
.B(net2069),
.Y(net2072)
);

BUFx24_ASAP7_75t_R c2069(
.A(net9202),
.Y(net2073)
);

BUFx2_ASAP7_75t_R c2070(
.A(net2069),
.Y(net2074)
);

NAND2xp33_ASAP7_75t_R c2071(
.A(net2052),
.B(net2055),
.Y(net2075)
);

NAND3xp33_ASAP7_75t_R c2072(
.A(net1111),
.B(net1896),
.C(net1905),
.Y(net2076)
);

BUFx3_ASAP7_75t_R c2073(
.A(net10479),
.Y(net2077)
);

BUFx4_ASAP7_75t_R c2074(
.A(net10453),
.Y(net2078)
);

BUFx4f_ASAP7_75t_R c2075(
.A(net9904),
.Y(net2079)
);

BUFx5_ASAP7_75t_R c2076(
.A(net224),
.Y(net2080)
);

BUFx6f_ASAP7_75t_R c2077(
.A(net10031),
.Y(net2081)
);

NAND2xp5_ASAP7_75t_R c2078(
.A(net1206),
.B(net1099),
.Y(net2082)
);

NAND2xp67_ASAP7_75t_R c2079(
.A(net2082),
.B(net2036),
.Y(net2083)
);

BUFx8_ASAP7_75t_R c2080(
.A(net298),
.Y(net2084)
);

NOR2x1_ASAP7_75t_R c2081(
.A(net1020),
.B(net1229),
.Y(net2085)
);

CKINVDCx10_ASAP7_75t_R c2082(
.A(net2002),
.Y(net2086)
);

CKINVDCx11_ASAP7_75t_R c2083(
.A(net1179),
.Y(net2087)
);

CKINVDCx12_ASAP7_75t_R c2084(
.A(net1201),
.Y(net2088)
);

NOR3x1_ASAP7_75t_R c2085(
.A(net1997),
.B(net1938),
.C(net2031),
.Y(net2089)
);

NOR2x1p5_ASAP7_75t_R c2086(
.A(net1100),
.B(net1833),
.Y(net2090)
);

CKINVDCx14_ASAP7_75t_R c2087(
.A(net2086),
.Y(net2091)
);

CKINVDCx16_ASAP7_75t_R c2088(
.A(net2082),
.Y(net2092)
);

CKINVDCx20_ASAP7_75t_R c2089(
.A(net2044),
.Y(net2093)
);

CKINVDCx5p33_ASAP7_75t_R c2090(
.A(net1132),
.Y(net2094)
);

CKINVDCx6p67_ASAP7_75t_R c2091(
.A(net1232),
.Y(net2095)
);

NOR2x2_ASAP7_75t_R c2092(
.A(net1204),
.B(net2079),
.Y(net2096)
);

CKINVDCx8_ASAP7_75t_R c2093(
.A(net2084),
.Y(net2097)
);

CKINVDCx9p33_ASAP7_75t_R c2094(
.A(net1938),
.Y(net2098)
);

HB1xp67_ASAP7_75t_R c2095(
.A(net10497),
.Y(net2099)
);

HB2xp67_ASAP7_75t_R c2096(
.A(net10031),
.Y(net2100)
);

SDFLx4_ASAP7_75t_R c2097(
.D(net1214),
.SE(net2049),
.SI(net10176),
.CLK(clk),
.QN(net2101)
);

NOR2xp33_ASAP7_75t_R c2098(
.A(net1996),
.B(net72),
.Y(net2102)
);

ICGx2p67DC_ASAP7_75t_R c2099(
.ENA(net1149),
.SE(net2060),
.CLK(clk),
.GCLK(net2103)
);

NOR2xp67_ASAP7_75t_R c2100(
.A(net2097),
.B(net1927),
.Y(net2104)
);

HB3xp67_ASAP7_75t_R c2101(
.A(net1999),
.Y(net2105)
);

HB4xp67_ASAP7_75t_R c2102(
.A(net2087),
.Y(net2106)
);

OR2x2_ASAP7_75t_R c2103(
.A(net1234),
.B(net2093),
.Y(net2107)
);

INVx11_ASAP7_75t_R c2104(
.A(net2102),
.Y(net2108)
);

AOI222xp33_ASAP7_75t_R c2105(
.A1(net2108),
.A2(net2097),
.B1(net2091),
.B2(net1999),
.C1(net1168),
.C2(net1160),
.Y(net2109)
);

INVx13_ASAP7_75t_R c2106(
.A(net1221),
.Y(net2110)
);

OR2x4_ASAP7_75t_R c2107(
.A(net2107),
.B(net9904),
.Y(net2111)
);

OR2x6_ASAP7_75t_R c2108(
.A(net1173),
.B(net1038),
.Y(net2112)
);

XNOR2x1_ASAP7_75t_R c2109(
.B(net1827),
.A(net2080),
.Y(net2113)
);

XNOR2x2_ASAP7_75t_R c2110(
.A(net2105),
.B(net2094),
.Y(net2114)
);

XNOR2xp5_ASAP7_75t_R c2111(
.A(net2093),
.B(net1944),
.Y(net2115)
);

XOR2x1_ASAP7_75t_R c2112(
.A(net2115),
.B(net2103),
.Y(net2116)
);

INVx1_ASAP7_75t_R c2113(
.A(net10006),
.Y(net2117)
);

NOR3x2_ASAP7_75t_R c2114(
.B(net2106),
.C(net2098),
.A(net2049),
.Y(net2118)
);

INVx2_ASAP7_75t_R c2115(
.A(net9225),
.Y(net2119)
);

INVx3_ASAP7_75t_R c2116(
.A(net9973),
.Y(net2120)
);

XOR2x2_ASAP7_75t_R c2117(
.A(net2054),
.B(net298),
.Y(net2121)
);

XOR2xp5_ASAP7_75t_R c2118(
.A(net2119),
.B(net2113),
.Y(net2122)
);

NOR3xp33_ASAP7_75t_R c2119(
.A(net1944),
.B(net1867),
.C(net9825),
.Y(net2123)
);

INVx4_ASAP7_75t_R c2120(
.A(net2099),
.Y(net2124)
);

INVx5_ASAP7_75t_R c2121(
.A(net2092),
.Y(net2125)
);

INVx6_ASAP7_75t_R c2122(
.A(net2080),
.Y(net2126)
);

AND2x2_ASAP7_75t_R c2123(
.A(net1183),
.B(net2125),
.Y(net2127)
);

OA21x2_ASAP7_75t_R c2124(
.A1(net241),
.A2(net1183),
.B(net298),
.Y(net2128)
);

OAI22xp33_ASAP7_75t_R c2125(
.A1(net2109),
.A2(net2100),
.B1(net1206),
.B2(net1915),
.Y(net2129)
);

AND2x4_ASAP7_75t_R c2126(
.A(net2128),
.B(net9904),
.Y(net2130)
);

OAI22xp5_ASAP7_75t_R c2127(
.A1(net299),
.A2(net2125),
.B1(net2100),
.B2(net2084),
.Y(net2131)
);

AND2x6_ASAP7_75t_R c2128(
.A(net2122),
.B(net2084),
.Y(net2132)
);

DFFASRHQNx1_ASAP7_75t_R c2129(
.D(net1184),
.RESETN(net2109),
.SETN(net2128),
.CLK(clk),
.QN(net2133)
);

INVx8_ASAP7_75t_R c2130(
.A(net10063),
.Y(net2134)
);

INVxp33_ASAP7_75t_R c2131(
.A(net9844),
.Y(net2135)
);

ICGx3_ASAP7_75t_R c2132(
.ENA(net2133),
.SE(net1140),
.CLK(clk),
.GCLK(net2136)
);

HAxp5_ASAP7_75t_R c2133(
.A(net2134),
.B(net2087),
.CON(net2138),
.SN(net2137)
);

NAND2x1_ASAP7_75t_R c2134(
.A(net2116),
.B(net2130),
.Y(net2139)
);

OAI31xp33_ASAP7_75t_R c2135(
.A1(net2101),
.A2(net2127),
.A3(net1205),
.B(net2130),
.Y(net2140)
);

NAND2x1p5_ASAP7_75t_R c2136(
.A(net2104),
.B(net2136),
.Y(net2141)
);

NAND2x2_ASAP7_75t_R c2137(
.A(net2112),
.B(net2141),
.Y(net2142)
);

OAI21x1_ASAP7_75t_R c2138(
.A1(net2094),
.A2(net2133),
.B(net2071),
.Y(net2143)
);

OAI21xp33_ASAP7_75t_R c2139(
.A1(net2139),
.A2(net2130),
.B(net2119),
.Y(net2144)
);

SDFHx1_ASAP7_75t_R c2140(
.D(net2135),
.SE(net2141),
.SI(net1149),
.CLK(clk),
.QN(net2145)
);

OAI21xp5_ASAP7_75t_R c2141(
.A1(net2120),
.A2(net2110),
.B(net2037),
.Y(net2146)
);

NAND2xp33_ASAP7_75t_R c2142(
.A(net2113),
.B(net2139),
.Y(net2147)
);

NAND2xp5_ASAP7_75t_R c2143(
.A(net1197),
.B(net2048),
.Y(net2148)
);

NAND2xp67_ASAP7_75t_R c2144(
.A(net2132),
.B(net2147),
.Y(net2149)
);

OR3x1_ASAP7_75t_R c2145(
.A(net276),
.B(net2138),
.C(net2131),
.Y(net2150)
);

OR3x2_ASAP7_75t_R c2146(
.A(net2098),
.B(net2140),
.C(net2145),
.Y(net2151)
);

OR3x4_ASAP7_75t_R c2147(
.A(net2137),
.B(net1867),
.C(net10095),
.Y(net2152)
);

NOR2x1_ASAP7_75t_R c2148(
.A(net2142),
.B(net1997),
.Y(net2153)
);

NOR2x1p5_ASAP7_75t_R c2149(
.A(net2100),
.B(net9977),
.Y(net2154)
);

AND3x1_ASAP7_75t_R c2150(
.A(net2138),
.B(net2127),
.C(net2080),
.Y(net2155)
);

NOR2x2_ASAP7_75t_R c2151(
.A(net2140),
.B(net2101),
.Y(net2156)
);

NOR2xp33_ASAP7_75t_R c2152(
.A(net2121),
.B(net1999),
.Y(net2157)
);

NOR2xp67_ASAP7_75t_R c2153(
.A(net2156),
.B(net2122),
.Y(net2158)
);

SDFHx2_ASAP7_75t_R c2154(
.D(net2157),
.SE(net2154),
.SI(net2158),
.CLK(clk),
.QN(net2159)
);

OR2x2_ASAP7_75t_R c2155(
.A(net1205),
.B(net2108),
.Y(net2160)
);

OR2x4_ASAP7_75t_R c2156(
.A(net1131),
.B(net2080),
.Y(net2161)
);

OR2x6_ASAP7_75t_R c2157(
.A(net2160),
.B(net2101),
.Y(net2162)
);

INVxp67_ASAP7_75t_R c2158(
.A(net1982),
.Y(net2163)
);

BUFx10_ASAP7_75t_R c2159(
.A(net188),
.Y(net2164)
);

XNOR2x1_ASAP7_75t_R c2160(
.B(net1298),
.A(net315),
.Y(net2165)
);

BUFx12_ASAP7_75t_R c2161(
.A(net34),
.Y(net2166)
);

BUFx12f_ASAP7_75t_R c2162(
.A(net2039),
.Y(net2167)
);

BUFx16f_ASAP7_75t_R c2163(
.A(net9120),
.Y(net2168)
);

XNOR2x2_ASAP7_75t_R c2164(
.A(net1170),
.B(net2126),
.Y(net2169)
);

AND3x2_ASAP7_75t_R c2165(
.A(net1222),
.B(net2031),
.C(net2166),
.Y(net2170)
);

BUFx24_ASAP7_75t_R c2166(
.A(net2165),
.Y(net2171)
);

XNOR2xp5_ASAP7_75t_R c2167(
.A(net2168),
.B(net1280),
.Y(net2172)
);

ICGx4DC_ASAP7_75t_R c2168(
.ENA(net1314),
.SE(net2148),
.CLK(clk),
.GCLK(net2173)
);

XOR2x1_ASAP7_75t_R c2169(
.A(net2164),
.B(net9996),
.Y(net2174)
);

XOR2x2_ASAP7_75t_R c2170(
.A(net2162),
.B(net276),
.Y(net2175)
);

XOR2xp5_ASAP7_75t_R c2171(
.A(net2136),
.B(net358),
.Y(net2176)
);

BUFx2_ASAP7_75t_R c2172(
.A(net9963),
.Y(net2177)
);

AND2x2_ASAP7_75t_R c2173(
.A(net2177),
.B(net1256),
.Y(net2178)
);

AND2x4_ASAP7_75t_R c2174(
.A(net2167),
.B(net1147),
.Y(net2179)
);

AND2x6_ASAP7_75t_R c2175(
.A(net1289),
.B(net1313),
.Y(net2180)
);

BUFx3_ASAP7_75t_R c2176(
.A(net10176),
.Y(net2181)
);

HAxp5_ASAP7_75t_R c2177(
.A(net9896),
.B(net10176),
.CON(net2183),
.SN(net2182)
);

BUFx4_ASAP7_75t_R c2178(
.A(net9120),
.Y(net2184)
);

NAND2x1_ASAP7_75t_R c2179(
.A(net2184),
.B(net2182),
.Y(net2185)
);

BUFx4f_ASAP7_75t_R c2180(
.A(net1299),
.Y(net2186)
);

NAND2x1p5_ASAP7_75t_R c2181(
.A(net332),
.B(net2163),
.Y(net2187)
);

BUFx5_ASAP7_75t_R c2182(
.A(net10527),
.Y(net2188)
);

AND3x4_ASAP7_75t_R c2183(
.A(net1157),
.B(net1290),
.C(net1135),
.Y(net2189)
);

NAND2x2_ASAP7_75t_R c2184(
.A(net2079),
.B(net1258),
.Y(net2190)
);

NAND2xp33_ASAP7_75t_R c2185(
.A(net2169),
.B(net1289),
.Y(net2191)
);

NAND2xp5_ASAP7_75t_R c2186(
.A(net2031),
.B(net2187),
.Y(net2192)
);

NAND2xp67_ASAP7_75t_R c2187(
.A(net1248),
.B(net1258),
.Y(net2193)
);

NOR2x1_ASAP7_75t_R c2188(
.A(net2171),
.B(net2191),
.Y(net2194)
);

BUFx6f_ASAP7_75t_R c2189(
.A(net10411),
.Y(net2195)
);

BUFx8_ASAP7_75t_R c2190(
.A(net1196),
.Y(net2196)
);

NOR2x1p5_ASAP7_75t_R c2191(
.A(net1051),
.B(net2188),
.Y(net2197)
);

NOR2x2_ASAP7_75t_R c2192(
.A(net1258),
.B(net315),
.Y(net2198)
);

CKINVDCx10_ASAP7_75t_R c2193(
.A(net365),
.Y(net2199)
);

NOR2xp33_ASAP7_75t_R c2194(
.A(net2194),
.B(net1282),
.Y(net2200)
);

CKINVDCx11_ASAP7_75t_R c2195(
.A(net2175),
.Y(net2201)
);

NOR2xp67_ASAP7_75t_R c2196(
.A(net2190),
.B(net2167),
.Y(net2202)
);

OR2x2_ASAP7_75t_R c2197(
.A(net1308),
.B(net2169),
.Y(net2203)
);

OR2x4_ASAP7_75t_R c2198(
.A(net2172),
.B(net2126),
.Y(net2204)
);

OR2x6_ASAP7_75t_R c2199(
.A(net2185),
.B(net2147),
.Y(net2205)
);

XNOR2x1_ASAP7_75t_R c2200(
.B(net2202),
.A(net2169),
.Y(net2206)
);

XNOR2x2_ASAP7_75t_R c2201(
.A(net9896),
.B(net9982),
.Y(net2207)
);

AO21x1_ASAP7_75t_R c2202(
.A1(net2190),
.A2(net2203),
.B(net9961),
.Y(net2208)
);

XNOR2xp5_ASAP7_75t_R c2203(
.A(net389),
.B(net2207),
.Y(net2209)
);

CKINVDCx12_ASAP7_75t_R c2204(
.A(net10457),
.Y(net2210)
);

AO21x2_ASAP7_75t_R c2205(
.A1(net2179),
.A2(net2201),
.B(net2191),
.Y(net2211)
);

XOR2x1_ASAP7_75t_R c2206(
.A(net1272),
.B(net2173),
.Y(net2212)
);

AND5x1_ASAP7_75t_R c2207(
.A(net2096),
.B(net2136),
.C(net1251),
.D(net2145),
.E(net1317),
.Y(net2213)
);

XOR2x2_ASAP7_75t_R c2208(
.A(net2181),
.B(net2210),
.Y(net2214)
);

AOI321xp33_ASAP7_75t_R c2209(
.A1(net1135),
.A2(net2178),
.A3(net2188),
.B1(net2163),
.B2(net2167),
.C(net10192),
.Y(net2215)
);

XOR2xp5_ASAP7_75t_R c2210(
.A(net2208),
.B(net9982),
.Y(net2216)
);

AND2x2_ASAP7_75t_R c2211(
.A(net1944),
.B(net2191),
.Y(net2217)
);

AND2x4_ASAP7_75t_R c2212(
.A(net1294),
.B(net2193),
.Y(net2218)
);

AND2x6_ASAP7_75t_R c2213(
.A(net2103),
.B(net2204),
.Y(net2219)
);

HAxp5_ASAP7_75t_R c2214(
.A(net2212),
.B(net2207),
.CON(net2221),
.SN(net2220)
);

AND5x2_ASAP7_75t_R c2215(
.A(net2217),
.B(net2195),
.C(net1287),
.D(net389),
.E(net10190),
.Y(net2222)
);

AOI21x1_ASAP7_75t_R c2216(
.A1(net2196),
.A2(net1167),
.B(net10161),
.Y(net2223)
);

NAND2x1_ASAP7_75t_R c2217(
.A(net2190),
.B(net10099),
.Y(net2224)
);

NAND2x1p5_ASAP7_75t_R c2218(
.A(net315),
.B(net1277),
.Y(net2225)
);

NAND2x2_ASAP7_75t_R c2219(
.A(net2209),
.B(net2224),
.Y(net2226)
);

AOI21xp33_ASAP7_75t_R c2220(
.A1(net2188),
.A2(net2190),
.B(net2163),
.Y(net2227)
);

SDFHx3_ASAP7_75t_R c2221(
.D(net2192),
.SE(net2188),
.SI(net9956),
.CLK(clk),
.QN(net2228)
);

NAND2xp33_ASAP7_75t_R c2222(
.A(net1167),
.B(net2130),
.Y(net2229)
);

NAND2xp5_ASAP7_75t_R c2223(
.A(net358),
.B(net2212),
.Y(net2230)
);

NAND2xp67_ASAP7_75t_R c2224(
.A(net1267),
.B(net1190),
.Y(net2231)
);

NOR2x1_ASAP7_75t_R c2225(
.A(net2207),
.B(net2173),
.Y(net2232)
);

ICGx4_ASAP7_75t_R c2226(
.ENA(net2192),
.SE(net2212),
.CLK(clk),
.GCLK(net2233)
);

NOR2x1p5_ASAP7_75t_R c2227(
.A(net2229),
.B(net2228),
.Y(net2234)
);

AOI21xp5_ASAP7_75t_R c2228(
.A1(net2166),
.A2(net270),
.B(net2220),
.Y(net2235)
);

AOI33xp33_ASAP7_75t_R c2229(
.A1(net2228),
.A2(net1212),
.A3(net2207),
.B1(net1190),
.B2(net2167),
.B3(net1170),
.Y(net2236)
);

FAx1_ASAP7_75t_R c2230(
.A(net2178),
.B(net1170),
.CI(net1314),
.SN(net2238),
.CON(net2237)
);

NOR2x2_ASAP7_75t_R c2231(
.A(net2238),
.B(net2221),
.Y(net2239)
);

OA222x2_ASAP7_75t_R c2232(
.A1(net2237),
.A2(net2173),
.B1(net1038),
.B2(net2235),
.C1(net9950),
.C2(net10208),
.Y(net2240)
);

SDFHx4_ASAP7_75t_R c2233(
.D(net2091),
.SE(net2208),
.SI(net2187),
.CLK(clk),
.QN(net2241)
);

SDFLx1_ASAP7_75t_R c2234(
.D(net2049),
.SE(net2241),
.SI(net2239),
.CLK(clk),
.QN(net2242)
);

MAJIxp5_ASAP7_75t_R c2235(
.A(net2234),
.B(net2242),
.C(net2039),
.Y(net2243)
);

MAJx2_ASAP7_75t_R c2236(
.A(net1287),
.B(net10106),
.C(net10208),
.Y(net2244)
);

SDFLx2_ASAP7_75t_R c2237(
.D(net2236),
.SE(net2239),
.SI(net1982),
.CLK(clk),
.QN(net2245)
);

OA33x2_ASAP7_75t_R c2238(
.A1(net2243),
.A2(net2221),
.A3(net1308),
.B1(net2239),
.B2(net2145),
.B3(net10208),
.Y(net2246)
);

OAI31xp67_ASAP7_75t_R c2239(
.A1(net2058),
.A2(net2214),
.A3(net2220),
.B(net1251),
.Y(net2247)
);

MAJx3_ASAP7_75t_R c2240(
.A(net1051),
.B(net2239),
.C(net10076),
.Y(net2248)
);

CKINVDCx14_ASAP7_75t_R c2241(
.A(net2187),
.Y(net2249)
);

CKINVDCx16_ASAP7_75t_R c2242(
.A(net10089),
.Y(net2250)
);

CKINVDCx20_ASAP7_75t_R c2243(
.A(net9948),
.Y(net2251)
);

CKINVDCx5p33_ASAP7_75t_R c2244(
.A(net2244),
.Y(net2252)
);

NOR2xp33_ASAP7_75t_R c2245(
.A(net2197),
.B(net2252),
.Y(net2253)
);

NAND3x1_ASAP7_75t_R c2246(
.A(net2148),
.B(net2197),
.C(net2241),
.Y(net2254)
);

CKINVDCx6p67_ASAP7_75t_R c2247(
.A(net2221),
.Y(net2255)
);

NAND3x2_ASAP7_75t_R c2248(
.B(net1360),
.C(net1317),
.A(net338),
.Y(net2256)
);

AO221x1_ASAP7_75t_R c2249(
.A1(net2225),
.A2(net2255),
.B1(net2145),
.B2(net1338),
.C(net1365),
.Y(net2257)
);

NOR2xp67_ASAP7_75t_R c2250(
.A(net2233),
.B(net411),
.Y(net2258)
);

CKINVDCx8_ASAP7_75t_R c2251(
.A(net10071),
.Y(net2259)
);

NAND3xp33_ASAP7_75t_R c2252(
.A(net2147),
.B(net1365),
.C(net10195),
.Y(net2260)
);

OR2x2_ASAP7_75t_R c2253(
.A(net1340),
.B(net9956),
.Y(net2261)
);

CKINVDCx9p33_ASAP7_75t_R c2254(
.A(net1099),
.Y(net2262)
);

HB1xp67_ASAP7_75t_R c2255(
.A(net2241),
.Y(net2263)
);

HB2xp67_ASAP7_75t_R c2256(
.A(net2263),
.Y(net2264)
);

OR2x4_ASAP7_75t_R c2257(
.A(net443),
.B(net1398),
.Y(net2265)
);

NOR3x1_ASAP7_75t_R c2258(
.A(net1395),
.B(net428),
.C(net1313),
.Y(net2266)
);

HB3xp67_ASAP7_75t_R c2259(
.A(net9150),
.Y(net2267)
);

HB4xp67_ASAP7_75t_R c2260(
.A(net2257),
.Y(net2268)
);

INVx11_ASAP7_75t_R c2261(
.A(net9150),
.Y(net2269)
);

INVx13_ASAP7_75t_R c2262(
.A(net2203),
.Y(net2270)
);

OR2x6_ASAP7_75t_R c2263(
.A(net2126),
.B(net2262),
.Y(net2271)
);

XNOR2x1_ASAP7_75t_R c2264(
.B(net2251),
.A(net2255),
.Y(net2272)
);

XNOR2x2_ASAP7_75t_R c2265(
.A(net2141),
.B(net404),
.Y(net2273)
);

XNOR2xp5_ASAP7_75t_R c2266(
.A(net2256),
.B(net2265),
.Y(net2274)
);

ICGx5_ASAP7_75t_R c2267(
.ENA(net2268),
.SE(net2148),
.CLK(clk),
.GCLK(net2275)
);

XOR2x1_ASAP7_75t_R c2268(
.A(net2273),
.B(net2167),
.Y(net2276)
);

INVx1_ASAP7_75t_R c2269(
.A(net1400),
.Y(net2277)
);

NOR3x2_ASAP7_75t_R c2270(
.B(net428),
.C(net1378),
.A(net2230),
.Y(net2278)
);

XOR2x2_ASAP7_75t_R c2271(
.A(net2259),
.B(net2264),
.Y(net2279)
);

XOR2xp5_ASAP7_75t_R c2272(
.A(net1379),
.B(net2145),
.Y(net2280)
);

AND2x2_ASAP7_75t_R c2273(
.A(net2279),
.B(net2174),
.Y(net2281)
);

AND2x4_ASAP7_75t_R c2274(
.A(net1317),
.B(net9726),
.Y(net2282)
);

AND2x6_ASAP7_75t_R c2275(
.A(net2269),
.B(net2272),
.Y(net2283)
);

HAxp5_ASAP7_75t_R c2276(
.A(net2283),
.B(net2272),
.CON(net2285),
.SN(net2284)
);

NAND2x1_ASAP7_75t_R c2277(
.A(net2281),
.B(net2227),
.Y(net2286)
);

NAND2x1p5_ASAP7_75t_R c2278(
.A(net2174),
.B(net1170),
.Y(net2287)
);

NAND2x2_ASAP7_75t_R c2279(
.A(net1317),
.B(net1371),
.Y(net2288)
);

NAND2xp33_ASAP7_75t_R c2280(
.A(net1282),
.B(net2281),
.Y(net2289)
);

SDFLx3_ASAP7_75t_R c2281(
.D(net2286),
.SE(net2258),
.SI(net1168),
.CLK(clk),
.QN(net2290)
);

INVx2_ASAP7_75t_R c2282(
.A(net411),
.Y(net2291)
);

INVx3_ASAP7_75t_R c2283(
.A(net10132),
.Y(net2292)
);

NAND2xp5_ASAP7_75t_R c2284(
.A(net2275),
.B(net2265),
.Y(net2293)
);

NAND2xp67_ASAP7_75t_R c2285(
.A(net2048),
.B(net2238),
.Y(net2294)
);

NOR2x1_ASAP7_75t_R c2286(
.A(net2288),
.B(net1398),
.Y(net2295)
);

NOR3xp33_ASAP7_75t_R c2287(
.A(net1381),
.B(net2275),
.C(net2292),
.Y(net2296)
);

NOR2x1p5_ASAP7_75t_R c2288(
.A(net2258),
.B(net2296),
.Y(net2297)
);

NOR2x2_ASAP7_75t_R c2289(
.A(net2297),
.B(net2272),
.Y(net2298)
);

NOR2xp33_ASAP7_75t_R c2290(
.A(net1331),
.B(net1282),
.Y(net2299)
);

AO221x2_ASAP7_75t_R c2291(
.A1(net2285),
.A2(net428),
.B1(net2131),
.B2(net2272),
.C(net10089),
.Y(net2300)
);

NOR2xp67_ASAP7_75t_R c2292(
.A(net2252),
.B(net10208),
.Y(net2301)
);

OR2x2_ASAP7_75t_R c2293(
.A(net2291),
.B(net9726),
.Y(net2302)
);

OR2x4_ASAP7_75t_R c2294(
.A(net2277),
.B(net1238),
.Y(net2303)
);

ICGx5p33DC_ASAP7_75t_R c2295(
.ENA(net2294),
.SE(net2249),
.CLK(clk),
.GCLK(net2304)
);

INVx4_ASAP7_75t_R c2296(
.A(net2303),
.Y(net2305)
);

OR2x6_ASAP7_75t_R c2297(
.A(net1038),
.B(net2274),
.Y(net2306)
);

INVx5_ASAP7_75t_R c2298(
.A(net10168),
.Y(net2307)
);

INVx6_ASAP7_75t_R c2299(
.A(net9985),
.Y(net2308)
);

XNOR2x1_ASAP7_75t_R c2300(
.B(net2306),
.A(net2292),
.Y(net2309)
);

XNOR2x2_ASAP7_75t_R c2301(
.A(net2274),
.B(net411),
.Y(net2310)
);

SDFLx4_ASAP7_75t_R c2302(
.D(net1367),
.SE(net407),
.SI(net2233),
.CLK(clk),
.QN(net2311)
);

INVx8_ASAP7_75t_R c2303(
.A(net2304),
.Y(net2312)
);

OA21x2_ASAP7_75t_R c2304(
.A1(net2310),
.A2(net2304),
.B(net2285),
.Y(net2313)
);

XNOR2xp5_ASAP7_75t_R c2305(
.A(net2289),
.B(net2256),
.Y(net2314)
);

XOR2x1_ASAP7_75t_R c2306(
.A(net1347),
.B(net2307),
.Y(net2315)
);

XOR2x2_ASAP7_75t_R c2307(
.A(net2299),
.B(net2293),
.Y(net2316)
);

XOR2xp5_ASAP7_75t_R c2308(
.A(net2255),
.B(net2274),
.Y(net2317)
);

DFFASRHQNx1_ASAP7_75t_R c2309(
.D(net2260),
.RESETN(net2316),
.SETN(net2317),
.CLK(clk),
.QN(net2318)
);

INVxp33_ASAP7_75t_R c2310(
.A(net10568),
.Y(net2319)
);

AND2x2_ASAP7_75t_R c2311(
.A(net2267),
.B(net2311),
.Y(net2320)
);

OR4x1_ASAP7_75t_R c2312(
.A(net2311),
.B(net1368),
.C(net2318),
.D(net2317),
.Y(net2321)
);

OAI222xp33_ASAP7_75t_R c2313(
.A1(net2145),
.A2(net2290),
.B1(net2320),
.B2(net2235),
.C1(net2316),
.C2(net2249),
.Y(net2322)
);

AND2x4_ASAP7_75t_R c2314(
.A(net1368),
.B(net2305),
.Y(net2323)
);

OR4x2_ASAP7_75t_R c2315(
.A(net2321),
.B(net2237),
.C(net2316),
.D(net9854),
.Y(net2324)
);

OAI21x1_ASAP7_75t_R c2316(
.A1(net2309),
.A2(net2314),
.B(net2318),
.Y(net2325)
);

OAI321xp33_ASAP7_75t_R c2317(
.A1(net2308),
.A2(net2318),
.A3(net2325),
.B1(net2311),
.B2(net2316),
.C(net1038),
.Y(net2326)
);

AO32x1_ASAP7_75t_R c2318(
.A1(net2316),
.A2(net2311),
.A3(net2315),
.B1(net2272),
.B2(net2317),
.Y(net2327)
);

OAI21xp33_ASAP7_75t_R c2319(
.A1(net1378),
.A2(net2316),
.B(net1250),
.Y(net2328)
);

A2O1A1Ixp33_ASAP7_75t_R c2320(
.A1(net2325),
.A2(net2307),
.B(net2316),
.C(net10211),
.Y(net2329)
);

AO32x2_ASAP7_75t_R c2321(
.A1(net2227),
.A2(net2321),
.A3(net2325),
.B1(net2316),
.B2(net2125),
.Y(net2330)
);

OAI33xp33_ASAP7_75t_R c2322(
.A1(net2233),
.A2(net2317),
.A3(net2325),
.B1(net2311),
.B2(net9844),
.B3(net10210),
.Y(net2331)
);

SDFHx1_ASAP7_75t_R c2323(
.D(net2319),
.SE(net2325),
.SI(net9764),
.CLK(clk),
.QN(net2332)
);

INVxp67_ASAP7_75t_R c2324(
.A(net1441),
.Y(net2333)
);

BUFx10_ASAP7_75t_R c2325(
.A(net10131),
.Y(net2334)
);

AND2x6_ASAP7_75t_R c2326(
.A(net2328),
.B(net2302),
.Y(net2335)
);

BUFx12_ASAP7_75t_R c2327(
.A(net510),
.Y(net2336)
);

BUFx12f_ASAP7_75t_R c2328(
.A(net2334),
.Y(net2337)
);

AO222x2_ASAP7_75t_R c2329(
.A1(net2250),
.A2(net1336),
.B1(net1458),
.B2(net1365),
.C1(net1446),
.C2(net9964),
.Y(net2338)
);

OAI21xp5_ASAP7_75t_R c2330(
.A1(net2238),
.A2(net2245),
.B(net1313),
.Y(net2339)
);

BUFx16f_ASAP7_75t_R c2331(
.A(net10112),
.Y(net2340)
);

BUFx24_ASAP7_75t_R c2332(
.A(net9682),
.Y(net2341)
);

BUFx2_ASAP7_75t_R c2333(
.A(net2320),
.Y(net2342)
);

HAxp5_ASAP7_75t_R c2334(
.A(net1462),
.B(net10082),
.CON(net2343)
);

NAND2x1_ASAP7_75t_R c2335(
.A(net2341),
.B(net2328),
.Y(net2344)
);

BUFx3_ASAP7_75t_R c2336(
.A(net9682),
.Y(net2345)
);

NAND2x1p5_ASAP7_75t_R c2337(
.A(net1433),
.B(net2338),
.Y(net2346)
);

NAND2x2_ASAP7_75t_R c2338(
.A(net2343),
.B(net10179),
.Y(net2347)
);

NAND2xp33_ASAP7_75t_R c2339(
.A(net1155),
.B(net1412),
.Y(net2348)
);

BUFx4_ASAP7_75t_R c2340(
.A(net2282),
.Y(net2349)
);

BUFx4f_ASAP7_75t_R c2341(
.A(net2345),
.Y(net2350)
);

NAND2xp5_ASAP7_75t_R c2342(
.A(net2349),
.B(net2034),
.Y(net2351)
);

NAND2xp67_ASAP7_75t_R c2343(
.A(net2230),
.B(net10209),
.Y(net2352)
);

BUFx5_ASAP7_75t_R c2344(
.A(net2351),
.Y(net2353)
);

NOR2x1_ASAP7_75t_R c2345(
.A(net2307),
.B(net2347),
.Y(net2354)
);

BUFx6f_ASAP7_75t_R c2346(
.A(net10563),
.Y(net2355)
);

NOR2x1p5_ASAP7_75t_R c2347(
.A(net2302),
.B(net2296),
.Y(net2356)
);

ICGx6p67DC_ASAP7_75t_R c2348(
.ENA(net2335),
.SE(net1457),
.CLK(clk),
.GCLK(net2357)
);

NOR2x2_ASAP7_75t_R c2349(
.A(net2340),
.B(net2357),
.Y(net2358)
);

ICGx8DC_ASAP7_75t_R c2350(
.ENA(net1485),
.SE(net2346),
.CLK(clk),
.GCLK(net2359)
);

NOR2xp33_ASAP7_75t_R c2351(
.A(net2336),
.B(net2340),
.Y(net2360)
);

NOR2xp67_ASAP7_75t_R c2352(
.A(net2360),
.B(net2352),
.Y(net2361)
);

OR3x1_ASAP7_75t_R c2353(
.A(net2357),
.B(net2199),
.C(net1458),
.Y(net2362)
);

BUFx8_ASAP7_75t_R c2354(
.A(net1451),
.Y(net2363)
);

OR2x2_ASAP7_75t_R c2355(
.A(net2342),
.B(net2360),
.Y(net2364)
);

CKINVDCx10_ASAP7_75t_R c2356(
.A(net2352),
.Y(net2365)
);

CKINVDCx11_ASAP7_75t_R c2357(
.A(net1464),
.Y(net2366)
);

SDFHx2_ASAP7_75t_R c2358(
.D(net1480),
.SE(net2351),
.SI(net1355),
.CLK(clk),
.QN(net2367)
);

AOI221x1_ASAP7_75t_R c2359(
.A1(net2242),
.A2(net2342),
.B1(net2361),
.B2(net2352),
.C(net1446),
.Y(net2368)
);

CKINVDCx12_ASAP7_75t_R c2360(
.A(net10024),
.Y(net2369)
);

OR2x4_ASAP7_75t_R c2361(
.A(net2338),
.B(net2355),
.Y(net2370)
);

ICGx1_ASAP7_75t_R c2362(
.ENA(net2355),
.SE(net2253),
.CLK(clk),
.GCLK(net2371)
);

OR2x6_ASAP7_75t_R c2363(
.A(net2296),
.B(net2328),
.Y(net2372)
);

XNOR2x1_ASAP7_75t_R c2364(
.B(net2348),
.A(net2367),
.Y(net2373)
);

CKINVDCx14_ASAP7_75t_R c2365(
.A(net9682),
.Y(net2374)
);

XNOR2x2_ASAP7_75t_R c2366(
.A(net2210),
.B(net2333),
.Y(net2375)
);

CKINVDCx16_ASAP7_75t_R c2367(
.A(net2295),
.Y(net2376)
);

XNOR2xp5_ASAP7_75t_R c2368(
.A(net2245),
.B(net10106),
.Y(net2377)
);

XOR2x1_ASAP7_75t_R c2369(
.A(net2358),
.B(net10196),
.Y(net2378)
);

OR3x2_ASAP7_75t_R c2370(
.A(net1401),
.B(net2357),
.C(net2250),
.Y(net2379)
);

XOR2x2_ASAP7_75t_R c2371(
.A(net2355),
.B(net327),
.Y(net2380)
);

XOR2xp5_ASAP7_75t_R c2372(
.A(net2368),
.B(net2296),
.Y(net2381)
);

CKINVDCx20_ASAP7_75t_R c2373(
.A(net2371),
.Y(net2382)
);

AND2x2_ASAP7_75t_R c2374(
.A(net1422),
.B(net2372),
.Y(net2383)
);

AND2x4_ASAP7_75t_R c2375(
.A(net2287),
.B(net2359),
.Y(net2384)
);

CKINVDCx5p33_ASAP7_75t_R c2376(
.A(net1473),
.Y(net2385)
);

AND2x6_ASAP7_75t_R c2377(
.A(net500),
.B(net10196),
.Y(net2386)
);

HAxp5_ASAP7_75t_R c2378(
.A(net1403),
.B(net2261),
.CON(net2388),
.SN(net2387)
);

CKINVDCx6p67_ASAP7_75t_R c2379(
.A(net2379),
.Y(net2389)
);

NAND2x1_ASAP7_75t_R c2380(
.A(net1478),
.B(net2352),
.Y(net2390)
);

CKINVDCx8_ASAP7_75t_R c2381(
.A(net10435),
.Y(net2391)
);

NAND2x1p5_ASAP7_75t_R c2382(
.A(net2374),
.B(net2371),
.Y(net2392)
);

AO33x2_ASAP7_75t_R c2383(
.A1(net2366),
.A2(net2362),
.A3(net2287),
.B1(net2355),
.B2(net1336),
.B3(net2358),
.Y(net2393)
);

OR3x4_ASAP7_75t_R c2384(
.A(net498),
.B(net2353),
.C(net1446),
.Y(net2394)
);

NAND2x2_ASAP7_75t_R c2385(
.A(net2388),
.B(net2386),
.Y(net2395)
);

CKINVDCx9p33_ASAP7_75t_R c2386(
.A(net9953),
.Y(net2396)
);

AND3x1_ASAP7_75t_R c2387(
.A(net2376),
.B(net2349),
.C(net2364),
.Y(net2397)
);

NAND2xp33_ASAP7_75t_R c2388(
.A(net2391),
.B(net2358),
.Y(net2398)
);

NAND2xp5_ASAP7_75t_R c2389(
.A(net2398),
.B(net2357),
.Y(net2399)
);

SDFHx3_ASAP7_75t_R c2390(
.D(net2397),
.SE(net2373),
.SI(net1473),
.CLK(clk),
.QN(net2400)
);

AND3x2_ASAP7_75t_R c2391(
.A(net2340),
.B(net2355),
.C(net2399),
.Y(net2401)
);

NAND2xp67_ASAP7_75t_R c2392(
.A(net2351),
.B(net2399),
.Y(net2402)
);

NOR2x1_ASAP7_75t_R c2393(
.A(net2389),
.B(net2396),
.Y(net2403)
);

NOR2x1p5_ASAP7_75t_R c2394(
.A(net2361),
.B(net445),
.Y(net2404)
);

NOR2x2_ASAP7_75t_R c2395(
.A(net2362),
.B(net2402),
.Y(net2405)
);

AOI221xp5_ASAP7_75t_R c2396(
.A1(net2356),
.A2(net2400),
.B1(net2401),
.B2(net1473),
.C(net2337),
.Y(net2406)
);

NOR2xp33_ASAP7_75t_R c2397(
.A(net2354),
.B(net2405),
.Y(net2407)
);

AOI222xp33_ASAP7_75t_R c2398(
.A1(net2384),
.A2(net2371),
.B1(net2399),
.B2(net1446),
.C1(net1313),
.C2(net10211),
.Y(net2408)
);

HB1xp67_ASAP7_75t_R c2399(
.A(net10112),
.Y(net2409)
);

NOR2xp67_ASAP7_75t_R c2400(
.A(net2409),
.B(net2355),
.Y(net2410)
);

AND3x4_ASAP7_75t_R c2401(
.A(net2403),
.B(net2191),
.C(net2337),
.Y(net2411)
);

AO21x1_ASAP7_75t_R c2402(
.A1(net2410),
.A2(net2367),
.B(net2372),
.Y(net2412)
);

HB2xp67_ASAP7_75t_R c2403(
.A(net9934),
.Y(net2413)
);

HB3xp67_ASAP7_75t_R c2404(
.A(net10522),
.Y(net2414)
);

SDFHx4_ASAP7_75t_R c2405(
.D(net2414),
.SE(net2395),
.SI(net2411),
.CLK(clk),
.QN(net2415)
);

AOI311xp33_ASAP7_75t_R c2406(
.A1(net2372),
.A2(net2394),
.A3(net1446),
.B(net2415),
.C(net2400),
.Y(net2416)
);

HB4xp67_ASAP7_75t_R c2407(
.A(net10413),
.Y(net2417)
);

INVx11_ASAP7_75t_R c2408(
.A(net1569),
.Y(net2418)
);

OR2x2_ASAP7_75t_R c2409(
.A(net1437),
.B(net2402),
.Y(net2419)
);

INVx13_ASAP7_75t_R c2410(
.A(net9130),
.Y(net2420)
);

INVx1_ASAP7_75t_R c2411(
.A(net1382),
.Y(net2421)
);

INVx2_ASAP7_75t_R c2412(
.A(net2419),
.Y(net2422)
);

INVx3_ASAP7_75t_R c2413(
.A(net9228),
.Y(net2423)
);

AO21x2_ASAP7_75t_R c2414(
.A1(net2034),
.A2(net2423),
.B(net1446),
.Y(net2424)
);

INVx4_ASAP7_75t_R c2415(
.A(net10470),
.Y(net2425)
);

INVx5_ASAP7_75t_R c2416(
.A(net1557),
.Y(net2426)
);

AOI21x1_ASAP7_75t_R c2417(
.A1(net2417),
.A2(net2425),
.B(net9854),
.Y(net2427)
);

INVx6_ASAP7_75t_R c2418(
.A(net568),
.Y(net2428)
);

INVx8_ASAP7_75t_R c2419(
.A(net1508),
.Y(net2429)
);

OR2x4_ASAP7_75t_R c2420(
.A(net2427),
.B(net1546),
.Y(net2430)
);

OR2x6_ASAP7_75t_R c2421(
.A(net1511),
.B(net2424),
.Y(net2431)
);

XNOR2x1_ASAP7_75t_R c2422(
.B(net2375),
.A(net10209),
.Y(net2432)
);

XNOR2x2_ASAP7_75t_R c2423(
.A(net2191),
.B(net2427),
.Y(net2433)
);

INVxp33_ASAP7_75t_R c2424(
.A(net9223),
.Y(net2434)
);

INVxp67_ASAP7_75t_R c2425(
.A(net2428),
.Y(net2435)
);

AND4x1_ASAP7_75t_R c2426(
.A(net2418),
.B(net1534),
.C(net1558),
.D(net2337),
.Y(net2436)
);

XNOR2xp5_ASAP7_75t_R c2427(
.A(net2435),
.B(net2425),
.Y(net2437)
);

XOR2x1_ASAP7_75t_R c2428(
.A(net2429),
.B(net1571),
.Y(net2438)
);

XOR2x2_ASAP7_75t_R c2429(
.A(net2401),
.B(net2382),
.Y(net2439)
);

XOR2xp5_ASAP7_75t_R c2430(
.A(net577),
.B(net2347),
.Y(net2440)
);

BUFx10_ASAP7_75t_R c2431(
.A(net626),
.Y(net2441)
);

BUFx12_ASAP7_75t_R c2432(
.A(net10485),
.Y(net2442)
);

AOI21xp33_ASAP7_75t_R c2433(
.A1(net2358),
.A2(net2433),
.B(net2333),
.Y(net2443)
);

BUFx12f_ASAP7_75t_R c2434(
.A(net10137),
.Y(net2444)
);

AND2x2_ASAP7_75t_R c2435(
.A(net2347),
.B(net2440),
.Y(net2445)
);

SDFLx1_ASAP7_75t_R c2436(
.D(net2433),
.SE(net2436),
.SI(net2437),
.CLK(clk),
.QN(net2446)
);

AND2x4_ASAP7_75t_R c2437(
.A(net588),
.B(net2423),
.Y(net2447)
);

AND2x6_ASAP7_75t_R c2438(
.A(net2442),
.B(net1521),
.Y(net2448)
);

BUFx16f_ASAP7_75t_R c2439(
.A(net10488),
.Y(net2449)
);

HAxp5_ASAP7_75t_R c2440(
.A(net2432),
.B(net2446),
.CON(net2451),
.SN(net2450)
);

NAND2x1_ASAP7_75t_R c2441(
.A(net2447),
.B(net2333),
.Y(net2452)
);

AOI21xp5_ASAP7_75t_R c2442(
.A1(net2448),
.A2(net2435),
.B(net2450),
.Y(net2453)
);

NAND2x1p5_ASAP7_75t_R c2443(
.A(net2350),
.B(net9644),
.Y(net2454)
);

NAND2x2_ASAP7_75t_R c2444(
.A(net2444),
.B(net2191),
.Y(net2455)
);

BUFx24_ASAP7_75t_R c2445(
.A(net9130),
.Y(net2456)
);

BUFx2_ASAP7_75t_R c2446(
.A(net10572),
.Y(net2457)
);

FAx1_ASAP7_75t_R c2447(
.A(net2423),
.B(net2417),
.CI(net1531),
.SN(net2458)
);

BUFx3_ASAP7_75t_R c2448(
.A(net10546),
.Y(net2459)
);

AND4x2_ASAP7_75t_R c2449(
.A(net1365),
.B(net2457),
.C(net2450),
.D(net2262),
.Y(net2460)
);

NAND2xp33_ASAP7_75t_R c2450(
.A(net2375),
.B(net1534),
.Y(net2461)
);

MAJIxp5_ASAP7_75t_R c2451(
.A(net2363),
.B(net2383),
.C(net9987),
.Y(net2462)
);

ICGx2_ASAP7_75t_R c2452(
.ENA(net2373),
.SE(net9934),
.CLK(clk),
.GCLK(net2463)
);

NAND2xp5_ASAP7_75t_R c2453(
.A(net2441),
.B(net445),
.Y(net2464)
);

NAND2xp67_ASAP7_75t_R c2454(
.A(net2446),
.B(net2401),
.Y(net2465)
);

NOR2x1_ASAP7_75t_R c2455(
.A(net2457),
.B(net2380),
.Y(net2466)
);

NOR2x1p5_ASAP7_75t_R c2456(
.A(net2451),
.B(net1572),
.Y(net2467)
);

NOR2x2_ASAP7_75t_R c2457(
.A(net2465),
.B(net2423),
.Y(net2468)
);

BUFx4_ASAP7_75t_R c2458(
.A(net2344),
.Y(net2469)
);

MAJx2_ASAP7_75t_R c2459(
.A(net2461),
.B(net2449),
.C(net2425),
.Y(net2470)
);

MAJx3_ASAP7_75t_R c2460(
.A(net2434),
.B(net2451),
.C(net1536),
.Y(net2471)
);

NOR2xp33_ASAP7_75t_R c2461(
.A(net1559),
.B(net1571),
.Y(net2472)
);

NOR2xp67_ASAP7_75t_R c2462(
.A(net2315),
.B(net1569),
.Y(net2473)
);

OR2x2_ASAP7_75t_R c2463(
.A(net1558),
.B(net1365),
.Y(net2474)
);

BUFx4f_ASAP7_75t_R c2464(
.A(net2473),
.Y(net2475)
);

OR2x4_ASAP7_75t_R c2465(
.A(net1545),
.B(net9970),
.Y(net2476)
);

OR2x6_ASAP7_75t_R c2466(
.A(net2468),
.B(net1561),
.Y(net2477)
);

BUFx5_ASAP7_75t_R c2467(
.A(net2454),
.Y(net2478)
);

XNOR2x1_ASAP7_75t_R c2468(
.B(net2417),
.A(net2451),
.Y(net2479)
);

BUFx6f_ASAP7_75t_R c2469(
.A(net9644),
.Y(net2480)
);

XNOR2x2_ASAP7_75t_R c2470(
.A(net2480),
.B(net609),
.Y(net2481)
);

XNOR2xp5_ASAP7_75t_R c2471(
.A(net2333),
.B(net1508),
.Y(net2482)
);

XOR2x1_ASAP7_75t_R c2472(
.A(net2481),
.B(net2479),
.Y(net2483)
);

XOR2x2_ASAP7_75t_R c2473(
.A(net338),
.B(net2262),
.Y(net2484)
);

XOR2xp5_ASAP7_75t_R c2474(
.A(net2382),
.B(net2446),
.Y(net2485)
);

AND2x2_ASAP7_75t_R c2475(
.A(net2476),
.B(net2473),
.Y(net2486)
);

AND2x4_ASAP7_75t_R c2476(
.A(net1545),
.B(net2449),
.Y(net2487)
);

AND2x6_ASAP7_75t_R c2477(
.A(net2485),
.B(net2473),
.Y(net2488)
);

AO211x2_ASAP7_75t_R c2478(
.A1(net622),
.A2(net2488),
.B(net2401),
.C(net1561),
.Y(net2489)
);

AO22x1_ASAP7_75t_R c2479(
.A1(net2482),
.A2(net1568),
.B1(net1561),
.B2(net10211),
.Y(net2490)
);

HAxp5_ASAP7_75t_R c2480(
.A(net2464),
.B(net2477),
.CON(net2492),
.SN(net2491)
);

BUFx8_ASAP7_75t_R c2481(
.A(net9285),
.Y(net2493)
);

NAND3x1_ASAP7_75t_R c2482(
.A(net2425),
.B(net2485),
.C(net2441),
.Y(net2494)
);

AO22x2_ASAP7_75t_R c2483(
.A1(net2490),
.A2(net2494),
.B1(net2463),
.B2(net10214),
.Y(net2495)
);

NAND2x1_ASAP7_75t_R c2484(
.A(net2467),
.B(net2477),
.Y(net2496)
);

AO31x2_ASAP7_75t_R c2485(
.A1(net2493),
.A2(net2479),
.A3(net2375),
.B(net626),
.Y(net2497)
);

NAND3x2_ASAP7_75t_R c2486(
.B(net2124),
.C(net2442),
.A(net2427),
.Y(net2498)
);

AOI211x1_ASAP7_75t_R c2487(
.A1(net2493),
.A2(net2487),
.B(net2498),
.C(net9813),
.Y(net2499)
);

NAND3xp33_ASAP7_75t_R c2488(
.A(net2484),
.B(net2492),
.C(net9970),
.Y(net2500)
);

NOR3x1_ASAP7_75t_R c2489(
.A(net2497),
.B(net2478),
.C(net9927),
.Y(net2501)
);

ICGx2p67DC_ASAP7_75t_R c2490(
.ENA(net716),
.SE(net2416),
.CLK(clk),
.GCLK(net2502)
);

NAND2x1p5_ASAP7_75t_R c2491(
.A(net1576),
.B(net1567),
.Y(net2503)
);

NAND2x2_ASAP7_75t_R c2492(
.A(net2430),
.B(net2424),
.Y(net2504)
);

CKINVDCx10_ASAP7_75t_R c2493(
.A(net2338),
.Y(net2505)
);

CKINVDCx11_ASAP7_75t_R c2494(
.A(net1618),
.Y(net2506)
);

NAND2xp33_ASAP7_75t_R c2495(
.A(net2477),
.B(net2426),
.Y(net2507)
);

NAND2xp5_ASAP7_75t_R c2496(
.A(net2369),
.B(net2392),
.Y(net2508)
);

CKINVDCx12_ASAP7_75t_R c2497(
.A(net9189),
.Y(net2509)
);

NOR3x2_ASAP7_75t_R c2498(
.B(net2507),
.C(net1526),
.A(net673),
.Y(net2510)
);

NAND2xp67_ASAP7_75t_R c2499(
.A(net2508),
.B(net1618),
.Y(net2511)
);

NOR2x1_ASAP7_75t_R c2500(
.A(net1569),
.B(net2511),
.Y(net2512)
);

NOR2x1p5_ASAP7_75t_R c2501(
.A(net2420),
.B(net2505),
.Y(net2513)
);

CKINVDCx14_ASAP7_75t_R c2502(
.A(net10124),
.Y(net2514)
);

NOR2x2_ASAP7_75t_R c2503(
.A(net2512),
.B(net2199),
.Y(net2515)
);

CKINVDCx16_ASAP7_75t_R c2504(
.A(net1312),
.Y(net2516)
);

CKINVDCx20_ASAP7_75t_R c2505(
.A(net1591),
.Y(net2517)
);

NOR2xp33_ASAP7_75t_R c2506(
.A(net1567),
.B(net673),
.Y(net2518)
);

NOR2xp67_ASAP7_75t_R c2507(
.A(net2199),
.B(net2477),
.Y(net2519)
);

OR2x2_ASAP7_75t_R c2508(
.A(net1626),
.B(net1652),
.Y(net2520)
);

NOR3xp33_ASAP7_75t_R c2509(
.A(net1455),
.B(net1561),
.C(net2353),
.Y(net2521)
);

CKINVDCx5p33_ASAP7_75t_R c2510(
.A(net10454),
.Y(net2522)
);

OR2x4_ASAP7_75t_R c2511(
.A(net2494),
.B(net9987),
.Y(net2523)
);

OR2x6_ASAP7_75t_R c2512(
.A(net2438),
.B(net2420),
.Y(net2524)
);

XNOR2x1_ASAP7_75t_R c2513(
.B(net651),
.A(net2494),
.Y(net2525)
);

XNOR2x2_ASAP7_75t_R c2514(
.A(net1610),
.B(net2358),
.Y(net2526)
);

XNOR2xp5_ASAP7_75t_R c2515(
.A(net2350),
.B(net2440),
.Y(net2527)
);

CKINVDCx6p67_ASAP7_75t_R c2516(
.A(net10003),
.Y(net2528)
);

CKINVDCx8_ASAP7_75t_R c2517(
.A(net10111),
.Y(net2529)
);

XOR2x1_ASAP7_75t_R c2518(
.A(net1620),
.B(net2517),
.Y(net2530)
);

XOR2x2_ASAP7_75t_R c2519(
.A(net1617),
.B(net1640),
.Y(net2531)
);

CKINVDCx9p33_ASAP7_75t_R c2520(
.A(net10469),
.Y(net2532)
);

OA21x2_ASAP7_75t_R c2521(
.A1(net2426),
.A2(net2506),
.B(net2515),
.Y(net2533)
);

XOR2xp5_ASAP7_75t_R c2522(
.A(net2522),
.B(net1621),
.Y(net2534)
);

AND2x2_ASAP7_75t_R c2523(
.A(net2524),
.B(net2438),
.Y(net2535)
);

HB1xp67_ASAP7_75t_R c2524(
.A(net9189),
.Y(net2536)
);

HB2xp67_ASAP7_75t_R c2525(
.A(net10378),
.Y(net2537)
);

HB3xp67_ASAP7_75t_R c2526(
.A(net2377),
.Y(net2538)
);

AND2x4_ASAP7_75t_R c2527(
.A(net1653),
.B(net2534),
.Y(net2539)
);

AOI211xp5_ASAP7_75t_R c2528(
.A1(net2516),
.A2(net1617),
.B(net2537),
.C(net2517),
.Y(net2540)
);

HB4xp67_ASAP7_75t_R c2529(
.A(net1614),
.Y(net2541)
);

AND2x6_ASAP7_75t_R c2530(
.A(net2541),
.B(net1655),
.Y(net2542)
);

HAxp5_ASAP7_75t_R c2531(
.A(net2534),
.B(net9679),
.CON(net2543)
);

INVx11_ASAP7_75t_R c2532(
.A(net10535),
.Y(net2544)
);

NAND2x1_ASAP7_75t_R c2533(
.A(net2543),
.B(net2337),
.Y(net2545)
);

AOI32xp33_ASAP7_75t_R c2534(
.A1(net2353),
.A2(net2538),
.A3(net2528),
.B1(net1653),
.B2(net1336),
.Y(net2546)
);

NAND2x1p5_ASAP7_75t_R c2535(
.A(net1546),
.B(net2424),
.Y(net2547)
);

OAI21x1_ASAP7_75t_R c2536(
.A1(net2504),
.A2(net2521),
.B(net651),
.Y(net2548)
);

NAND2x2_ASAP7_75t_R c2537(
.A(net671),
.B(net2508),
.Y(net2549)
);

NAND2xp33_ASAP7_75t_R c2538(
.A(net2545),
.B(net2538),
.Y(net2550)
);

NAND2xp5_ASAP7_75t_R c2539(
.A(net2392),
.B(net2538),
.Y(net2551)
);

NAND2xp67_ASAP7_75t_R c2540(
.A(net2532),
.B(net2526),
.Y(net2552)
);

ICGx3_ASAP7_75t_R c2541(
.ENA(net2528),
.SE(net1627),
.CLK(clk),
.GCLK(net2553)
);

OAI21xp33_ASAP7_75t_R c2542(
.A1(net2440),
.A2(net1614),
.B(net2553),
.Y(net2554)
);

ICGx4DC_ASAP7_75t_R c2543(
.ENA(net2515),
.SE(net671),
.CLK(clk),
.GCLK(net2555)
);

NOR2x1_ASAP7_75t_R c2544(
.A(net2290),
.B(net2547),
.Y(net2556)
);

NOR2x1p5_ASAP7_75t_R c2545(
.A(net1585),
.B(net2553),
.Y(net2557)
);

INVx13_ASAP7_75t_R c2546(
.A(net9994),
.Y(net2558)
);

NOR2x2_ASAP7_75t_R c2547(
.A(net2424),
.B(net2553),
.Y(net2559)
);

OAI21xp5_ASAP7_75t_R c2548(
.A1(net2559),
.A2(net2532),
.B(net2547),
.Y(net2560)
);

NOR2xp33_ASAP7_75t_R c2549(
.A(net1587),
.B(net2512),
.Y(net2561)
);

INVx1_ASAP7_75t_R c2550(
.A(net10056),
.Y(net2562)
);

NOR2xp67_ASAP7_75t_R c2551(
.A(net2527),
.B(net2554),
.Y(net2563)
);

OR2x2_ASAP7_75t_R c2552(
.A(net950),
.B(net2553),
.Y(net2564)
);

OR2x4_ASAP7_75t_R c2553(
.A(net1629),
.B(net2547),
.Y(net2565)
);

OR2x6_ASAP7_75t_R c2554(
.A(net1634),
.B(net2539),
.Y(net2566)
);

XNOR2x1_ASAP7_75t_R c2555(
.B(net2555),
.A(net10002),
.Y(net2567)
);

XNOR2x2_ASAP7_75t_R c2556(
.A(net2514),
.B(net1625),
.Y(net2568)
);

SDFLx2_ASAP7_75t_R c2557(
.D(net2540),
.SE(net2522),
.SI(net10107),
.CLK(clk),
.QN(net2569)
);

INVx2_ASAP7_75t_R c2558(
.A(net10541),
.Y(net2570)
);

XNOR2xp5_ASAP7_75t_R c2559(
.A(net2536),
.B(net2557),
.Y(net2571)
);

NAND5xp2_ASAP7_75t_R c2560(
.A(net2570),
.B(net2571),
.C(net2358),
.D(net665),
.E(net2538),
.Y(net2572)
);

INVx3_ASAP7_75t_R c2561(
.A(net10469),
.Y(net2573)
);

OR3x1_ASAP7_75t_R c2562(
.A(net2573),
.B(net598),
.C(net10034),
.Y(net2574)
);

XOR2x1_ASAP7_75t_R c2563(
.A(net2563),
.B(net2562),
.Y(net2575)
);

OR3x2_ASAP7_75t_R c2564(
.A(net2575),
.B(net2574),
.C(net2558),
.Y(net2576)
);

AOI321xp33_ASAP7_75t_R c2565(
.A1(net2526),
.A2(net2571),
.A3(net722),
.B1(net1526),
.B2(net2563),
.C(net2574),
.Y(net2577)
);

OR3x4_ASAP7_75t_R c2566(
.A(net2445),
.B(net2569),
.C(net10034),
.Y(net2578)
);

AND3x1_ASAP7_75t_R c2567(
.A(net2550),
.B(net2577),
.C(net10162),
.Y(net2579)
);

XOR2x2_ASAP7_75t_R c2568(
.A(net2553),
.B(net2522),
.Y(net2580)
);

AND3x2_ASAP7_75t_R c2569(
.A(net2573),
.B(net2574),
.C(net1651),
.Y(net2581)
);

NOR5xp2_ASAP7_75t_R c2570(
.A(net2574),
.B(net2558),
.C(net2517),
.D(net9842),
.E(net10162),
.Y(net2582)
);

XOR2xp5_ASAP7_75t_R c2571(
.A(net2577),
.B(net2551),
.Y(net2583)
);

INVx4_ASAP7_75t_R c2572(
.A(net10561),
.Y(net2584)
);

INVx5_ASAP7_75t_R c2573(
.A(net10097),
.Y(net2585)
);

AND2x2_ASAP7_75t_R c2574(
.A(net1718),
.B(net2506),
.Y(net2586)
);

INVx6_ASAP7_75t_R c2575(
.A(net10153),
.Y(net2587)
);

INVx8_ASAP7_75t_R c2576(
.A(net777),
.Y(net2588)
);

INVxp33_ASAP7_75t_R c2577(
.A(net2546),
.Y(net2589)
);

INVxp67_ASAP7_75t_R c2578(
.A(net2520),
.Y(net2590)
);

AOI22x1_ASAP7_75t_R c2579(
.A1(net1719),
.A2(net1730),
.B1(net2449),
.B2(net2558),
.Y(net2591)
);

AND2x4_ASAP7_75t_R c2580(
.A(net1740),
.B(net2539),
.Y(net2592)
);

AND2x6_ASAP7_75t_R c2581(
.A(net2572),
.B(net1718),
.Y(net2593)
);

BUFx10_ASAP7_75t_R c2582(
.A(net1729),
.Y(net2594)
);

AND3x4_ASAP7_75t_R c2583(
.A(net2586),
.B(net1625),
.C(net1730),
.Y(net2595)
);

BUFx12_ASAP7_75t_R c2584(
.A(net10558),
.Y(net2596)
);

BUFx12f_ASAP7_75t_R c2585(
.A(net9153),
.Y(net2597)
);

BUFx16f_ASAP7_75t_R c2586(
.A(net2509),
.Y(net2598)
);

BUFx24_ASAP7_75t_R c2587(
.A(net10508),
.Y(net2599)
);

HAxp5_ASAP7_75t_R c2588(
.A(net1432),
.B(net10213),
.CON(net2601),
.SN(net2600)
);

NAND2x1_ASAP7_75t_R c2589(
.A(net2558),
.B(net1672),
.Y(net2602)
);

BUFx2_ASAP7_75t_R c2590(
.A(net2592),
.Y(net2603)
);

BUFx3_ASAP7_75t_R c2591(
.A(net2557),
.Y(net2604)
);

BUFx4_ASAP7_75t_R c2592(
.A(net2567),
.Y(net2605)
);

AO21x1_ASAP7_75t_R c2593(
.A1(net2588),
.A2(net2590),
.B(net2605),
.Y(net2606)
);

BUFx4f_ASAP7_75t_R c2594(
.A(net2506),
.Y(net2607)
);

BUFx5_ASAP7_75t_R c2595(
.A(net10117),
.Y(net2608)
);

NAND2x1p5_ASAP7_75t_R c2596(
.A(net2448),
.B(net10200),
.Y(net2609)
);

NAND2x2_ASAP7_75t_R c2597(
.A(net2608),
.B(net2558),
.Y(net2610)
);

BUFx6f_ASAP7_75t_R c2598(
.A(net10087),
.Y(net2611)
);

BUFx8_ASAP7_75t_R c2599(
.A(net9679),
.Y(net2612)
);

NAND2xp33_ASAP7_75t_R c2600(
.A(net2602),
.B(net1718),
.Y(net2613)
);

AO21x2_ASAP7_75t_R c2601(
.A1(net2416),
.A2(net2555),
.B(net2589),
.Y(net2614)
);

NAND2xp5_ASAP7_75t_R c2602(
.A(net2596),
.B(net1522),
.Y(net2615)
);

NAND2xp67_ASAP7_75t_R c2603(
.A(net1658),
.B(net775),
.Y(net2616)
);

NOR2x1_ASAP7_75t_R c2604(
.A(net798),
.B(net2448),
.Y(net2617)
);

NOR2x1p5_ASAP7_75t_R c2605(
.A(net1721),
.B(net2617),
.Y(net2618)
);

CKINVDCx10_ASAP7_75t_R c2606(
.A(net1710),
.Y(net2619)
);

NOR2x2_ASAP7_75t_R c2607(
.A(net2612),
.B(net1694),
.Y(net2620)
);

NOR2xp33_ASAP7_75t_R c2608(
.A(net1672),
.B(net2574),
.Y(net2621)
);

NOR2xp67_ASAP7_75t_R c2609(
.A(net2586),
.B(net10102),
.Y(net2622)
);

OR2x2_ASAP7_75t_R c2610(
.A(net2580),
.B(net1611),
.Y(net2623)
);

CKINVDCx11_ASAP7_75t_R c2611(
.A(net9153),
.Y(net2624)
);

OR2x4_ASAP7_75t_R c2612(
.A(net2623),
.B(net665),
.Y(net2625)
);

CKINVDCx12_ASAP7_75t_R c2613(
.A(net9952),
.Y(net2626)
);

OR2x6_ASAP7_75t_R c2614(
.A(net2611),
.B(net2449),
.Y(net2627)
);

XNOR2x1_ASAP7_75t_R c2615(
.B(net2505),
.A(net1658),
.Y(net2628)
);

XNOR2x2_ASAP7_75t_R c2616(
.A(net2624),
.B(net10105),
.Y(net2629)
);

ICGx4_ASAP7_75t_R c2617(
.ENA(net1738),
.SE(net2624),
.CLK(clk),
.GCLK(net2630)
);

XNOR2xp5_ASAP7_75t_R c2618(
.A(net2587),
.B(net2624),
.Y(net2631)
);

XOR2x1_ASAP7_75t_R c2619(
.A(net2534),
.B(net2631),
.Y(net2632)
);

XOR2x2_ASAP7_75t_R c2620(
.A(net1735),
.B(net598),
.Y(net2633)
);

XOR2xp5_ASAP7_75t_R c2621(
.A(net2603),
.B(net2618),
.Y(net2634)
);

AND2x2_ASAP7_75t_R c2622(
.A(net2618),
.B(net2539),
.Y(net2635)
);

AOI22xp33_ASAP7_75t_R c2623(
.A1(net2604),
.A2(net2617),
.B1(net2629),
.B2(net2619),
.Y(net2636)
);

AND2x4_ASAP7_75t_R c2624(
.A(net2635),
.B(net2634),
.Y(net2637)
);

AND2x6_ASAP7_75t_R c2625(
.A(net2523),
.B(net1729),
.Y(net2638)
);

OA221x2_ASAP7_75t_R c2626(
.A1(net2633),
.A2(net2593),
.B1(net1718),
.B2(net1664),
.C(net2615),
.Y(net2639)
);

AOI21x1_ASAP7_75t_R c2627(
.A1(net2593),
.A2(net2624),
.B(net10022),
.Y(net2640)
);

HAxp5_ASAP7_75t_R c2628(
.A(net2627),
.B(net2634),
.CON(net2641)
);

NAND2x1_ASAP7_75t_R c2629(
.A(net1712),
.B(net2558),
.Y(net2642)
);

NAND2x1p5_ASAP7_75t_R c2630(
.A(net2609),
.B(net2607),
.Y(net2643)
);

AOI21xp33_ASAP7_75t_R c2631(
.A1(net2640),
.A2(net2624),
.B(net2588),
.Y(net2644)
);

SDFLx3_ASAP7_75t_R c2632(
.D(net2641),
.SE(net2637),
.SI(net2643),
.CLK(clk),
.QN(net2645)
);

NAND2x2_ASAP7_75t_R c2633(
.A(net2606),
.B(net2605),
.Y(net2646)
);

NAND2xp33_ASAP7_75t_R c2634(
.A(net2646),
.B(net2645),
.Y(net2647)
);

NAND2xp5_ASAP7_75t_R c2635(
.A(net2607),
.B(net2625),
.Y(net2648)
);

CKINVDCx14_ASAP7_75t_R c2636(
.A(net9952),
.Y(net2649)
);

NAND2xp67_ASAP7_75t_R c2637(
.A(net2622),
.B(net10105),
.Y(net2650)
);

AOI22xp5_ASAP7_75t_R c2638(
.A1(net2650),
.A2(net2630),
.B1(net2638),
.B2(net2624),
.Y(net2651)
);

AOI21xp5_ASAP7_75t_R c2639(
.A1(net2647),
.A2(net2380),
.B(net2448),
.Y(net2652)
);

NOR2x1_ASAP7_75t_R c2640(
.A(net2245),
.B(net10215),
.Y(net2653)
);

AOI31xp33_ASAP7_75t_R c2641(
.A1(net2564),
.A2(net2539),
.A3(net2620),
.B(net10215),
.Y(net2654)
);

NOR2x1p5_ASAP7_75t_R c2642(
.A(net2622),
.B(net2654),
.Y(net2655)
);

OAI221xp5_ASAP7_75t_R c2643(
.A1(net673),
.A2(net2463),
.B1(net2619),
.B2(net2615),
.C(net10102),
.Y(net2656)
);

NOR2x2_ASAP7_75t_R c2644(
.A(net2593),
.B(net2650),
.Y(net2657)
);

NOR2xp33_ASAP7_75t_R c2645(
.A(net2656),
.B(net1592),
.Y(net2658)
);

ICGx5_ASAP7_75t_R c2646(
.ENA(net2631),
.SE(net2657),
.CLK(clk),
.GCLK(net2659)
);

CKINVDCx16_ASAP7_75t_R c2647(
.A(net10102),
.Y(net2660)
);

NOR2xp67_ASAP7_75t_R c2648(
.A(net2660),
.B(net10215),
.Y(net2661)
);

OAI311xp33_ASAP7_75t_R c2649(
.A1(net2652),
.A2(net2650),
.A3(net2646),
.B1(net2661),
.C1(net2615),
.Y(net2662)
);

OR2x2_ASAP7_75t_R c2650(
.A(net2648),
.B(net2618),
.Y(net2663)
);

OR2x4_ASAP7_75t_R c2651(
.A(net2655),
.B(net2657),
.Y(net2664)
);

OR2x6_ASAP7_75t_R c2652(
.A(net2639),
.B(net2659),
.Y(net2665)
);

XNOR2x1_ASAP7_75t_R c2653(
.B(net2625),
.A(net2659),
.Y(net2666)
);

XNOR2x2_ASAP7_75t_R c2654(
.A(net1490),
.B(net9897),
.Y(net2667)
);

XNOR2xp5_ASAP7_75t_R c2655(
.A(net2659),
.B(net10105),
.Y(net2668)
);

XOR2x1_ASAP7_75t_R c2656(
.A(net1815),
.B(net1777),
.Y(net2669)
);

XOR2x2_ASAP7_75t_R c2657(
.A(net1680),
.B(net1757),
.Y(net2670)
);

XOR2xp5_ASAP7_75t_R c2658(
.A(net1750),
.B(net2634),
.Y(net2671)
);

FAx1_ASAP7_75t_R c2659(
.A(net2599),
.B(net1803),
.CI(net1671),
.SN(net2672)
);

OAI32xp33_ASAP7_75t_R c2660(
.A1(net1640),
.A2(net897),
.A3(net824),
.B1(net2617),
.B2(net749),
.Y(net2673)
);

ICGx5p33DC_ASAP7_75t_R c2661(
.ENA(net2491),
.SE(net9782),
.CLK(clk),
.GCLK(net2674)
);

AND2x2_ASAP7_75t_R c2662(
.A(net893),
.B(net2670),
.Y(net2675)
);

CKINVDCx20_ASAP7_75t_R c2663(
.A(net10343),
.Y(net2676)
);

AND2x4_ASAP7_75t_R c2664(
.A(net1788),
.B(net2674),
.Y(net2677)
);

AND2x6_ASAP7_75t_R c2665(
.A(net2675),
.B(net1787),
.Y(net2678)
);

HAxp5_ASAP7_75t_R c2666(
.A(net1540),
.B(net860),
.CON(net2680),
.SN(net2679)
);

ICGx6p67DC_ASAP7_75t_R c2667(
.ENA(net743),
.SE(net2492),
.CLK(clk),
.GCLK(net2681)
);

ICGx8DC_ASAP7_75t_R c2668(
.ENA(net2680),
.SE(net1763),
.CLK(clk),
.GCLK(net2682)
);

NAND2x1_ASAP7_75t_R c2669(
.A(net842),
.B(net849),
.Y(net2683)
);

NAND2x1p5_ASAP7_75t_R c2670(
.A(net2262),
.B(net860),
.Y(net2684)
);

NAND2x2_ASAP7_75t_R c2671(
.A(net897),
.B(net1774),
.Y(net2685)
);

NAND2xp33_ASAP7_75t_R c2672(
.A(net2659),
.B(net1727),
.Y(net2686)
);

NAND2xp5_ASAP7_75t_R c2673(
.A(net892),
.B(net860),
.Y(net2687)
);

NAND2xp67_ASAP7_75t_R c2674(
.A(net765),
.B(net1777),
.Y(net2688)
);

MAJIxp5_ASAP7_75t_R c2675(
.A(net665),
.B(net2649),
.C(net873),
.Y(net2689)
);

NOR2x1_ASAP7_75t_R c2676(
.A(net861),
.B(net2679),
.Y(net2690)
);

NOR2x1p5_ASAP7_75t_R c2677(
.A(net871),
.B(net2674),
.Y(net2691)
);

NOR2x2_ASAP7_75t_R c2678(
.A(net2674),
.B(net2686),
.Y(net2692)
);

NOR2xp33_ASAP7_75t_R c2679(
.A(net1592),
.B(net2675),
.Y(net2693)
);

NOR2xp67_ASAP7_75t_R c2680(
.A(net2632),
.B(net893),
.Y(net2694)
);

OR2x2_ASAP7_75t_R c2681(
.A(net1797),
.B(net2673),
.Y(net2695)
);

CKINVDCx5p33_ASAP7_75t_R c2682(
.A(net2621),
.Y(net2696)
);

OR2x4_ASAP7_75t_R c2683(
.A(net2521),
.B(net2673),
.Y(net2697)
);

CKINVDCx6p67_ASAP7_75t_R c2684(
.A(net10538),
.Y(net2698)
);

OR2x6_ASAP7_75t_R c2685(
.A(net1780),
.B(net2689),
.Y(net2699)
);

XNOR2x1_ASAP7_75t_R c2686(
.B(net2684),
.A(net10200),
.Y(net2700)
);

XNOR2x2_ASAP7_75t_R c2687(
.A(net2676),
.B(net10215),
.Y(net2701)
);

XNOR2xp5_ASAP7_75t_R c2688(
.A(net836),
.B(net9651),
.Y(net2702)
);

SDFLx4_ASAP7_75t_R c2689(
.D(net2685),
.SE(net1785),
.SI(net1788),
.CLK(clk),
.QN(net2703)
);

XOR2x1_ASAP7_75t_R c2690(
.A(net891),
.B(net1727),
.Y(net2704)
);

MAJx2_ASAP7_75t_R c2691(
.A(net2653),
.B(net1759),
.C(net10201),
.Y(net2705)
);

XOR2x2_ASAP7_75t_R c2692(
.A(net1803),
.B(net2705),
.Y(net2706)
);

XOR2xp5_ASAP7_75t_R c2693(
.A(net860),
.B(net2698),
.Y(net2707)
);

AND2x2_ASAP7_75t_R c2694(
.A(net2701),
.B(net2699),
.Y(net2708)
);

AND2x4_ASAP7_75t_R c2695(
.A(net885),
.B(net2705),
.Y(net2709)
);

OR5x1_ASAP7_75t_R c2696(
.A(net2653),
.B(net1784),
.C(net1671),
.D(net2699),
.E(net2707),
.Y(net2710)
);

DFFASRHQNx1_ASAP7_75t_R c2697(
.D(net2710),
.RESETN(net2687),
.SETN(net885),
.CLK(clk),
.QN(net2711)
);

AND2x6_ASAP7_75t_R c2698(
.A(net1760),
.B(net2711),
.Y(net2712)
);

HAxp5_ASAP7_75t_R c2699(
.A(net787),
.B(net1787),
.CON(net2714),
.SN(net2713)
);

NAND2x1_ASAP7_75t_R c2700(
.A(net2706),
.B(net842),
.Y(net2715)
);

MAJx3_ASAP7_75t_R c2701(
.A(net2634),
.B(net2696),
.C(net10200),
.Y(net2716)
);

NAND2x1p5_ASAP7_75t_R c2702(
.A(net868),
.B(net1680),
.Y(net2717)
);

OR5x2_ASAP7_75t_R c2703(
.A(net881),
.B(net2492),
.C(net2645),
.D(net2675),
.E(net1787),
.Y(net2718)
);

ICGx1_ASAP7_75t_R c2704(
.ENA(net2555),
.SE(net2716),
.CLK(clk),
.GCLK(net2719)
);

NAND3x1_ASAP7_75t_R c2705(
.A(net2694),
.B(net2719),
.C(net824),
.Y(net2720)
);

AOI31xp67_ASAP7_75t_R c2706(
.A1(net2717),
.A2(net1807),
.A3(net892),
.B(net2708),
.Y(net2721)
);

NAND2x2_ASAP7_75t_R c2707(
.A(net2698),
.B(net9920),
.Y(net2722)
);

CKINVDCx8_ASAP7_75t_R c2708(
.A(net10364),
.Y(net2723)
);

CKINVDCx9p33_ASAP7_75t_R c2709(
.A(net10536),
.Y(net2724)
);

ICGx2_ASAP7_75t_R c2710(
.ENA(net2690),
.SE(net2709),
.CLK(clk),
.GCLK(net2725)
);

NAND2xp33_ASAP7_75t_R c2711(
.A(net2666),
.B(net2722),
.Y(net2726)
);

NAND4xp25_ASAP7_75t_R c2712(
.A(net2725),
.B(net2705),
.C(net1807),
.D(net10211),
.Y(net2727)
);

NAND2xp5_ASAP7_75t_R c2713(
.A(net2624),
.B(net2726),
.Y(net2728)
);

ICGx2p67DC_ASAP7_75t_R c2714(
.ENA(net1763),
.SE(net2727),
.CLK(clk),
.GCLK(net2729)
);

NAND3x2_ASAP7_75t_R c2715(
.B(net810),
.C(net1823),
.A(net2706),
.Y(net2730)
);

NAND3xp33_ASAP7_75t_R c2716(
.A(net749),
.B(net2722),
.C(net873),
.Y(net2731)
);

NAND2xp67_ASAP7_75t_R c2717(
.A(net1621),
.B(net2713),
.Y(net2732)
);

NOR3x1_ASAP7_75t_R c2718(
.A(net2692),
.B(net1822),
.C(net2599),
.Y(net2733)
);

HB1xp67_ASAP7_75t_R c2719(
.A(net10483),
.Y(net2734)
);

NOR2x1_ASAP7_75t_R c2720(
.A(net2649),
.B(net2724),
.Y(net2735)
);

NOR2x1p5_ASAP7_75t_R c2721(
.A(net1521),
.B(net2677),
.Y(net2736)
);

NAND4xp75_ASAP7_75t_R c2722(
.A(net2730),
.B(net2732),
.C(net2719),
.D(net849),
.Y(net2737)
);

NOR2x2_ASAP7_75t_R c2723(
.A(net2449),
.B(net2683),
.Y(net2738)
);

NOR2xp33_ASAP7_75t_R c2724(
.A(net2738),
.B(net2463),
.Y(net2739)
);

SDFHx1_ASAP7_75t_R c2725(
.D(net2739),
.SE(net2732),
.SI(net10217),
.CLK(clk),
.QN(net2740)
);

A2O1A1O1Ixp25_ASAP7_75t_R c2726(
.A1(net2697),
.A2(net885),
.B(net2735),
.C(net2740),
.D(net2719),
.Y(net2741)
);

HB2xp67_ASAP7_75t_R c2727(
.A(net10343),
.Y(net2742)
);

NOR3x2_ASAP7_75t_R c2728(
.B(net2715),
.C(net2702),
.A(net1621),
.Y(net2743)
);

NOR2xp67_ASAP7_75t_R c2729(
.A(net2740),
.B(net9801),
.Y(net2744)
);

OR2x2_ASAP7_75t_R c2730(
.A(net2688),
.B(net2743),
.Y(net2745)
);

NOR3xp33_ASAP7_75t_R c2731(
.A(net1671),
.B(net2740),
.C(net2733),
.Y(net2746)
);

OR2x4_ASAP7_75t_R c2732(
.A(net1572),
.B(net9801),
.Y(net2747)
);

SDFHx2_ASAP7_75t_R c2733(
.D(net2727),
.SE(net1798),
.SI(net2747),
.CLK(clk),
.QN(net2748)
);

NOR4xp25_ASAP7_75t_R c2734(
.A(net1757),
.B(net2732),
.C(net2747),
.D(net10216),
.Y(net2749)
);

OA21x2_ASAP7_75t_R c2735(
.A1(net2722),
.A2(net2735),
.B(net2744),
.Y(net2750)
);

OAI21x1_ASAP7_75t_R c2736(
.A1(net2750),
.A2(net2742),
.B(net2748),
.Y(net2751)
);

OAI21xp33_ASAP7_75t_R c2737(
.A1(net2751),
.A2(net2746),
.B(net2621),
.Y(net2752)
);

AOI33xp33_ASAP7_75t_R c2738(
.A1(net1727),
.A2(net2751),
.A3(net2747),
.B1(net824),
.B2(net2732),
.B3(net9651),
.Y(net2753)
);

HB3xp67_ASAP7_75t_R c2739(
.A(net1900),
.Y(net2754)
);

HB4xp67_ASAP7_75t_R c2740(
.A(net1879),
.Y(net2755)
);

INVx11_ASAP7_75t_R c2741(
.A(net922),
.Y(net2756)
);

ICGx3_ASAP7_75t_R c2742(
.ENA(in24),
.SE(net982),
.CLK(clk),
.GCLK(net2757)
);

INVx13_ASAP7_75t_R c2743(
.A(net2756),
.Y(net2758)
);

INVx1_ASAP7_75t_R c2744(
.A(net1842),
.Y(net2759)
);

INVx2_ASAP7_75t_R c2745(
.A(net2755),
.Y(net2760)
);

INVx3_ASAP7_75t_R c2746(
.A(net2754),
.Y(net2761)
);

OR2x6_ASAP7_75t_R c2747(
.A(net919),
.B(net10204),
.Y(net2762)
);

XNOR2x1_ASAP7_75t_R c2748(
.B(net927),
.A(net2756),
.Y(net2763)
);

XNOR2x2_ASAP7_75t_R c2749(
.A(net1835),
.B(in7),
.Y(net2764)
);

XNOR2xp5_ASAP7_75t_R c2750(
.A(net1865),
.B(net1897),
.Y(net2765)
);

INVx4_ASAP7_75t_R c2751(
.A(net15),
.Y(net2766)
);

INVx5_ASAP7_75t_R c2752(
.A(net928),
.Y(net2767)
);

XOR2x1_ASAP7_75t_R c2753(
.A(net922),
.B(net1886),
.Y(net2768)
);

OAI21xp5_ASAP7_75t_R c2754(
.A1(net2761),
.A2(net2762),
.B(net2767),
.Y(net2769)
);

XOR2x2_ASAP7_75t_R c2755(
.A(net2764),
.B(net1845),
.Y(net2770)
);

INVx6_ASAP7_75t_R c2756(
.A(net2764),
.Y(net2771)
);

INVx8_ASAP7_75t_R c2757(
.A(net1857),
.Y(net2772)
);

XOR2xp5_ASAP7_75t_R c2758(
.A(net2767),
.B(net10204),
.Y(net2773)
);

AND2x2_ASAP7_75t_R c2759(
.A(net2773),
.B(net2755),
.Y(net2774)
);

INVxp33_ASAP7_75t_R c2760(
.A(net964),
.Y(net2775)
);

OR3x1_ASAP7_75t_R c2761(
.A(net2772),
.B(net1842),
.C(net959),
.Y(net2776)
);

INVxp67_ASAP7_75t_R c2762(
.A(net1886),
.Y(net2777)
);

BUFx10_ASAP7_75t_R c2763(
.A(net1884),
.Y(net2778)
);

OR3x2_ASAP7_75t_R c2764(
.A(net2768),
.B(net2775),
.C(net34),
.Y(net2779)
);

AND2x4_ASAP7_75t_R c2765(
.A(net1900),
.B(net2773),
.Y(net2780)
);

BUFx12_ASAP7_75t_R c2766(
.A(net9095),
.Y(net2781)
);

ICGx4DC_ASAP7_75t_R c2767(
.ENA(net2776),
.SE(net1848),
.CLK(clk),
.GCLK(net2782)
);

BUFx12f_ASAP7_75t_R c2768(
.A(net9095),
.Y(net2783)
);

OR3x4_ASAP7_75t_R c2769(
.A(net2783),
.B(net2770),
.C(in24),
.Y(net2784)
);

BUFx16f_ASAP7_75t_R c2770(
.A(net1842),
.Y(net2785)
);

AND2x6_ASAP7_75t_R c2771(
.A(net2767),
.B(net1875),
.Y(net2786)
);

AND3x1_ASAP7_75t_R c2772(
.A(net2784),
.B(net2771),
.C(net2777),
.Y(net2787)
);

HAxp5_ASAP7_75t_R c2773(
.A(net2763),
.B(net2757),
.CON(net2788)
);

BUFx24_ASAP7_75t_R c2774(
.A(net2762),
.Y(net2789)
);

NAND2x1_ASAP7_75t_R c2775(
.A(net1842),
.B(net9744),
.Y(net2790)
);

NAND2x1p5_ASAP7_75t_R c2776(
.A(net2788),
.B(net947),
.Y(net2791)
);

BUFx2_ASAP7_75t_R c2777(
.A(net2781),
.Y(net2792)
);

NAND2x2_ASAP7_75t_R c2778(
.A(net1897),
.B(net1857),
.Y(net2793)
);

BUFx3_ASAP7_75t_R c2779(
.A(net964),
.Y(net2794)
);

NAND2xp33_ASAP7_75t_R c2780(
.A(net2771),
.B(net2760),
.Y(net2795)
);

NAND2xp5_ASAP7_75t_R c2781(
.A(net2759),
.B(net2770),
.Y(net2796)
);

BUFx4_ASAP7_75t_R c2782(
.A(net2765),
.Y(net2797)
);

BUFx4f_ASAP7_75t_R c2783(
.A(net2773),
.Y(net2798)
);

NAND2xp67_ASAP7_75t_R c2784(
.A(net2778),
.B(net2781),
.Y(net2799)
);

NOR2x1_ASAP7_75t_R c2785(
.A(net2795),
.B(net2783),
.Y(net2800)
);

NOR2x1p5_ASAP7_75t_R c2786(
.A(net2800),
.B(net9717),
.Y(net2801)
);

NOR2x2_ASAP7_75t_R c2787(
.A(net1845),
.B(net9717),
.Y(net2802)
);

BUFx5_ASAP7_75t_R c2788(
.A(net2769),
.Y(net2803)
);

NOR2xp33_ASAP7_75t_R c2789(
.A(net2802),
.B(net2796),
.Y(net2804)
);

BUFx6f_ASAP7_75t_R c2790(
.A(net2801),
.Y(net2805)
);

SDFHx3_ASAP7_75t_R c2791(
.D(net2789),
.SE(net2780),
.SI(net2782),
.CLK(clk),
.QN(net2806)
);

NOR2xp67_ASAP7_75t_R c2792(
.A(net2797),
.B(net2786),
.Y(net2807)
);

AND3x2_ASAP7_75t_R c2793(
.A(net2790),
.B(net2781),
.C(net2783),
.Y(net2808)
);

ICGx4_ASAP7_75t_R c2794(
.ENA(net2798),
.SE(net2782),
.CLK(clk),
.GCLK(net2809)
);

SDFHx4_ASAP7_75t_R c2795(
.D(net2806),
.SE(net2797),
.SI(net2807),
.CLK(clk),
.QN(net2810)
);

OR2x2_ASAP7_75t_R c2796(
.A(net1831),
.B(net2805),
.Y(net2811)
);

SDFLx1_ASAP7_75t_R c2797(
.D(net2770),
.SE(net2803),
.SI(net2763),
.CLK(clk),
.QN(net2812)
);

OR2x4_ASAP7_75t_R c2798(
.A(net2786),
.B(net2776),
.Y(net2813)
);

SDFLx2_ASAP7_75t_R c2799(
.D(net2800),
.SE(net2810),
.SI(net2807),
.CLK(clk),
.QN(net2814)
);

ICGx5_ASAP7_75t_R c2800(
.ENA(net2808),
.SE(net2813),
.CLK(clk),
.GCLK(net2815)
);

OR2x6_ASAP7_75t_R c2801(
.A(net2796),
.B(net919),
.Y(net2816)
);

SDFLx3_ASAP7_75t_R c2802(
.D(net2782),
.SE(net2803),
.SI(net2806),
.CLK(clk),
.QN(net2817)
);

AND3x4_ASAP7_75t_R c2803(
.A(net2793),
.B(net2815),
.C(net2781),
.Y(net2818)
);

AO21x1_ASAP7_75t_R c2804(
.A1(net2805),
.A2(net2761),
.B(net2814),
.Y(net2819)
);

AO21x2_ASAP7_75t_R c2805(
.A1(net2787),
.A2(net2794),
.B(net2768),
.Y(net2820)
);

AOI21x1_ASAP7_75t_R c2806(
.A1(net2775),
.A2(net2814),
.B(net2817),
.Y(net2821)
);

XNOR2x1_ASAP7_75t_R c2807(
.B(net2772),
.A(net2765),
.Y(net2822)
);

NOR4xp75_ASAP7_75t_R c2808(
.A(net2814),
.B(net2818),
.C(net2766),
.D(net1827),
.Y(net2823)
);

SDFLx4_ASAP7_75t_R c2809(
.D(net2803),
.SE(net2818),
.SI(net2820),
.CLK(clk),
.QN(net2824)
);

XNOR2x2_ASAP7_75t_R c2810(
.A(net2785),
.B(net2820),
.Y(net2825)
);

XNOR2xp5_ASAP7_75t_R c2811(
.A(net2818),
.B(net1886),
.Y(net2826)
);

AOI21xp33_ASAP7_75t_R c2812(
.A1(net2817),
.A2(net2824),
.B(net2821),
.Y(net2827)
);

XOR2x1_ASAP7_75t_R c2813(
.A(net2820),
.B(net2822),
.Y(net2828)
);

XOR2x2_ASAP7_75t_R c2814(
.A(net2784),
.B(net2821),
.Y(net2829)
);

ICGx5p33DC_ASAP7_75t_R c2815(
.ENA(net982),
.SE(net1883),
.CLK(clk),
.GCLK(net2830)
);

XOR2xp5_ASAP7_75t_R c2816(
.A(net2821),
.B(net2826),
.Y(net2831)
);

DFFASRHQNx1_ASAP7_75t_R c2817(
.D(net1879),
.RESETN(net2808),
.SETN(net2807),
.CLK(clk),
.QN(net2832)
);

AND2x2_ASAP7_75t_R c2818(
.A(net2824),
.B(net2826),
.Y(net2833)
);

AND5x1_ASAP7_75t_R c2819(
.A(net2789),
.B(net2781),
.C(net2820),
.D(net2811),
.E(net2829),
.Y(net2834)
);

AND5x2_ASAP7_75t_R c2820(
.A(net2833),
.B(net2820),
.C(net2830),
.D(net2829),
.E(net2823),
.Y(net2835)
);

AND2x4_ASAP7_75t_R c2821(
.A(net2833),
.B(net9717),
.Y(net2836)
);

AND2x6_ASAP7_75t_R c2822(
.A(net2766),
.B(net1972),
.Y(net2837)
);

BUFx8_ASAP7_75t_R c2823(
.A(net996),
.Y(net2838)
);

CKINVDCx10_ASAP7_75t_R c2824(
.A(net2816),
.Y(net2839)
);

ICGx6p67DC_ASAP7_75t_R c2825(
.ENA(net1059),
.SE(net1915),
.CLK(clk),
.GCLK(net2840)
);

CKINVDCx11_ASAP7_75t_R c2826(
.A(net1022),
.Y(net2841)
);

CKINVDCx12_ASAP7_75t_R c2827(
.A(net2830),
.Y(net2842)
);

HAxp5_ASAP7_75t_R c2828(
.A(net1875),
.B(net2791),
.CON(net2843)
);

CKINVDCx14_ASAP7_75t_R c2829(
.A(net1926),
.Y(net2844)
);

CKINVDCx16_ASAP7_75t_R c2830(
.A(net1008),
.Y(net2845)
);

CKINVDCx20_ASAP7_75t_R c2831(
.A(net9107),
.Y(net2846)
);

CKINVDCx5p33_ASAP7_75t_R c2832(
.A(net10219),
.Y(net2847)
);

CKINVDCx6p67_ASAP7_75t_R c2833(
.A(net9889),
.Y(net2848)
);

CKINVDCx8_ASAP7_75t_R c2834(
.A(net2809),
.Y(net2849)
);

CKINVDCx9p33_ASAP7_75t_R c2835(
.A(net9702),
.Y(net2850)
);

HB1xp67_ASAP7_75t_R c2836(
.A(net1919),
.Y(net2851)
);

HB2xp67_ASAP7_75t_R c2837(
.A(net2794),
.Y(net2852)
);

HB3xp67_ASAP7_75t_R c2838(
.A(net2841),
.Y(net2853)
);

HB4xp67_ASAP7_75t_R c2839(
.A(net2851),
.Y(net2854)
);

INVx11_ASAP7_75t_R c2840(
.A(net2850),
.Y(net2855)
);

NAND2x1_ASAP7_75t_R c2841(
.A(net2827),
.B(net2839),
.Y(net2856)
);

INVx13_ASAP7_75t_R c2842(
.A(net2832),
.Y(net2857)
);

INVx1_ASAP7_75t_R c2843(
.A(net9107),
.Y(net2858)
);

INVx2_ASAP7_75t_R c2844(
.A(net30),
.Y(net2859)
);

INVx3_ASAP7_75t_R c2845(
.A(net2853),
.Y(net2860)
);

NAND2x1p5_ASAP7_75t_R c2846(
.A(net2791),
.B(net2853),
.Y(net2861)
);

NAND2x2_ASAP7_75t_R c2847(
.A(net2844),
.B(net950),
.Y(net2862)
);

INVx4_ASAP7_75t_R c2848(
.A(net2815),
.Y(net2863)
);

NAND2xp33_ASAP7_75t_R c2849(
.A(net1966),
.B(net2853),
.Y(net2864)
);

AOI21xp5_ASAP7_75t_R c2850(
.A1(net1952),
.A2(net2859),
.B(net2832),
.Y(net2865)
);

FAx1_ASAP7_75t_R c2851(
.A(net2760),
.B(net2840),
.CI(net2859),
.SN(net2867),
.CON(net2866)
);

MAJIxp5_ASAP7_75t_R c2852(
.A(net2854),
.B(net1988),
.C(net1911),
.Y(net2868)
);

NAND2xp5_ASAP7_75t_R c2853(
.A(net2863),
.B(net1861),
.Y(net2869)
);

NAND2xp67_ASAP7_75t_R c2854(
.A(net2850),
.B(net1963),
.Y(net2870)
);

INVx5_ASAP7_75t_R c2855(
.A(net2859),
.Y(net2871)
);

NOR2x1_ASAP7_75t_R c2856(
.A(net1986),
.B(net2811),
.Y(net2872)
);

INVx6_ASAP7_75t_R c2857(
.A(net1981),
.Y(net2873)
);

INVx8_ASAP7_75t_R c2858(
.A(net2852),
.Y(net2874)
);

INVxp33_ASAP7_75t_R c2859(
.A(net9257),
.Y(net2875)
);

INVxp67_ASAP7_75t_R c2860(
.A(net2845),
.Y(net2876)
);

MAJx2_ASAP7_75t_R c2861(
.A(net2871),
.B(net2853),
.C(net1844),
.Y(net2877)
);

BUFx10_ASAP7_75t_R c2862(
.A(net9244),
.Y(net2878)
);

NOR2x1p5_ASAP7_75t_R c2863(
.A(net2876),
.B(net79),
.Y(net2879)
);

BUFx12_ASAP7_75t_R c2864(
.A(net2862),
.Y(net2880)
);

BUFx12f_ASAP7_75t_R c2865(
.A(net2879),
.Y(net2881)
);

BUFx16f_ASAP7_75t_R c2866(
.A(net2858),
.Y(net2882)
);

ICGx8DC_ASAP7_75t_R c2867(
.ENA(net2869),
.SE(net2807),
.CLK(clk),
.GCLK(net2883)
);

ICGx1_ASAP7_75t_R c2868(
.ENA(net2864),
.SE(net1971),
.CLK(clk),
.GCLK(net2884)
);

NOR2x2_ASAP7_75t_R c2869(
.A(net2880),
.B(net2875),
.Y(net2885)
);

NOR2xp33_ASAP7_75t_R c2870(
.A(net2857),
.B(net9725),
.Y(net2886)
);

NOR2xp67_ASAP7_75t_R c2871(
.A(net2838),
.B(net2875),
.Y(net2887)
);

OR2x2_ASAP7_75t_R c2872(
.A(net2873),
.B(net2884),
.Y(net2888)
);

BUFx24_ASAP7_75t_R c2873(
.A(net2881),
.Y(net2889)
);

BUFx2_ASAP7_75t_R c2874(
.A(net9238),
.Y(net2890)
);

OR2x4_ASAP7_75t_R c2875(
.A(net2868),
.B(net2857),
.Y(net2891)
);

BUFx3_ASAP7_75t_R c2876(
.A(net1865),
.Y(net2892)
);

BUFx4_ASAP7_75t_R c2877(
.A(net2889),
.Y(net2893)
);

OR2x6_ASAP7_75t_R c2878(
.A(net2849),
.B(net2880),
.Y(net2894)
);

O2A1O1Ixp33_ASAP7_75t_R c2879(
.A1(net2886),
.A2(net1941),
.B(net2877),
.C(net10189),
.Y(net2895)
);

XNOR2x1_ASAP7_75t_R c2880(
.B(net2846),
.A(net2809),
.Y(net2896)
);

XNOR2x2_ASAP7_75t_R c2881(
.A(net2888),
.B(net2875),
.Y(net2897)
);

XNOR2xp5_ASAP7_75t_R c2882(
.A(net945),
.B(net1961),
.Y(net2898)
);

BUFx4f_ASAP7_75t_R c2883(
.A(net10422),
.Y(net2899)
);

XOR2x1_ASAP7_75t_R c2884(
.A(net2892),
.B(net10220),
.Y(net2900)
);

XOR2x2_ASAP7_75t_R c2885(
.A(net2839),
.B(net2900),
.Y(net2901)
);

MAJx3_ASAP7_75t_R c2886(
.A(net2901),
.B(net2890),
.C(net1972),
.Y(net2902)
);

XOR2xp5_ASAP7_75t_R c2887(
.A(net2878),
.B(net2900),
.Y(net2903)
);

NAND3x1_ASAP7_75t_R c2888(
.A(net2837),
.B(net2870),
.C(net2875),
.Y(net2904)
);

AND2x2_ASAP7_75t_R c2889(
.A(net1883),
.B(net2903),
.Y(net2905)
);

NAND3x2_ASAP7_75t_R c2890(
.B(net2904),
.C(net2874),
.A(net2757),
.Y(net2906)
);

AND2x4_ASAP7_75t_R c2891(
.A(net2890),
.B(net2905),
.Y(net2907)
);

ICGx2_ASAP7_75t_R c2892(
.ENA(net2840),
.SE(net1976),
.CLK(clk),
.GCLK(net2908)
);

AND2x6_ASAP7_75t_R c2893(
.A(net1941),
.B(net2897),
.Y(net2909)
);

NAND3xp33_ASAP7_75t_R c2894(
.A(net2902),
.B(net1927),
.C(net2903),
.Y(net2910)
);

HAxp5_ASAP7_75t_R c2895(
.A(net2875),
.B(net9821),
.CON(net2911)
);

SDFHx1_ASAP7_75t_R c2896(
.D(net1936),
.SE(net2907),
.SI(net2810),
.CLK(clk),
.QN(net2912)
);

NAND2x1_ASAP7_75t_R c2897(
.A(net2910),
.B(net2866),
.Y(net2913)
);

NAND2x1p5_ASAP7_75t_R c2898(
.A(net2912),
.B(net2908),
.Y(net2914)
);

NOR3x1_ASAP7_75t_R c2899(
.A(net1931),
.B(net2908),
.C(net2914),
.Y(net2915)
);

O2A1O1Ixp5_ASAP7_75t_R c2900(
.A1(net2915),
.A2(net2860),
.B(net2908),
.C(net2914),
.Y(net2916)
);

NAND2x2_ASAP7_75t_R c2901(
.A(net2912),
.B(net9756),
.Y(net2917)
);

OA222x2_ASAP7_75t_R c2902(
.A1(net2914),
.A2(net2908),
.B1(net2884),
.B2(net2907),
.C1(net2899),
.C2(net2842),
.Y(net2918)
);

OA33x2_ASAP7_75t_R c2903(
.A1(net2911),
.A2(net2855),
.A3(net2909),
.B1(net1898),
.B2(net2918),
.B3(net10220),
.Y(net2919)
);

NOR3x2_ASAP7_75t_R c2904(
.B(net2894),
.C(net2914),
.A(net2918),
.Y(net2920)
);

NAND2xp33_ASAP7_75t_R c2905(
.A(net2883),
.B(net2918),
.Y(net2921)
);

OA211x2_ASAP7_75t_R c2906(
.A1(net2061),
.A2(net2836),
.B(net2071),
.C(net34),
.Y(net2922)
);

BUFx5_ASAP7_75t_R c2907(
.A(net1994),
.Y(net2923)
);

BUFx6f_ASAP7_75t_R c2908(
.A(net2006),
.Y(net2924)
);

BUFx8_ASAP7_75t_R c2909(
.A(net9174),
.Y(net2925)
);

NAND2xp5_ASAP7_75t_R c2910(
.A(net2893),
.B(net2755),
.Y(net2926)
);

CKINVDCx10_ASAP7_75t_R c2911(
.A(net9174),
.Y(net2927)
);

CKINVDCx11_ASAP7_75t_R c2912(
.A(net2924),
.Y(net2928)
);

NAND2xp67_ASAP7_75t_R c2913(
.A(net2923),
.B(net2014),
.Y(net2929)
);

NOR3xp33_ASAP7_75t_R c2914(
.A(net2055),
.B(net1102),
.C(net2857),
.Y(net2930)
);

CKINVDCx12_ASAP7_75t_R c2915(
.A(net2018),
.Y(net2931)
);

CKINVDCx14_ASAP7_75t_R c2916(
.A(net1947),
.Y(net2932)
);

NOR2x1_ASAP7_75t_R c2917(
.A(net2932),
.B(net1138),
.Y(net2933)
);

NOR2x1p5_ASAP7_75t_R c2918(
.A(net2931),
.B(net1947),
.Y(net2934)
);

NOR2x2_ASAP7_75t_R c2919(
.A(net2928),
.B(net2903),
.Y(net2935)
);

CKINVDCx16_ASAP7_75t_R c2920(
.A(net9907),
.Y(net2936)
);

CKINVDCx20_ASAP7_75t_R c2921(
.A(net10071),
.Y(net2937)
);

CKINVDCx5p33_ASAP7_75t_R c2922(
.A(net2935),
.Y(net2938)
);

NOR2xp33_ASAP7_75t_R c2923(
.A(net2062),
.B(net1980),
.Y(net2939)
);

CKINVDCx6p67_ASAP7_75t_R c2924(
.A(net1972),
.Y(net2940)
);

CKINVDCx8_ASAP7_75t_R c2925(
.A(net2075),
.Y(net2941)
);

CKINVDCx9p33_ASAP7_75t_R c2926(
.A(net10108),
.Y(net2942)
);

NOR2xp67_ASAP7_75t_R c2927(
.A(net2929),
.B(net2938),
.Y(net2943)
);

OR2x2_ASAP7_75t_R c2928(
.A(net2907),
.B(net2062),
.Y(net2944)
);

HB1xp67_ASAP7_75t_R c2929(
.A(net10013),
.Y(net2945)
);

HB2xp67_ASAP7_75t_R c2930(
.A(net2934),
.Y(net2946)
);

HB3xp67_ASAP7_75t_R c2931(
.A(net2944),
.Y(net2947)
);

HB4xp67_ASAP7_75t_R c2932(
.A(net2937),
.Y(net2948)
);

INVx11_ASAP7_75t_R c2933(
.A(net2945),
.Y(net2949)
);

OR2x4_ASAP7_75t_R c2934(
.A(net2949),
.B(net2909),
.Y(net2950)
);

INVx13_ASAP7_75t_R c2935(
.A(net2943),
.Y(net2951)
);

OR2x6_ASAP7_75t_R c2936(
.A(net1102),
.B(net2075),
.Y(net2952)
);

INVx1_ASAP7_75t_R c2937(
.A(net10136),
.Y(net2953)
);

XNOR2x1_ASAP7_75t_R c2938(
.B(net1945),
.A(net1898),
.Y(net2954)
);

INVx2_ASAP7_75t_R c2939(
.A(net9752),
.Y(net2955)
);

XNOR2x2_ASAP7_75t_R c2940(
.A(net1114),
.B(net2946),
.Y(net2956)
);

INVx3_ASAP7_75t_R c2941(
.A(net2936),
.Y(net2957)
);

XNOR2xp5_ASAP7_75t_R c2942(
.A(net2758),
.B(net10047),
.Y(net2958)
);

XOR2x1_ASAP7_75t_R c2943(
.A(net2955),
.B(net2883),
.Y(net2959)
);

INVx4_ASAP7_75t_R c2944(
.A(net1898),
.Y(net2960)
);

INVx5_ASAP7_75t_R c2945(
.A(net9202),
.Y(net2961)
);

XOR2x2_ASAP7_75t_R c2946(
.A(net2957),
.B(net2954),
.Y(net2962)
);

XOR2xp5_ASAP7_75t_R c2947(
.A(net2925),
.B(net2071),
.Y(net2963)
);

AND2x2_ASAP7_75t_R c2948(
.A(net2903),
.B(net2962),
.Y(net2964)
);

AND2x4_ASAP7_75t_R c2949(
.A(net2836),
.B(net2963),
.Y(net2965)
);

INVx6_ASAP7_75t_R c2950(
.A(net2964),
.Y(net2966)
);

INVx8_ASAP7_75t_R c2951(
.A(net2887),
.Y(net2967)
);

AND2x6_ASAP7_75t_R c2952(
.A(net2807),
.B(net180),
.Y(net2968)
);

INVxp33_ASAP7_75t_R c2953(
.A(net9992),
.Y(net2969)
);

INVxp67_ASAP7_75t_R c2954(
.A(net9950),
.Y(net2970)
);

BUFx10_ASAP7_75t_R c2955(
.A(net9926),
.Y(net2971)
);

OA21x2_ASAP7_75t_R c2956(
.A1(net2961),
.A2(net2960),
.B(net2962),
.Y(net2972)
);

HAxp5_ASAP7_75t_R c2957(
.A(net2972),
.B(net2971),
.CON(net2974),
.SN(net2973)
);

NAND2x1_ASAP7_75t_R c2958(
.A(net2962),
.B(net2955),
.Y(net2975)
);

OAI21x1_ASAP7_75t_R c2959(
.A1(net2969),
.A2(net2947),
.B(net2909),
.Y(net2976)
);

NAND2x1p5_ASAP7_75t_R c2960(
.A(net2971),
.B(net2938),
.Y(net2977)
);

BUFx12_ASAP7_75t_R c2961(
.A(net1052),
.Y(net2978)
);

NAND2x2_ASAP7_75t_R c2962(
.A(net2970),
.B(net2961),
.Y(net2979)
);

NAND2xp33_ASAP7_75t_R c2963(
.A(net2940),
.B(net2947),
.Y(net2980)
);

NAND2xp5_ASAP7_75t_R c2964(
.A(net2959),
.B(net2963),
.Y(net2981)
);

NAND2xp67_ASAP7_75t_R c2965(
.A(net1005),
.B(net2963),
.Y(net2982)
);

NOR2x1_ASAP7_75t_R c2966(
.A(net2965),
.B(net2959),
.Y(net2983)
);

BUFx12f_ASAP7_75t_R c2967(
.A(net9980),
.Y(net2984)
);

BUFx16f_ASAP7_75t_R c2968(
.A(net10422),
.Y(net2985)
);

OAI21xp33_ASAP7_75t_R c2969(
.A1(net2939),
.A2(net2907),
.B(net2942),
.Y(net2986)
);

OAI21xp5_ASAP7_75t_R c2970(
.A1(net2857),
.A2(net2985),
.B(net2861),
.Y(net2987)
);

NOR2x1p5_ASAP7_75t_R c2971(
.A(net1093),
.B(net2052),
.Y(net2988)
);

AO221x1_ASAP7_75t_R c2972(
.A1(net2988),
.A2(net2075),
.B1(net2836),
.B2(net2036),
.C(net2963),
.Y(net2989)
);

NOR2x2_ASAP7_75t_R c2973(
.A(net2947),
.B(net2989),
.Y(net2990)
);

BUFx24_ASAP7_75t_R c2974(
.A(net2983),
.Y(net2991)
);

NOR2xp33_ASAP7_75t_R c2975(
.A(net2975),
.B(net2985),
.Y(net2992)
);

OA22x2_ASAP7_75t_R c2976(
.A1(net178),
.A2(net2989),
.B1(net2991),
.B2(net2071),
.Y(net2993)
);

NOR2xp67_ASAP7_75t_R c2977(
.A(net2982),
.B(net2954),
.Y(net2994)
);

OR2x2_ASAP7_75t_R c2978(
.A(net2976),
.B(net2990),
.Y(net2995)
);

BUFx2_ASAP7_75t_R c2979(
.A(net10064),
.Y(net2996)
);

SDFHx2_ASAP7_75t_R c2980(
.D(net2909),
.SE(net2974),
.SI(net2991),
.CLK(clk),
.QN(net2997)
);

OR3x1_ASAP7_75t_R c2981(
.A(net2980),
.B(net2984),
.C(net2997),
.Y(net2998)
);

OR3x2_ASAP7_75t_R c2982(
.A(net2986),
.B(net1827),
.C(net2980),
.Y(net2999)
);

AO221x2_ASAP7_75t_R c2983(
.A1(net2950),
.A2(net2967),
.B1(net2977),
.B2(net2962),
.C(net2942),
.Y(net3000)
);

AO32x1_ASAP7_75t_R c2984(
.A1(net2941),
.A2(net2967),
.A3(net2996),
.B1(net2917),
.B2(net2942),
.Y(net3001)
);

OR3x4_ASAP7_75t_R c2985(
.A(net2978),
.B(net2985),
.C(net2971),
.Y(net3002)
);

SDFHx3_ASAP7_75t_R c2986(
.D(net2995),
.SE(net2962),
.SI(net9725),
.CLK(clk),
.QN(net3003)
);

AND3x1_ASAP7_75t_R c2987(
.A(net2994),
.B(net2983),
.C(net3003),
.Y(net3004)
);

OR2x4_ASAP7_75t_R c2988(
.A(net2151),
.B(net2060),
.Y(net3005)
);

OR2x6_ASAP7_75t_R c2989(
.A(net2948),
.B(net2117),
.Y(net3006)
);

BUFx3_ASAP7_75t_R c2990(
.A(net2905),
.Y(net3007)
);

BUFx4_ASAP7_75t_R c2991(
.A(net2089),
.Y(net3008)
);

XNOR2x1_ASAP7_75t_R c2992(
.B(net1984),
.A(net2128),
.Y(net3009)
);

XNOR2x2_ASAP7_75t_R c2993(
.A(net259),
.B(net1172),
.Y(net3010)
);

XNOR2xp5_ASAP7_75t_R c2994(
.A(net3008),
.B(net2081),
.Y(net3011)
);

BUFx4f_ASAP7_75t_R c2995(
.A(net2979),
.Y(net3012)
);

BUFx5_ASAP7_75t_R c2996(
.A(net2977),
.Y(net3013)
);

XOR2x1_ASAP7_75t_R c2997(
.A(net1229),
.B(net10047),
.Y(net3014)
);

BUFx6f_ASAP7_75t_R c2998(
.A(net10482),
.Y(net3015)
);

BUFx8_ASAP7_75t_R c2999(
.A(net10083),
.Y(net3016)
);

AND3x2_ASAP7_75t_R c3000(
.A(net3013),
.B(net2977),
.C(net3003),
.Y(net3017)
);

XOR2x2_ASAP7_75t_R c3001(
.A(net2060),
.B(net2905),
.Y(net3018)
);

AND3x4_ASAP7_75t_R c3002(
.A(net3005),
.B(net1172),
.C(net10088),
.Y(net3019)
);

XOR2xp5_ASAP7_75t_R c3003(
.A(net1833),
.B(net2997),
.Y(net3020)
);

AND2x2_ASAP7_75t_R c3004(
.A(net2084),
.B(net79),
.Y(net3021)
);

AND2x4_ASAP7_75t_R c3005(
.A(net994),
.B(net3004),
.Y(net3022)
);

AND2x6_ASAP7_75t_R c3006(
.A(net3018),
.B(net3015),
.Y(net3023)
);

CKINVDCx10_ASAP7_75t_R c3007(
.A(net10083),
.Y(net3024)
);

HAxp5_ASAP7_75t_R c3008(
.A(net2088),
.B(net1163),
.CON(net3026),
.SN(net3025)
);

CKINVDCx11_ASAP7_75t_R c3009(
.A(net3009),
.Y(net3027)
);

NAND2x1_ASAP7_75t_R c3010(
.A(net2981),
.B(net1922),
.Y(net3028)
);

NAND2x1p5_ASAP7_75t_R c3011(
.A(net2128),
.B(net10063),
.Y(net3029)
);

NAND2x2_ASAP7_75t_R c3012(
.A(net2144),
.B(net2089),
.Y(net3030)
);

NAND2xp33_ASAP7_75t_R c3013(
.A(net3030),
.B(net1229),
.Y(net3031)
);

CKINVDCx12_ASAP7_75t_R c3014(
.A(net10508),
.Y(net3032)
);

ICGx2p67DC_ASAP7_75t_R c3015(
.ENA(net2992),
.SE(net3032),
.CLK(clk),
.GCLK(net3033)
);

CKINVDCx14_ASAP7_75t_R c3016(
.A(net10569),
.Y(net3034)
);

NAND2xp5_ASAP7_75t_R c3017(
.A(net2128),
.B(net2997),
.Y(net3035)
);

CKINVDCx16_ASAP7_75t_R c3018(
.A(net3016),
.Y(net3036)
);

CKINVDCx20_ASAP7_75t_R c3019(
.A(net10091),
.Y(net3037)
);

AO21x1_ASAP7_75t_R c3020(
.A1(net958),
.A2(net2993),
.B(net3001),
.Y(net3038)
);

SDFHx4_ASAP7_75t_R c3021(
.D(net2989),
.SE(net2131),
.SI(net9996),
.CLK(clk),
.QN(net3039)
);

NAND2xp67_ASAP7_75t_R c3022(
.A(net1140),
.B(net272),
.Y(net3040)
);

CKINVDCx5p33_ASAP7_75t_R c3023(
.A(net9315),
.Y(net3041)
);

CKINVDCx6p67_ASAP7_75t_R c3024(
.A(net9973),
.Y(net3042)
);

NOR2x1_ASAP7_75t_R c3025(
.A(net3014),
.B(net10063),
.Y(net3043)
);

CKINVDCx8_ASAP7_75t_R c3026(
.A(net10063),
.Y(net3044)
);

AO32x2_ASAP7_75t_R c3027(
.A1(net3036),
.A2(net3035),
.A3(net2997),
.B1(net2842),
.B2(net2084),
.Y(net3045)
);

NOR2x1p5_ASAP7_75t_R c3028(
.A(net2081),
.B(net3045),
.Y(net3046)
);

NOR2x2_ASAP7_75t_R c3029(
.A(net3021),
.B(net3042),
.Y(net3047)
);

NOR2xp33_ASAP7_75t_R c3030(
.A(net3037),
.B(net2917),
.Y(net3048)
);

NOR2xp67_ASAP7_75t_R c3031(
.A(net2755),
.B(net2991),
.Y(net3049)
);

AOI221x1_ASAP7_75t_R c3032(
.A1(net3023),
.A2(net270),
.B1(net3049),
.B2(net3034),
.C(net10088),
.Y(net3050)
);

CKINVDCx9p33_ASAP7_75t_R c3033(
.A(net180),
.Y(net3051)
);

OR2x2_ASAP7_75t_R c3034(
.A(net2161),
.B(net3048),
.Y(net3052)
);

OR2x4_ASAP7_75t_R c3035(
.A(net3035),
.B(net3032),
.Y(net3053)
);

OR2x6_ASAP7_75t_R c3036(
.A(net2917),
.B(net10221),
.Y(net3054)
);

AO21x2_ASAP7_75t_R c3037(
.A1(net3044),
.A2(net2036),
.B(net1915),
.Y(net3055)
);

XNOR2x1_ASAP7_75t_R c3038(
.B(net3045),
.A(net3039),
.Y(net3056)
);

AOI21x1_ASAP7_75t_R c3039(
.A1(net3052),
.A2(net2128),
.B(net3054),
.Y(net3057)
);

XNOR2x2_ASAP7_75t_R c3040(
.A(net3051),
.B(net10221),
.Y(net3058)
);

XNOR2xp5_ASAP7_75t_R c3041(
.A(net3028),
.B(net3033),
.Y(net3059)
);

AOI21xp33_ASAP7_75t_R c3042(
.A1(net3055),
.A2(net3049),
.B(net3034),
.Y(net3060)
);

XOR2x1_ASAP7_75t_R c3043(
.A(net3006),
.B(net1195),
.Y(net3061)
);

XOR2x2_ASAP7_75t_R c3044(
.A(net2960),
.B(net3051),
.Y(net3062)
);

XOR2xp5_ASAP7_75t_R c3045(
.A(net3047),
.B(net3004),
.Y(net3063)
);

AND2x2_ASAP7_75t_R c3046(
.A(net3053),
.B(net3044),
.Y(net3064)
);

AOI21xp5_ASAP7_75t_R c3047(
.A1(net3061),
.A2(net3039),
.B(net10028),
.Y(net3065)
);

FAx1_ASAP7_75t_R c3048(
.A(net1927),
.B(net3045),
.CI(net2981),
.SN(net3067),
.CON(net3066)
);

MAJIxp5_ASAP7_75t_R c3049(
.A(net1195),
.B(net3062),
.C(net3034),
.Y(net3068)
);

AND2x4_ASAP7_75t_R c3050(
.A(net3029),
.B(net3067),
.Y(net3069)
);

HB1xp67_ASAP7_75t_R c3051(
.A(net9961),
.Y(net3070)
);

MAJx2_ASAP7_75t_R c3052(
.A(net3065),
.B(net1963),
.C(net3070),
.Y(net3071)
);

AOI221xp5_ASAP7_75t_R c3053(
.A1(net3042),
.A2(net3049),
.B1(net2905),
.B2(net2084),
.C(net2963),
.Y(net3072)
);

SDFLx1_ASAP7_75t_R c3054(
.D(net3058),
.SE(net3069),
.SI(net10222),
.CLK(clk),
.QN(net3073)
);

MAJx3_ASAP7_75t_R c3055(
.A(net3020),
.B(net3051),
.C(net3006),
.Y(net3074)
);

AND2x6_ASAP7_75t_R c3056(
.A(net3064),
.B(net3048),
.Y(net3075)
);

AOI311xp33_ASAP7_75t_R c3057(
.A1(net3074),
.A2(net3061),
.A3(net3059),
.B(net3015),
.C(net3073),
.Y(net3076)
);

HAxp5_ASAP7_75t_R c3058(
.A(net3059),
.B(net10028),
.CON(net3078),
.SN(net3077)
);

NAND3x1_ASAP7_75t_R c3059(
.A(net3071),
.B(net3010),
.C(net2917),
.Y(net3079)
);

SDFLx2_ASAP7_75t_R c3060(
.D(net3068),
.SE(net3078),
.SI(net2755),
.CLK(clk),
.QN(net3080)
);

AOI32xp33_ASAP7_75t_R c3061(
.A1(net3032),
.A2(net3037),
.A3(net1195),
.B1(net3049),
.B2(net10222),
.Y(net3081)
);

NAND3x2_ASAP7_75t_R c3062(
.B(net3062),
.C(net3003),
.A(net3054),
.Y(net3082)
);

OAI222xp33_ASAP7_75t_R c3063(
.A1(net3080),
.A2(net3070),
.B1(net3068),
.B2(net3073),
.C1(net2891),
.C2(net3034),
.Y(net3083)
);

NAND3xp33_ASAP7_75t_R c3064(
.A(net3080),
.B(net3069),
.C(net10221),
.Y(net3084)
);

NOR3x1_ASAP7_75t_R c3065(
.A(net3056),
.B(net2977),
.C(net3062),
.Y(net3085)
);

ICGx3_ASAP7_75t_R c3066(
.ENA(net3083),
.SE(net3069),
.CLK(clk),
.GCLK(net3086)
);

HB2xp67_ASAP7_75t_R c3067(
.A(net10066),
.Y(net3087)
);

OAI321xp33_ASAP7_75t_R c3068(
.A1(net3046),
.A2(net1827),
.A3(net3085),
.B1(net3087),
.B2(net3080),
.C(net10223),
.Y(net3088)
);

NAND2x1_ASAP7_75t_R c3069(
.A(net3012),
.B(net3087),
.Y(net3089)
);

OAI33xp33_ASAP7_75t_R c3070(
.A1(net3076),
.A2(net3002),
.A3(net3086),
.B1(net3087),
.B2(net3032),
.B3(net10099),
.Y(net3090)
);

HB3xp67_ASAP7_75t_R c3071(
.A(net2218),
.Y(net3091)
);

HB4xp67_ASAP7_75t_R c3072(
.A(net10163),
.Y(net3092)
);

INVx11_ASAP7_75t_R c3073(
.A(net9961),
.Y(net3093)
);

INVx13_ASAP7_75t_R c3074(
.A(net2130),
.Y(net3094)
);

INVx1_ASAP7_75t_R c3075(
.A(net2958),
.Y(net3095)
);

NAND2x1p5_ASAP7_75t_R c3076(
.A(net2193),
.B(net10222),
.Y(net3096)
);

INVx2_ASAP7_75t_R c3077(
.A(net2071),
.Y(net3097)
);

NOR3x2_ASAP7_75t_R c3078(
.B(net353),
.C(net1922),
.A(net2125),
.Y(net3098)
);

NAND2x2_ASAP7_75t_R c3079(
.A(net333),
.B(net10206),
.Y(net3099)
);

INVx3_ASAP7_75t_R c3080(
.A(net10206),
.Y(net3100)
);

NAND2xp33_ASAP7_75t_R c3081(
.A(net2239),
.B(net2143),
.Y(net3101)
);

NAND2xp5_ASAP7_75t_R c3082(
.A(net2231),
.B(net1922),
.Y(net3102)
);

INVx4_ASAP7_75t_R c3083(
.A(net1290),
.Y(net3103)
);

INVx5_ASAP7_75t_R c3084(
.A(net9096),
.Y(net3104)
);

NAND2xp67_ASAP7_75t_R c3085(
.A(net2224),
.B(net3073),
.Y(net3105)
);

NOR2x1_ASAP7_75t_R c3086(
.A(net3010),
.B(net10222),
.Y(net3106)
);

NOR2x1p5_ASAP7_75t_R c3087(
.A(net3099),
.B(net2125),
.Y(net3107)
);

INVx6_ASAP7_75t_R c3088(
.A(net3094),
.Y(net3108)
);

INVx8_ASAP7_75t_R c3089(
.A(net3100),
.Y(net3109)
);

INVxp33_ASAP7_75t_R c3090(
.A(net9096),
.Y(net3110)
);

INVxp67_ASAP7_75t_R c3091(
.A(net3095),
.Y(net3111)
);

NOR3xp33_ASAP7_75t_R c3092(
.A(net3073),
.B(net3104),
.C(net10067),
.Y(net3112)
);

BUFx10_ASAP7_75t_R c3093(
.A(net1963),
.Y(net3113)
);

NOR2x2_ASAP7_75t_R c3094(
.A(net10161),
.B(net10208),
.Y(net3114)
);

BUFx12_ASAP7_75t_R c3095(
.A(net10045),
.Y(net3115)
);

BUFx12f_ASAP7_75t_R c3096(
.A(net3045),
.Y(net3116)
);

NOR2xp33_ASAP7_75t_R c3097(
.A(net2083),
.B(net3093),
.Y(net3117)
);

OA21x2_ASAP7_75t_R c3098(
.A1(net3103),
.A2(net2960),
.B(net1963),
.Y(net3118)
);

BUFx16f_ASAP7_75t_R c3099(
.A(net10545),
.Y(net3119)
);

NOR2xp67_ASAP7_75t_R c3100(
.A(net3011),
.B(net2125),
.Y(net3120)
);

BUFx24_ASAP7_75t_R c3101(
.A(net3115),
.Y(net3121)
);

OAI21x1_ASAP7_75t_R c3102(
.A1(net3102),
.A2(net2210),
.B(net3026),
.Y(net3122)
);

OA31x2_ASAP7_75t_R c3103(
.A1(net3113),
.A2(net3026),
.A3(net10206),
.B1(net10207),
.Y(net3123)
);

BUFx2_ASAP7_75t_R c3104(
.A(net9225),
.Y(net3124)
);

OAI21xp33_ASAP7_75t_R c3105(
.A1(net3097),
.A2(net2083),
.B(net2218),
.Y(net3125)
);

OAI21xp5_ASAP7_75t_R c3106(
.A1(net2779),
.A2(net2163),
.B(net10080),
.Y(net3126)
);

OR3x1_ASAP7_75t_R c3107(
.A(net1212),
.B(net3114),
.C(net3119),
.Y(net3127)
);

OR3x2_ASAP7_75t_R c3108(
.A(net3127),
.B(net2218),
.C(net3115),
.Y(net3128)
);

OR2x2_ASAP7_75t_R c3109(
.A(net2231),
.B(net10012),
.Y(net3129)
);

BUFx3_ASAP7_75t_R c3110(
.A(net3004),
.Y(net3130)
);

BUFx4_ASAP7_75t_R c3111(
.A(net9210),
.Y(net3131)
);

ICGx4DC_ASAP7_75t_R c3112(
.ENA(net3075),
.SE(net3095),
.CLK(clk),
.GCLK(net3132)
);

BUFx4f_ASAP7_75t_R c3113(
.A(net1922),
.Y(net3133)
);

BUFx5_ASAP7_75t_R c3114(
.A(net3110),
.Y(net3134)
);

OR2x4_ASAP7_75t_R c3115(
.A(net3131),
.B(net2164),
.Y(net3135)
);

OR2x6_ASAP7_75t_R c3116(
.A(net3116),
.B(net3119),
.Y(net3136)
);

ICGx4_ASAP7_75t_R c3117(
.ENA(net3125),
.SE(net3069),
.CLK(clk),
.GCLK(net3137)
);

BUFx6f_ASAP7_75t_R c3118(
.A(net3107),
.Y(net3138)
);

XNOR2x1_ASAP7_75t_R c3119(
.B(net3138),
.A(net3133),
.Y(net3139)
);

XNOR2x2_ASAP7_75t_R c3120(
.A(net3114),
.B(net3139),
.Y(net3140)
);

OR3x4_ASAP7_75t_R c3121(
.A(net2226),
.B(net1160),
.C(net3107),
.Y(net3141)
);

OAI211xp5_ASAP7_75t_R c3122(
.A1(net3140),
.A2(net3059),
.B(net3094),
.C(net3134),
.Y(net3142)
);

XNOR2xp5_ASAP7_75t_R c3123(
.A(net3111),
.B(net1238),
.Y(net3143)
);

ICGx5_ASAP7_75t_R c3124(
.ENA(net3117),
.SE(net3142),
.CLK(clk),
.GCLK(net3144)
);

BUFx8_ASAP7_75t_R c3125(
.A(net2176),
.Y(net3145)
);

AND3x1_ASAP7_75t_R c3126(
.A(net3112),
.B(net2219),
.C(net3138),
.Y(net3146)
);

AND3x2_ASAP7_75t_R c3127(
.A(net1277),
.B(net3115),
.C(net3134),
.Y(net3147)
);

CKINVDCx10_ASAP7_75t_R c3128(
.A(net9982),
.Y(net3148)
);

AND3x4_ASAP7_75t_R c3129(
.A(net3143),
.B(net3034),
.C(net3110),
.Y(net3149)
);

SDFLx3_ASAP7_75t_R c3130(
.D(net3126),
.SE(net1190),
.SI(net2224),
.CLK(clk),
.QN(net3150)
);

XOR2x1_ASAP7_75t_R c3131(
.A(net3093),
.B(net3133),
.Y(net3151)
);

XOR2x2_ASAP7_75t_R c3132(
.A(net3106),
.B(net3107),
.Y(net3152)
);

AO21x1_ASAP7_75t_R c3133(
.A1(net3118),
.A2(net3034),
.B(net3144),
.Y(net3153)
);

AO21x2_ASAP7_75t_R c3134(
.A1(net3133),
.A2(net3148),
.B(net3126),
.Y(net3154)
);

XOR2xp5_ASAP7_75t_R c3135(
.A(net3148),
.B(net1212),
.Y(net3155)
);

AND2x2_ASAP7_75t_R c3136(
.A(net3128),
.B(net3124),
.Y(net3156)
);

AND2x4_ASAP7_75t_R c3137(
.A(net2195),
.B(net10012),
.Y(net3157)
);

AOI21x1_ASAP7_75t_R c3138(
.A1(net3155),
.A2(net3151),
.B(net2235),
.Y(net3158)
);

SDFLx4_ASAP7_75t_R c3139(
.D(net3130),
.SE(net2167),
.SI(net3099),
.CLK(clk),
.QN(net3159)
);

AND2x6_ASAP7_75t_R c3140(
.A(net3141),
.B(net3124),
.Y(net3160)
);

HAxp5_ASAP7_75t_R c3141(
.A(net3145),
.B(net10051),
.CON(net3161)
);

NAND2x1_ASAP7_75t_R c3142(
.A(net3147),
.B(net3004),
.Y(net3162)
);

NAND2x1p5_ASAP7_75t_R c3143(
.A(net3134),
.B(net3152),
.Y(net3163)
);

AOI21xp33_ASAP7_75t_R c3144(
.A1(net3161),
.A2(net3159),
.B(net3147),
.Y(net3164)
);

AOI21xp5_ASAP7_75t_R c3145(
.A1(net3164),
.A2(net3137),
.B(net10224),
.Y(net3165)
);

NAND2x2_ASAP7_75t_R c3146(
.A(net3129),
.B(net3059),
.Y(net3166)
);

DFFASRHQNx1_ASAP7_75t_R c3147(
.D(net3166),
.RESETN(net3165),
.SETN(net10223),
.CLK(clk),
.QN(net3167)
);

FAx1_ASAP7_75t_R c3148(
.A(net3165),
.B(net3144),
.CI(net3099),
.SN(net3168)
);

MAJIxp5_ASAP7_75t_R c3149(
.A(net3109),
.B(net3094),
.C(net3163),
.Y(net3169)
);

MAJx2_ASAP7_75t_R c3150(
.A(net3159),
.B(net3167),
.C(net3129),
.Y(net3170)
);

NAND2xp33_ASAP7_75t_R c3151(
.A(net3152),
.B(net3169),
.Y(net3171)
);

AO222x2_ASAP7_75t_R c3152(
.A1(net3171),
.A2(net3153),
.B1(net3170),
.B2(net3134),
.C1(net3144),
.C2(net3163),
.Y(net3172)
);

OAI22x1_ASAP7_75t_R c3153(
.A1(net3169),
.A2(net3159),
.B1(net3155),
.B2(net3163),
.Y(net3173)
);

CKINVDCx11_ASAP7_75t_R c3154(
.A(net10170),
.Y(net3174)
);

CKINVDCx12_ASAP7_75t_R c3155(
.A(net2125),
.Y(net3175)
);

NAND2xp5_ASAP7_75t_R c3156(
.A(net1168),
.B(net2963),
.Y(net3176)
);

CKINVDCx14_ASAP7_75t_R c3157(
.A(net10035),
.Y(net3177)
);

CKINVDCx16_ASAP7_75t_R c3158(
.A(net9961),
.Y(net3178)
);

NAND2xp67_ASAP7_75t_R c3159(
.A(net325),
.B(net3144),
.Y(net3179)
);

CKINVDCx20_ASAP7_75t_R c3160(
.A(net10031),
.Y(net3180)
);

MAJx3_ASAP7_75t_R c3161(
.A(net2291),
.B(net3155),
.C(net3179),
.Y(net3181)
);

CKINVDCx5p33_ASAP7_75t_R c3162(
.A(net10519),
.Y(net3182)
);

CKINVDCx6p67_ASAP7_75t_R c3163(
.A(net3181),
.Y(net3183)
);

NOR2x1_ASAP7_75t_R c3164(
.A(net2271),
.B(net2317),
.Y(net3184)
);

NOR2x1p5_ASAP7_75t_R c3165(
.A(net407),
.B(net2232),
.Y(net3185)
);

CKINVDCx8_ASAP7_75t_R c3166(
.A(net2232),
.Y(net3186)
);

NOR2x2_ASAP7_75t_R c3167(
.A(net2293),
.B(net3177),
.Y(net3187)
);

NOR2xp33_ASAP7_75t_R c3168(
.A(net2321),
.B(net3177),
.Y(net3188)
);

NOR2xp67_ASAP7_75t_R c3169(
.A(net3184),
.B(net10192),
.Y(net3189)
);

CKINVDCx9p33_ASAP7_75t_R c3170(
.A(net3187),
.Y(net3190)
);

HB1xp67_ASAP7_75t_R c3171(
.A(net3178),
.Y(net3191)
);

NAND3x1_ASAP7_75t_R c3172(
.A(net1398),
.B(net3184),
.C(net3010),
.Y(net3192)
);

HB2xp67_ASAP7_75t_R c3173(
.A(net9134),
.Y(net3193)
);

HB3xp67_ASAP7_75t_R c3174(
.A(net3121),
.Y(net3194)
);

HB4xp67_ASAP7_75t_R c3175(
.A(net3191),
.Y(net3195)
);

INVx11_ASAP7_75t_R c3176(
.A(net2319),
.Y(net3196)
);

NAND3x2_ASAP7_75t_R c3177(
.B(net3010),
.C(net2301),
.A(net10210),
.Y(net3197)
);

OR2x2_ASAP7_75t_R c3178(
.A(net3160),
.B(net3146),
.Y(net3198)
);

INVx13_ASAP7_75t_R c3179(
.A(net3179),
.Y(net3199)
);

INVx1_ASAP7_75t_R c3180(
.A(net2313),
.Y(net3200)
);

INVx2_ASAP7_75t_R c3181(
.A(net3190),
.Y(net3201)
);

NAND3xp33_ASAP7_75t_R c3182(
.A(net2312),
.B(net3157),
.C(net2291),
.Y(net3202)
);

INVx3_ASAP7_75t_R c3183(
.A(net9469),
.Y(net3203)
);

INVx4_ASAP7_75t_R c3184(
.A(net10207),
.Y(net3204)
);

OR2x4_ASAP7_75t_R c3185(
.A(net3174),
.B(net3146),
.Y(net3205)
);

AO33x2_ASAP7_75t_R c3186(
.A1(net2230),
.A2(net3175),
.A3(net3167),
.B1(net3204),
.B2(net2235),
.B3(net2268),
.Y(net3206)
);

NOR3x1_ASAP7_75t_R c3187(
.A(net350),
.B(net2261),
.C(net10073),
.Y(net3207)
);

INVx5_ASAP7_75t_R c3188(
.A(net10389),
.Y(net3208)
);

INVx6_ASAP7_75t_R c3189(
.A(net10416),
.Y(net3209)
);

OR2x6_ASAP7_75t_R c3190(
.A(net2204),
.B(net3196),
.Y(net3210)
);

XNOR2x1_ASAP7_75t_R c3191(
.B(net3201),
.A(net3191),
.Y(net3211)
);

XNOR2x2_ASAP7_75t_R c3192(
.A(net3198),
.B(net2313),
.Y(net3212)
);

INVx8_ASAP7_75t_R c3193(
.A(net9210),
.Y(net3213)
);

XNOR2xp5_ASAP7_75t_R c3194(
.A(net3196),
.B(net2313),
.Y(net3214)
);

INVxp33_ASAP7_75t_R c3195(
.A(net10065),
.Y(net3215)
);

XOR2x1_ASAP7_75t_R c3196(
.A(net3205),
.B(net3204),
.Y(net3216)
);

XOR2x2_ASAP7_75t_R c3197(
.A(net3215),
.B(net3197),
.Y(net3217)
);

XOR2xp5_ASAP7_75t_R c3198(
.A(net3217),
.B(net3205),
.Y(net3218)
);

AND2x2_ASAP7_75t_R c3199(
.A(net3213),
.B(net2272),
.Y(net3219)
);

INVxp67_ASAP7_75t_R c3200(
.A(net3204),
.Y(net3220)
);

AND2x4_ASAP7_75t_R c3201(
.A(net3208),
.B(net407),
.Y(net3221)
);

AND2x6_ASAP7_75t_R c3202(
.A(net3197),
.B(net3204),
.Y(net3222)
);

HAxp5_ASAP7_75t_R c3203(
.A(net3210),
.B(net3203),
.CON(net3223)
);

BUFx10_ASAP7_75t_R c3204(
.A(net9907),
.Y(net3224)
);

OAI22xp33_ASAP7_75t_R c3205(
.A1(net3222),
.A2(net3180),
.B1(net2270),
.B2(net3218),
.Y(net3225)
);

BUFx12_ASAP7_75t_R c3206(
.A(net9788),
.Y(net3226)
);

BUFx12f_ASAP7_75t_R c3207(
.A(net3207),
.Y(net3227)
);

NAND2x1_ASAP7_75t_R c3208(
.A(net3209),
.B(net2318),
.Y(net3228)
);

NAND2x1p5_ASAP7_75t_R c3209(
.A(net3216),
.B(net1292),
.Y(net3229)
);

OAI22xp5_ASAP7_75t_R c3210(
.A1(net3026),
.A2(net3222),
.B1(net3057),
.B2(net3134),
.Y(net3230)
);

BUFx16f_ASAP7_75t_R c3211(
.A(net3223),
.Y(net3231)
);

NAND2x2_ASAP7_75t_R c3212(
.A(net1338),
.B(net3210),
.Y(net3232)
);

BUFx24_ASAP7_75t_R c3213(
.A(net3219),
.Y(net3233)
);

NAND5xp2_ASAP7_75t_R c3214(
.A(net3224),
.B(net3229),
.C(net3181),
.D(net3167),
.E(net3190),
.Y(net3234)
);

BUFx2_ASAP7_75t_R c3215(
.A(net10064),
.Y(net3235)
);

AOI222xp33_ASAP7_75t_R c3216(
.A1(net3233),
.A2(net3235),
.B1(net2313),
.B2(net1338),
.C1(net2131),
.C2(net3163),
.Y(net3236)
);

NOR3x2_ASAP7_75t_R c3217(
.B(net2327),
.C(net9763),
.A(net10065),
.Y(net3237)
);

NAND2xp33_ASAP7_75t_R c3218(
.A(net407),
.B(net10073),
.Y(net3238)
);

BUFx3_ASAP7_75t_R c3219(
.A(net3202),
.Y(net3239)
);

BUFx4_ASAP7_75t_R c3220(
.A(net9469),
.Y(net3240)
);

BUFx4f_ASAP7_75t_R c3221(
.A(net3146),
.Y(net3241)
);

NOR3xp33_ASAP7_75t_R c3222(
.A(net3240),
.B(net3198),
.C(net3191),
.Y(net3242)
);

NAND2xp5_ASAP7_75t_R c3223(
.A(net3242),
.B(net9996),
.Y(net3243)
);

NAND2xp67_ASAP7_75t_R c3224(
.A(net3227),
.B(net10165),
.Y(net3244)
);

BUFx5_ASAP7_75t_R c3225(
.A(net9134),
.Y(net3245)
);

NOR2x1_ASAP7_75t_R c3226(
.A(net3168),
.B(net3207),
.Y(net3246)
);

NOR2x1p5_ASAP7_75t_R c3227(
.A(net3242),
.B(net3241),
.Y(net3247)
);

BUFx6f_ASAP7_75t_R c3228(
.A(net3182),
.Y(net3248)
);

NOR2x2_ASAP7_75t_R c3229(
.A(net3241),
.B(net3010),
.Y(net3249)
);

OA21x2_ASAP7_75t_R c3230(
.A1(net3248),
.A2(net2272),
.B(net325),
.Y(net3250)
);

BUFx8_ASAP7_75t_R c3231(
.A(net10035),
.Y(net3251)
);

OAI21x1_ASAP7_75t_R c3232(
.A1(net3250),
.A2(net3134),
.B(net10210),
.Y(net3252)
);

CKINVDCx10_ASAP7_75t_R c3233(
.A(net10039),
.Y(net3253)
);

OAI21xp33_ASAP7_75t_R c3234(
.A1(net3220),
.A2(net3253),
.B(net3226),
.Y(net3254)
);

NOR2xp33_ASAP7_75t_R c3235(
.A(net3251),
.B(net3253),
.Y(net3255)
);

NOR2xp67_ASAP7_75t_R c3236(
.A(net3255),
.B(net10080),
.Y(net3256)
);

CKINVDCx11_ASAP7_75t_R c3237(
.A(net3195),
.Y(net3257)
);

CKINVDCx12_ASAP7_75t_R c3238(
.A(net3006),
.Y(net3258)
);

OR2x2_ASAP7_75t_R c3239(
.A(net3144),
.B(net2317),
.Y(net3259)
);

OR2x4_ASAP7_75t_R c3240(
.A(net2387),
.B(net2365),
.Y(net3260)
);

OR2x6_ASAP7_75t_R c3241(
.A(net1313),
.B(net3258),
.Y(net3261)
);

CKINVDCx14_ASAP7_75t_R c3242(
.A(net1447),
.Y(net3262)
);

CKINVDCx16_ASAP7_75t_R c3243(
.A(net1324),
.Y(net3263)
);

XNOR2x1_ASAP7_75t_R c3244(
.B(net3259),
.A(net1408),
.Y(net3264)
);

CKINVDCx20_ASAP7_75t_R c3245(
.A(net3257),
.Y(net3265)
);

XNOR2x2_ASAP7_75t_R c3246(
.A(net3108),
.B(net2261),
.Y(net3266)
);

CKINVDCx5p33_ASAP7_75t_R c3247(
.A(net10512),
.Y(net3267)
);

OAI21xp5_ASAP7_75t_R c3248(
.A1(net3183),
.A2(net2405),
.B(net3162),
.Y(net3268)
);

XNOR2xp5_ASAP7_75t_R c3249(
.A(net3167),
.B(net3226),
.Y(net3269)
);

XOR2x1_ASAP7_75t_R c3250(
.A(net3265),
.B(net3092),
.Y(net3270)
);

CKINVDCx6p67_ASAP7_75t_R c3251(
.A(net2378),
.Y(net3271)
);

SDFHx1_ASAP7_75t_R c3252(
.D(net3196),
.SE(net3244),
.SI(net3175),
.CLK(clk),
.QN(net3272)
);

XOR2x2_ASAP7_75t_R c3253(
.A(net2272),
.B(net1424),
.Y(net3273)
);

CKINVDCx8_ASAP7_75t_R c3254(
.A(net2159),
.Y(net3274)
);

CKINVDCx9p33_ASAP7_75t_R c3255(
.A(net9955),
.Y(net3275)
);

HB1xp67_ASAP7_75t_R c3256(
.A(net9158),
.Y(net3276)
);

HB2xp67_ASAP7_75t_R c3257(
.A(net10051),
.Y(net3277)
);

XOR2xp5_ASAP7_75t_R c3258(
.A(net3193),
.B(net10212),
.Y(net3278)
);

AND2x2_ASAP7_75t_R c3259(
.A(net3270),
.B(net3269),
.Y(net3279)
);

HB3xp67_ASAP7_75t_R c3260(
.A(net10024),
.Y(net3280)
);

HB4xp67_ASAP7_75t_R c3261(
.A(net9682),
.Y(net3281)
);

AND2x4_ASAP7_75t_R c3262(
.A(net3281),
.B(net3274),
.Y(net3282)
);

INVx11_ASAP7_75t_R c3263(
.A(net3259),
.Y(net3283)
);

AND2x6_ASAP7_75t_R c3264(
.A(net3199),
.B(net10212),
.Y(net3284)
);

INVx13_ASAP7_75t_R c3265(
.A(net3282),
.Y(net3285)
);

HAxp5_ASAP7_75t_R c3266(
.A(net2415),
.B(net1459),
.CON(net3286)
);

NAND2x1_ASAP7_75t_R c3267(
.A(net2210),
.B(net3249),
.Y(net3287)
);

NAND2x1p5_ASAP7_75t_R c3268(
.A(net3144),
.B(net3274),
.Y(net3288)
);

INVx1_ASAP7_75t_R c3269(
.A(net2367),
.Y(net3289)
);

NAND2x2_ASAP7_75t_R c3270(
.A(net3260),
.B(net1348),
.Y(net3290)
);

INVx2_ASAP7_75t_R c3271(
.A(net10560),
.Y(net3291)
);

NAND2xp33_ASAP7_75t_R c3272(
.A(net3285),
.B(net3284),
.Y(net3292)
);

NAND2xp5_ASAP7_75t_R c3273(
.A(net3258),
.B(net2413),
.Y(net3293)
);

NAND2xp67_ASAP7_75t_R c3274(
.A(net327),
.B(net3259),
.Y(net3294)
);

NOR2x1_ASAP7_75t_R c3275(
.A(net3149),
.B(net3269),
.Y(net3295)
);

NOR2x1p5_ASAP7_75t_R c3276(
.A(net3276),
.B(net2390),
.Y(net3296)
);

NOR2x2_ASAP7_75t_R c3277(
.A(net3292),
.B(net10213),
.Y(net3297)
);

INVx3_ASAP7_75t_R c3278(
.A(net10435),
.Y(net3298)
);

OR3x1_ASAP7_75t_R c3279(
.A(net3287),
.B(net2364),
.C(net3214),
.Y(net3299)
);

NOR2xp33_ASAP7_75t_R c3280(
.A(net3262),
.B(net9764),
.Y(net3300)
);

INVx4_ASAP7_75t_R c3281(
.A(net2317),
.Y(net3301)
);

OR3x2_ASAP7_75t_R c3282(
.A(net3288),
.B(net2159),
.C(net3290),
.Y(net3302)
);

NOR2xp67_ASAP7_75t_R c3283(
.A(net3301),
.B(net2415),
.Y(net3303)
);

INVx5_ASAP7_75t_R c3284(
.A(net9158),
.Y(net3304)
);

OR3x4_ASAP7_75t_R c3285(
.A(net3249),
.B(net2378),
.C(net3297),
.Y(net3305)
);

AND3x1_ASAP7_75t_R c3286(
.A(net3295),
.B(net3269),
.C(net512),
.Y(net3306)
);

AND3x2_ASAP7_75t_R c3287(
.A(net3305),
.B(net1408),
.C(net1324),
.Y(net3307)
);

OAI31xp33_ASAP7_75t_R c3288(
.A1(net3306),
.A2(net3273),
.A3(net3239),
.B(net3167),
.Y(net3308)
);

AND3x4_ASAP7_75t_R c3289(
.A(net512),
.B(net3297),
.C(net10225),
.Y(net3309)
);

OR2x2_ASAP7_75t_R c3290(
.A(net1408),
.B(net3258),
.Y(net3310)
);

OR2x4_ASAP7_75t_R c3291(
.A(net2399),
.B(net10112),
.Y(net3311)
);

INVx6_ASAP7_75t_R c3292(
.A(net10563),
.Y(net3312)
);

INVx8_ASAP7_75t_R c3293(
.A(net10505),
.Y(net3313)
);

AO21x1_ASAP7_75t_R c3294(
.A1(net3303),
.A2(net3273),
.B(net3280),
.Y(net3314)
);

OR2x6_ASAP7_75t_R c3295(
.A(net3271),
.B(net1447),
.Y(net3315)
);

INVxp33_ASAP7_75t_R c3296(
.A(net3300),
.Y(net3316)
);

XNOR2x1_ASAP7_75t_R c3297(
.B(net3279),
.A(net1437),
.Y(net3317)
);

XNOR2x2_ASAP7_75t_R c3298(
.A(net2378),
.B(net10054),
.Y(net3318)
);

INVxp67_ASAP7_75t_R c3299(
.A(net10515),
.Y(net3319)
);

XNOR2xp5_ASAP7_75t_R c3300(
.A(net3319),
.B(net3317),
.Y(net3320)
);

OAI31xp67_ASAP7_75t_R c3301(
.A1(net1412),
.A2(net3239),
.A3(net3274),
.B(net3317),
.Y(net3321)
);

XOR2x1_ASAP7_75t_R c3302(
.A(net3304),
.B(net3320),
.Y(net3322)
);

SDFHx2_ASAP7_75t_R c3303(
.D(net3226),
.SE(net3307),
.SI(net3290),
.CLK(clk),
.QN(net3323)
);

XOR2x2_ASAP7_75t_R c3304(
.A(net3292),
.B(net9917),
.Y(net3324)
);

AO21x2_ASAP7_75t_R c3305(
.A1(net3304),
.A2(net3092),
.B(net10225),
.Y(net3325)
);

XOR2xp5_ASAP7_75t_R c3306(
.A(net2261),
.B(net3297),
.Y(net3326)
);

BUFx10_ASAP7_75t_R c3307(
.A(net10080),
.Y(net3327)
);

AOI321xp33_ASAP7_75t_R c3308(
.A1(net3307),
.A2(net3235),
.A3(net3326),
.B1(net3291),
.B2(net3194),
.C(net2045),
.Y(net3328)
);

AOI21x1_ASAP7_75t_R c3309(
.A1(net3293),
.A2(net3305),
.B(net2345),
.Y(net3329)
);

AOI21xp33_ASAP7_75t_R c3310(
.A1(net3320),
.A2(net3270),
.B(net3327),
.Y(net3330)
);

AOI21xp5_ASAP7_75t_R c3311(
.A1(net3324),
.A2(net2261),
.B(net10212),
.Y(net3331)
);

AND2x2_ASAP7_75t_R c3312(
.A(net3283),
.B(net10225),
.Y(net3332)
);

OR4x1_ASAP7_75t_R c3313(
.A(net3313),
.B(net3194),
.C(net3330),
.D(net3327),
.Y(net3333)
);

FAx1_ASAP7_75t_R c3314(
.A(net3323),
.B(net3317),
.CI(net10076),
.SN(net3335),
.CON(net3334)
);

BUFx12_ASAP7_75t_R c3315(
.A(net10421),
.Y(net3336)
);

MAJIxp5_ASAP7_75t_R c3316(
.A(net3336),
.B(net3320),
.C(net10226),
.Y(net3337)
);

AOI33xp33_ASAP7_75t_R c3317(
.A1(net3331),
.A2(net3330),
.A3(net3335),
.B1(net1292),
.B2(net3239),
.B3(net3290),
.Y(net3338)
);

MAJx2_ASAP7_75t_R c3318(
.A(net3291),
.B(net3284),
.C(net9763),
.Y(net3339)
);

MAJx3_ASAP7_75t_R c3319(
.A(net2318),
.B(net2317),
.C(net3336),
.Y(net3340)
);

BUFx12f_ASAP7_75t_R c3320(
.A(net9086),
.Y(net3341)
);

BUFx16f_ASAP7_75t_R c3321(
.A(net2470),
.Y(net3342)
);

AND2x4_ASAP7_75t_R c3322(
.A(net2478),
.B(net2262),
.Y(net3343)
);

BUFx24_ASAP7_75t_R c3323(
.A(net2405),
.Y(net3344)
);

AND2x6_ASAP7_75t_R c3324(
.A(net2219),
.B(net3335),
.Y(net3345)
);

HAxp5_ASAP7_75t_R c3325(
.A(net2396),
.B(net3194),
.CON(net3347),
.SN(net3346)
);

BUFx2_ASAP7_75t_R c3326(
.A(net2472),
.Y(net3348)
);

BUFx3_ASAP7_75t_R c3327(
.A(net10100),
.Y(net3349)
);

BUFx4_ASAP7_75t_R c3328(
.A(net598),
.Y(net3350)
);

BUFx4f_ASAP7_75t_R c3329(
.A(net10414),
.Y(net3351)
);

NAND2x1_ASAP7_75t_R c3330(
.A(net2332),
.B(net2259),
.Y(net3352)
);

BUFx5_ASAP7_75t_R c3331(
.A(net10393),
.Y(net3353)
);

BUFx6f_ASAP7_75t_R c3332(
.A(net2439),
.Y(net3354)
);

BUFx8_ASAP7_75t_R c3333(
.A(net3352),
.Y(net3355)
);

ICGx5p33DC_ASAP7_75t_R c3334(
.ENA(net2471),
.SE(net3194),
.CLK(clk),
.GCLK(net3356)
);

NAND2x1p5_ASAP7_75t_R c3335(
.A(net3289),
.B(net2470),
.Y(net3357)
);

CKINVDCx10_ASAP7_75t_R c3336(
.A(net3342),
.Y(net3358)
);

CKINVDCx11_ASAP7_75t_R c3337(
.A(net3358),
.Y(net3359)
);

NAND2x2_ASAP7_75t_R c3338(
.A(net3357),
.B(net3291),
.Y(net3360)
);

NAND2xp33_ASAP7_75t_R c3339(
.A(net2045),
.B(net1534),
.Y(net3361)
);

CKINVDCx12_ASAP7_75t_R c3340(
.A(net9252),
.Y(net3362)
);

NAND3x1_ASAP7_75t_R c3341(
.A(net3341),
.B(net3350),
.C(net3346),
.Y(net3363)
);

CKINVDCx14_ASAP7_75t_R c3342(
.A(net3326),
.Y(net3364)
);

NAND2xp5_ASAP7_75t_R c3343(
.A(net3284),
.B(net3327),
.Y(net3365)
);

SDFHx3_ASAP7_75t_R c3344(
.D(net2479),
.SE(net2332),
.SI(net3162),
.CLK(clk),
.QN(net3366)
);

NAND2xp67_ASAP7_75t_R c3345(
.A(net3356),
.B(net3362),
.Y(net3367)
);

CKINVDCx16_ASAP7_75t_R c3346(
.A(net9252),
.Y(net3368)
);

NOR2x1_ASAP7_75t_R c3347(
.A(net3350),
.B(net3292),
.Y(net3369)
);

NAND3x2_ASAP7_75t_R c3348(
.B(net2483),
.C(net3350),
.A(net2404),
.Y(net3370)
);

NOR2x1p5_ASAP7_75t_R c3349(
.A(net3270),
.B(net3356),
.Y(net3371)
);

CKINVDCx20_ASAP7_75t_R c3350(
.A(net3365),
.Y(net3372)
);

CKINVDCx5p33_ASAP7_75t_R c3351(
.A(net10373),
.Y(net3373)
);

NOR2x2_ASAP7_75t_R c3352(
.A(net2460),
.B(net2478),
.Y(net3374)
);

NOR2xp33_ASAP7_75t_R c3353(
.A(net1534),
.B(net3372),
.Y(net3375)
);

CKINVDCx6p67_ASAP7_75t_R c3354(
.A(net10432),
.Y(net3376)
);

CKINVDCx8_ASAP7_75t_R c3355(
.A(net2456),
.Y(net3377)
);

CKINVDCx9p33_ASAP7_75t_R c3356(
.A(net3374),
.Y(net3378)
);

HB1xp67_ASAP7_75t_R c3357(
.A(net10490),
.Y(net3379)
);

NOR2xp67_ASAP7_75t_R c3358(
.A(net3377),
.B(net3292),
.Y(net3380)
);

OR2x2_ASAP7_75t_R c3359(
.A(net3368),
.B(net3379),
.Y(net3381)
);

HB2xp67_ASAP7_75t_R c3360(
.A(net3323),
.Y(net3382)
);

OR2x4_ASAP7_75t_R c3361(
.A(net1340),
.B(net3355),
.Y(net3383)
);

OR2x6_ASAP7_75t_R c3362(
.A(net2466),
.B(net3379),
.Y(net3384)
);

XNOR2x1_ASAP7_75t_R c3363(
.B(net3372),
.A(net3256),
.Y(net3385)
);

XNOR2x2_ASAP7_75t_R c3364(
.A(net3370),
.B(net3382),
.Y(net3386)
);

XNOR2xp5_ASAP7_75t_R c3365(
.A(net3344),
.B(net3375),
.Y(net3387)
);

XOR2x1_ASAP7_75t_R c3366(
.A(net3378),
.B(net3347),
.Y(net3388)
);

HB3xp67_ASAP7_75t_R c3367(
.A(net3379),
.Y(net3389)
);

XOR2x2_ASAP7_75t_R c3368(
.A(net3353),
.B(net2427),
.Y(net3390)
);

OA222x2_ASAP7_75t_R c3369(
.A1(net3252),
.A2(net3382),
.B1(net2498),
.B2(net3273),
.C1(net2427),
.C2(net1446),
.Y(net3391)
);

HB4xp67_ASAP7_75t_R c3370(
.A(net10152),
.Y(net3392)
);

NAND3xp33_ASAP7_75t_R c3371(
.A(net3356),
.B(net3379),
.C(net10198),
.Y(net3393)
);

INVx11_ASAP7_75t_R c3372(
.A(net10148),
.Y(net3394)
);

XOR2xp5_ASAP7_75t_R c3373(
.A(net3388),
.B(net3379),
.Y(net3395)
);

INVx13_ASAP7_75t_R c3374(
.A(net10440),
.Y(net3396)
);

INVx1_ASAP7_75t_R c3375(
.A(net3371),
.Y(net3397)
);

INVx2_ASAP7_75t_R c3376(
.A(net3380),
.Y(net3398)
);

NOR5xp2_ASAP7_75t_R c3377(
.A(net1437),
.B(net3382),
.C(net3392),
.D(net2459),
.E(net2498),
.Y(net3399)
);

NOR3x1_ASAP7_75t_R c3378(
.A(net3347),
.B(net3398),
.C(net2779),
.Y(net3400)
);

NOR3x2_ASAP7_75t_R c3379(
.B(net2335),
.C(net3272),
.A(net3398),
.Y(net3401)
);

AND2x2_ASAP7_75t_R c3380(
.A(net3396),
.B(net3379),
.Y(net3402)
);

AND2x4_ASAP7_75t_R c3381(
.A(net3376),
.B(net3382),
.Y(net3403)
);

NOR3xp33_ASAP7_75t_R c3382(
.A(net3292),
.B(net3386),
.C(net3382),
.Y(net3404)
);

INVx3_ASAP7_75t_R c3383(
.A(net10076),
.Y(net3405)
);

AND2x6_ASAP7_75t_R c3384(
.A(net3263),
.B(net2470),
.Y(net3406)
);

HAxp5_ASAP7_75t_R c3385(
.A(net3399),
.B(net3398),
.CON(net3407)
);

NAND2x1_ASAP7_75t_R c3386(
.A(net3382),
.B(net3396),
.Y(net3408)
);

OA21x2_ASAP7_75t_R c3387(
.A1(net3392),
.A2(net3363),
.B(net2404),
.Y(net3409)
);

NAND2x1p5_ASAP7_75t_R c3388(
.A(net3405),
.B(net3342),
.Y(net3410)
);

OAI21x1_ASAP7_75t_R c3389(
.A1(net3394),
.A2(net3364),
.B(net3372),
.Y(net3411)
);

INVx4_ASAP7_75t_R c3390(
.A(net9086),
.Y(net3412)
);

NAND2x2_ASAP7_75t_R c3391(
.A(net3402),
.B(net3412),
.Y(net3413)
);

NAND2xp33_ASAP7_75t_R c3392(
.A(net3375),
.B(net3402),
.Y(net3414)
);

OAI21xp33_ASAP7_75t_R c3393(
.A1(net3384),
.A2(net3413),
.B(net3414),
.Y(net3415)
);

NAND2xp5_ASAP7_75t_R c3394(
.A(net3407),
.B(net3414),
.Y(net3416)
);

OAI21xp5_ASAP7_75t_R c3395(
.A1(net3397),
.A2(net3398),
.B(net3412),
.Y(net3417)
);

SDFHx4_ASAP7_75t_R c3396(
.D(net3398),
.SE(net3395),
.SI(net3417),
.CLK(clk),
.QN(net3418)
);

NAND2xp67_ASAP7_75t_R c3397(
.A(net3409),
.B(net9634),
.Y(net3419)
);

OR3x1_ASAP7_75t_R c3398(
.A(net2501),
.B(net1250),
.C(net3418),
.Y(net3420)
);

OR3x2_ASAP7_75t_R c3399(
.A(net3420),
.B(net3413),
.C(net3398),
.Y(net3421)
);

OR3x4_ASAP7_75t_R c3400(
.A(net2402),
.B(net3408),
.C(net3421),
.Y(net3422)
);

NOR2x1_ASAP7_75t_R c3401(
.A(net3418),
.B(net9634),
.Y(net3423)
);

AND3x1_ASAP7_75t_R c3402(
.A(net3423),
.B(net3412),
.C(net9855),
.Y(net3424)
);

NOR2x1p5_ASAP7_75t_R c3403(
.A(net2517),
.B(net662),
.Y(net3425)
);

NOR2x2_ASAP7_75t_R c3404(
.A(net3349),
.B(net3393),
.Y(net3426)
);

NOR2xp33_ASAP7_75t_R c3405(
.A(net1292),
.B(net10214),
.Y(net3427)
);

NOR2xp67_ASAP7_75t_R c3406(
.A(net1536),
.B(net2459),
.Y(net3428)
);

OR2x2_ASAP7_75t_R c3407(
.A(net483),
.B(net3386),
.Y(net3429)
);

INVx5_ASAP7_75t_R c3408(
.A(net9994),
.Y(net3430)
);

INVx6_ASAP7_75t_R c3409(
.A(net9898),
.Y(net3431)
);

INVx8_ASAP7_75t_R c3410(
.A(net3354),
.Y(net3432)
);

INVxp33_ASAP7_75t_R c3411(
.A(net3311),
.Y(net3433)
);

ICGx6p67DC_ASAP7_75t_R c3412(
.ENA(net3317),
.SE(net2474),
.CLK(clk),
.GCLK(net3434)
);

INVxp67_ASAP7_75t_R c3413(
.A(net9994),
.Y(net3435)
);

BUFx10_ASAP7_75t_R c3414(
.A(net3415),
.Y(net3436)
);

OR2x4_ASAP7_75t_R c3415(
.A(net3359),
.B(net2517),
.Y(net3437)
);

OR2x6_ASAP7_75t_R c3416(
.A(net3417),
.B(net3363),
.Y(net3438)
);

BUFx12_ASAP7_75t_R c3417(
.A(net3262),
.Y(net3439)
);

AND3x2_ASAP7_75t_R c3418(
.A(net3175),
.B(net3383),
.C(net2517),
.Y(net3440)
);

BUFx12f_ASAP7_75t_R c3419(
.A(net10495),
.Y(net3441)
);

XNOR2x1_ASAP7_75t_R c3420(
.B(net3369),
.A(net3410),
.Y(net3442)
);

BUFx16f_ASAP7_75t_R c3421(
.A(net10107),
.Y(net3443)
);

BUFx24_ASAP7_75t_R c3422(
.A(net3355),
.Y(net3444)
);

XNOR2x2_ASAP7_75t_R c3423(
.A(net3434),
.B(net3355),
.Y(net3445)
);

SDFLx1_ASAP7_75t_R c3424(
.D(net1457),
.SE(net3317),
.SI(net624),
.CLK(clk),
.QN(net3446)
);

XNOR2xp5_ASAP7_75t_R c3425(
.A(net3312),
.B(net3446),
.Y(net3447)
);

XOR2x1_ASAP7_75t_R c3426(
.A(net2358),
.B(net2578),
.Y(net3448)
);

XOR2x2_ASAP7_75t_R c3427(
.A(net722),
.B(net2459),
.Y(net3449)
);

XOR2xp5_ASAP7_75t_R c3428(
.A(net3410),
.B(net3417),
.Y(net3450)
);

AND2x2_ASAP7_75t_R c3429(
.A(net1570),
.B(net3317),
.Y(net3451)
);

AND2x4_ASAP7_75t_R c3430(
.A(net3442),
.B(net10214),
.Y(net3452)
);

BUFx2_ASAP7_75t_R c3431(
.A(net9994),
.Y(net3453)
);

AND3x4_ASAP7_75t_R c3432(
.A(net3440),
.B(net3449),
.C(net1651),
.Y(net3454)
);

AND2x6_ASAP7_75t_R c3433(
.A(net3351),
.B(net2427),
.Y(net3455)
);

HAxp5_ASAP7_75t_R c3434(
.A(net3446),
.B(net10208),
.CON(net3456)
);

BUFx3_ASAP7_75t_R c3435(
.A(net10078),
.Y(net3457)
);

BUFx4_ASAP7_75t_R c3436(
.A(net10003),
.Y(net3458)
);

NAND2x1_ASAP7_75t_R c3437(
.A(net3451),
.B(net10214),
.Y(net3459)
);

BUFx4f_ASAP7_75t_R c3438(
.A(net3439),
.Y(net3460)
);

NAND2x1p5_ASAP7_75t_R c3439(
.A(net1454),
.B(net3443),
.Y(net3461)
);

BUFx5_ASAP7_75t_R c3440(
.A(net10520),
.Y(net3462)
);

NAND2x2_ASAP7_75t_R c3441(
.A(net3431),
.B(net2517),
.Y(net3463)
);

BUFx6f_ASAP7_75t_R c3442(
.A(net9926),
.Y(net3464)
);

NAND2xp33_ASAP7_75t_R c3443(
.A(net3444),
.B(net2529),
.Y(net3465)
);

NAND2xp5_ASAP7_75t_R c3444(
.A(net3447),
.B(net3452),
.Y(net3466)
);

BUFx8_ASAP7_75t_R c3445(
.A(net10367),
.Y(net3467)
);

NAND2xp67_ASAP7_75t_R c3446(
.A(net2544),
.B(net3448),
.Y(net3468)
);

CKINVDCx10_ASAP7_75t_R c3447(
.A(net10056),
.Y(net3469)
);

AO21x1_ASAP7_75t_R c3448(
.A1(net3462),
.A2(net2045),
.B(net3453),
.Y(net3470)
);

NOR2x1_ASAP7_75t_R c3449(
.A(net3441),
.B(net3459),
.Y(net3471)
);

NOR2x1p5_ASAP7_75t_R c3450(
.A(net3430),
.B(net3363),
.Y(net3472)
);

NOR2x2_ASAP7_75t_R c3451(
.A(net3460),
.B(net10015),
.Y(net3473)
);

CKINVDCx11_ASAP7_75t_R c3452(
.A(net10160),
.Y(net3474)
);

NOR2xp33_ASAP7_75t_R c3453(
.A(net3465),
.B(net10015),
.Y(net3475)
);

NOR2xp67_ASAP7_75t_R c3454(
.A(net3393),
.B(net3427),
.Y(net3476)
);

OR2x2_ASAP7_75t_R c3455(
.A(net3453),
.B(net3473),
.Y(net3477)
);

OR2x4_ASAP7_75t_R c3456(
.A(net3386),
.B(net2502),
.Y(net3478)
);

OR2x6_ASAP7_75t_R c3457(
.A(net2250),
.B(net3429),
.Y(net3479)
);

XNOR2x1_ASAP7_75t_R c3458(
.B(net3446),
.A(net9986),
.Y(net3480)
);

AO21x2_ASAP7_75t_R c3459(
.A1(net3367),
.A2(net3480),
.B(net3453),
.Y(net3481)
);

XNOR2x2_ASAP7_75t_R c3460(
.A(net3470),
.B(net3355),
.Y(net3482)
);

XNOR2xp5_ASAP7_75t_R c3461(
.A(net3473),
.B(net3445),
.Y(net3483)
);

XOR2x1_ASAP7_75t_R c3462(
.A(net3474),
.B(net3445),
.Y(net3484)
);

XOR2x2_ASAP7_75t_R c3463(
.A(net3426),
.B(net3484),
.Y(net3485)
);

XOR2xp5_ASAP7_75t_R c3464(
.A(net3391),
.B(net3485),
.Y(net3486)
);

AOI21x1_ASAP7_75t_R c3465(
.A1(net3472),
.A2(net2569),
.B(net3481),
.Y(net3487)
);

OA33x2_ASAP7_75t_R c3466(
.A1(net3456),
.A2(net3343),
.A3(net3429),
.B1(net3481),
.B2(net2517),
.B3(net3432),
.Y(net3488)
);

OA221x2_ASAP7_75t_R c3467(
.A1(net3487),
.A2(net1625),
.B1(net3449),
.B2(net3447),
.C(net3481),
.Y(net3489)
);

AND2x2_ASAP7_75t_R c3468(
.A(net3458),
.B(net1612),
.Y(net3490)
);

CKINVDCx12_ASAP7_75t_R c3469(
.A(net10003),
.Y(net3491)
);

CKINVDCx14_ASAP7_75t_R c3470(
.A(net9957),
.Y(net3492)
);

AOI21xp33_ASAP7_75t_R c3471(
.A1(net3193),
.A2(net3483),
.B(net3434),
.Y(net3493)
);

CKINVDCx16_ASAP7_75t_R c3472(
.A(net10388),
.Y(net3494)
);

AND2x4_ASAP7_75t_R c3473(
.A(net3494),
.B(net659),
.Y(net3495)
);

AND2x6_ASAP7_75t_R c3474(
.A(net3495),
.B(net10002),
.Y(net3496)
);

HAxp5_ASAP7_75t_R c3475(
.A(net3414),
.B(net3432),
.CON(net3498),
.SN(net3497)
);

NAND2x1_ASAP7_75t_R c3476(
.A(net3473),
.B(net10002),
.Y(net3499)
);

NAND2x1p5_ASAP7_75t_R c3477(
.A(net2525),
.B(net3499),
.Y(net3500)
);

AOI21xp5_ASAP7_75t_R c3478(
.A1(net3500),
.A2(net3447),
.B(net3485),
.Y(net3501)
);

FAx1_ASAP7_75t_R c3479(
.A(net3500),
.B(net3434),
.CI(net9986),
.SN(net3502)
);

OAI221xp5_ASAP7_75t_R c3480(
.A1(net3499),
.A2(net3415),
.B1(net3481),
.B2(net3432),
.C(net1526),
.Y(net3503)
);

NAND2x2_ASAP7_75t_R c3481(
.A(net3498),
.B(net3427),
.Y(net3504)
);

NAND2xp33_ASAP7_75t_R c3482(
.A(net3493),
.B(net3497),
.Y(net3505)
);

NAND2xp5_ASAP7_75t_R c3483(
.A(net2386),
.B(net3493),
.Y(net3506)
);

OAI311xp33_ASAP7_75t_R c3484(
.A1(net3505),
.A2(net3493),
.A3(net3500),
.B1(net3272),
.C1(net3481),
.Y(net3507)
);

OR4x2_ASAP7_75t_R c3485(
.A(net2531),
.B(net3500),
.C(net3481),
.D(net10228),
.Y(net3508)
);

CKINVDCx20_ASAP7_75t_R c3486(
.A(net805),
.Y(net3509)
);

CKINVDCx5p33_ASAP7_75t_R c3487(
.A(net10022),
.Y(net3510)
);

NAND2xp67_ASAP7_75t_R c3488(
.A(net2633),
.B(net2615),
.Y(net3511)
);

CKINVDCx6p67_ASAP7_75t_R c3489(
.A(net10227),
.Y(net3512)
);

NOR2x1_ASAP7_75t_R c3490(
.A(net2610),
.B(net2668),
.Y(net3513)
);

NOR2x1p5_ASAP7_75t_R c3491(
.A(net2645),
.B(net10179),
.Y(net3514)
);

CKINVDCx8_ASAP7_75t_R c3492(
.A(net9087),
.Y(net3515)
);

NOR2x2_ASAP7_75t_R c3493(
.A(net3448),
.B(net2667),
.Y(net3516)
);

NOR2xp33_ASAP7_75t_R c3494(
.A(net1700),
.B(net738),
.Y(net3517)
);

CKINVDCx9p33_ASAP7_75t_R c3495(
.A(net10087),
.Y(net3518)
);

MAJIxp5_ASAP7_75t_R c3496(
.A(net1600),
.B(net3490),
.C(net3481),
.Y(net3519)
);

NOR2xp67_ASAP7_75t_R c3497(
.A(net2597),
.B(net3519),
.Y(net3520)
);

HB1xp67_ASAP7_75t_R c3498(
.A(net9657),
.Y(net3521)
);

OR2x2_ASAP7_75t_R c3499(
.A(net2616),
.B(net3361),
.Y(net3522)
);

HB2xp67_ASAP7_75t_R c3500(
.A(net1616),
.Y(net3523)
);

A2O1A1Ixp33_ASAP7_75t_R c3501(
.A1(net754),
.A2(net2581),
.B(net3519),
.C(net9941),
.Y(net3524)
);

HB3xp67_ASAP7_75t_R c3502(
.A(net2658),
.Y(net3525)
);

MAJx2_ASAP7_75t_R c3503(
.A(net2663),
.B(net3523),
.C(net2620),
.Y(net3526)
);

HB4xp67_ASAP7_75t_R c3504(
.A(net9087),
.Y(net3527)
);

MAJx3_ASAP7_75t_R c3505(
.A(net446),
.B(net3360),
.C(net2620),
.Y(net3528)
);

SDFLx2_ASAP7_75t_R c3506(
.D(net3457),
.SE(net2663),
.SI(net3523),
.CLK(clk),
.QN(net3529)
);

OR2x4_ASAP7_75t_R c3507(
.A(net3518),
.B(net3445),
.Y(net3530)
);

AND4x1_ASAP7_75t_R c3508(
.A(net3509),
.B(net2590),
.C(net3529),
.D(net3481),
.Y(net3531)
);

NAND3x1_ASAP7_75t_R c3509(
.A(net2619),
.B(net3510),
.C(net9647),
.Y(net3532)
);

OR2x6_ASAP7_75t_R c3510(
.A(net3194),
.B(net1664),
.Y(net3533)
);

XNOR2x1_ASAP7_75t_R c3511(
.B(net3446),
.A(net803),
.Y(net3534)
);

INVx11_ASAP7_75t_R c3512(
.A(net10109),
.Y(net3535)
);

NAND3x2_ASAP7_75t_R c3513(
.B(net1700),
.C(net3527),
.A(net10054),
.Y(net3536)
);

INVx13_ASAP7_75t_R c3514(
.A(net10568),
.Y(net3537)
);

XNOR2x2_ASAP7_75t_R c3515(
.A(net2667),
.B(net2630),
.Y(net3538)
);

INVx1_ASAP7_75t_R c3516(
.A(net10545),
.Y(net3539)
);

XNOR2xp5_ASAP7_75t_R c3517(
.A(net2574),
.B(net3523),
.Y(net3540)
);

XOR2x1_ASAP7_75t_R c3518(
.A(net3521),
.B(net803),
.Y(net3541)
);

XOR2x2_ASAP7_75t_R c3519(
.A(net1611),
.B(net3539),
.Y(net3542)
);

XOR2xp5_ASAP7_75t_R c3520(
.A(net3527),
.B(net3539),
.Y(net3543)
);

AND2x2_ASAP7_75t_R c3521(
.A(net3534),
.B(net1709),
.Y(net3544)
);

INVx2_ASAP7_75t_R c3522(
.A(net3536),
.Y(net3545)
);

AND2x4_ASAP7_75t_R c3523(
.A(net3545),
.B(net3537),
.Y(net3546)
);

AND2x6_ASAP7_75t_R c3524(
.A(net3383),
.B(net3519),
.Y(net3547)
);

HAxp5_ASAP7_75t_R c3525(
.A(net2552),
.B(net3545),
.CON(net3549),
.SN(net3548)
);

NAND3xp33_ASAP7_75t_R c3526(
.A(net1694),
.B(net2633),
.C(net10062),
.Y(net3550)
);

NAND2x1_ASAP7_75t_R c3527(
.A(net2630),
.B(net2581),
.Y(net3551)
);

NAND2x1p5_ASAP7_75t_R c3528(
.A(net2613),
.B(net3541),
.Y(net3552)
);

NOR3x1_ASAP7_75t_R c3529(
.A(net3546),
.B(net3535),
.C(net3532),
.Y(net3553)
);

INVx3_ASAP7_75t_R c3530(
.A(net9952),
.Y(net3554)
);

NAND2x2_ASAP7_75t_R c3531(
.A(net3511),
.B(net2581),
.Y(net3555)
);

NOR3x2_ASAP7_75t_R c3532(
.B(net2598),
.C(net3546),
.A(net3523),
.Y(net3556)
);

NAND2xp33_ASAP7_75t_R c3533(
.A(net3553),
.B(net3512),
.Y(net3557)
);

NAND2xp5_ASAP7_75t_R c3534(
.A(net3539),
.B(net10227),
.Y(net3558)
);

NAND2xp67_ASAP7_75t_R c3535(
.A(net799),
.B(net2661),
.Y(net3559)
);

NOR2x1_ASAP7_75t_R c3536(
.A(net3544),
.B(net3432),
.Y(net3560)
);

INVx4_ASAP7_75t_R c3537(
.A(net10102),
.Y(net3561)
);

NOR2x1p5_ASAP7_75t_R c3538(
.A(net3520),
.B(net3546),
.Y(net3562)
);

INVx5_ASAP7_75t_R c3539(
.A(net10556),
.Y(net3563)
);

ICGx8DC_ASAP7_75t_R c3540(
.ENA(net3524),
.SE(net3546),
.CLK(clk),
.GCLK(net3564)
);

NOR2x2_ASAP7_75t_R c3541(
.A(net3559),
.B(net2337),
.Y(net3565)
);

NOR2xp33_ASAP7_75t_R c3542(
.A(net3530),
.B(net3541),
.Y(net3566)
);

NOR2xp67_ASAP7_75t_R c3543(
.A(net3540),
.B(net1600),
.Y(net3567)
);

NOR3xp33_ASAP7_75t_R c3544(
.A(net3549),
.B(net3550),
.C(net2474),
.Y(net3568)
);

OAI222xp33_ASAP7_75t_R c3545(
.A1(net3558),
.A2(net3548),
.B1(net659),
.B2(net2574),
.C1(net3547),
.C2(net3537),
.Y(net3569)
);

OR2x2_ASAP7_75t_R c3546(
.A(net3567),
.B(net3565),
.Y(net3570)
);

ICGx1_ASAP7_75t_R c3547(
.ENA(net3533),
.SE(net2474),
.CLK(clk),
.GCLK(net3571)
);

OR2x4_ASAP7_75t_R c3548(
.A(net3528),
.B(net3527),
.Y(net3572)
);

OA21x2_ASAP7_75t_R c3549(
.A1(net3563),
.A2(net3571),
.B(net3550),
.Y(net3573)
);

OR2x6_ASAP7_75t_R c3550(
.A(net3570),
.B(net2337),
.Y(net3574)
);

OAI321xp33_ASAP7_75t_R c3551(
.A1(net3531),
.A2(net3570),
.A3(net3546),
.B1(net3557),
.B2(net3564),
.C(net10227),
.Y(net3575)
);

XNOR2x1_ASAP7_75t_R c3552(
.B(net3547),
.A(net3531),
.Y(net3576)
);

OAI21x1_ASAP7_75t_R c3553(
.A1(net711),
.A2(net3560),
.B(net10213),
.Y(net3577)
);

INVx6_ASAP7_75t_R c3554(
.A(net3523),
.Y(net3578)
);

OAI32xp33_ASAP7_75t_R c3555(
.A1(net2585),
.A2(net3572),
.A3(net3553),
.B1(net3537),
.B2(net1664),
.Y(net3579)
);

SDFLx3_ASAP7_75t_R c3556(
.D(net3576),
.SE(net3524),
.SI(net3315),
.CLK(clk),
.QN(net3580)
);

XNOR2x2_ASAP7_75t_R c3557(
.A(net3445),
.B(net3539),
.Y(net3581)
);

OAI21xp33_ASAP7_75t_R c3558(
.A1(net3571),
.A2(net3536),
.B(net9842),
.Y(net3582)
);

AND4x2_ASAP7_75t_R c3559(
.A(net3574),
.B(net3547),
.C(net3538),
.D(net3580),
.Y(net3583)
);

OR5x1_ASAP7_75t_R c3560(
.A(net2636),
.B(net3564),
.C(net2620),
.D(net3537),
.E(net10105),
.Y(net3584)
);

OAI21xp5_ASAP7_75t_R c3561(
.A1(net3581),
.A2(net1653),
.B(net2581),
.Y(net3585)
);

INVx8_ASAP7_75t_R c3562(
.A(net10511),
.Y(net3586)
);

OR5x2_ASAP7_75t_R c3563(
.A(net3515),
.B(net3545),
.C(net3586),
.D(net3537),
.E(net1611),
.Y(net3587)
);

OR3x1_ASAP7_75t_R c3564(
.A(net1568),
.B(net3580),
.C(net1726),
.Y(net3588)
);

OR3x2_ASAP7_75t_R c3565(
.A(net3584),
.B(net3586),
.C(net10097),
.Y(net3589)
);

AO211x2_ASAP7_75t_R c3566(
.A1(net3550),
.A2(net2380),
.B(net2589),
.C(net3529),
.Y(net3590)
);

AO22x1_ASAP7_75t_R c3567(
.A1(net3589),
.A2(net3519),
.B1(net10097),
.B2(net10229),
.Y(net3591)
);

A2O1A1O1Ixp25_ASAP7_75t_R c3568(
.A1(net3538),
.A2(net2661),
.B(net3586),
.C(net9986),
.D(net10229),
.Y(net3592)
);

AO22x2_ASAP7_75t_R c3569(
.A1(net3361),
.A2(net1807),
.B1(net3481),
.B2(net1774),
.Y(net3593)
);

XNOR2xp5_ASAP7_75t_R c3570(
.A(net866),
.B(net3484),
.Y(net3594)
);

XOR2x1_ASAP7_75t_R c3571(
.A(net1807),
.B(net738),
.Y(net3595)
);

XOR2x2_ASAP7_75t_R c3572(
.A(net1791),
.B(net2744),
.Y(net3596)
);

XOR2xp5_ASAP7_75t_R c3573(
.A(net2711),
.B(net2708),
.Y(net3597)
);

INVxp33_ASAP7_75t_R c3574(
.A(net10330),
.Y(net3598)
);

AND2x2_ASAP7_75t_R c3575(
.A(net2744),
.B(net1720),
.Y(net3599)
);

INVxp67_ASAP7_75t_R c3576(
.A(net10349),
.Y(net3600)
);

OR3x4_ASAP7_75t_R c3577(
.A(net836),
.B(net2638),
.C(net1787),
.Y(net3601)
);

ICGx2_ASAP7_75t_R c3578(
.ENA(net2671),
.SE(net3519),
.CLK(clk),
.GCLK(net3602)
);

AND2x4_ASAP7_75t_R c3579(
.A(net1744),
.B(net2712),
.Y(net3603)
);

AND2x6_ASAP7_75t_R c3580(
.A(net2673),
.B(net3529),
.Y(net3604)
);

HAxp5_ASAP7_75t_R c3581(
.A(net876),
.B(net10160),
.CON(net3605)
);

AND3x1_ASAP7_75t_R c3582(
.A(net3529),
.B(net3604),
.C(net3602),
.Y(net3606)
);

NAND2x1_ASAP7_75t_R c3583(
.A(net2669),
.B(net9984),
.Y(net3607)
);

NAND2x1p5_ASAP7_75t_R c3584(
.A(net3607),
.B(net10228),
.Y(net3608)
);

NAND2x2_ASAP7_75t_R c3585(
.A(net2729),
.B(net2619),
.Y(net3609)
);

NAND2xp33_ASAP7_75t_R c3586(
.A(net1748),
.B(net1720),
.Y(net3610)
);

SDFLx4_ASAP7_75t_R c3587(
.D(net873),
.SE(net2615),
.SI(net2708),
.CLK(clk),
.QN(net3611)
);

NAND2xp5_ASAP7_75t_R c3588(
.A(net3595),
.B(net1787),
.Y(net3612)
);

AND3x2_ASAP7_75t_R c3589(
.A(net2700),
.B(net1720),
.C(net2719),
.Y(net3613)
);

NAND2xp67_ASAP7_75t_R c3590(
.A(net1561),
.B(net9858),
.Y(net3614)
);

BUFx10_ASAP7_75t_R c3591(
.A(net10495),
.Y(net3615)
);

ICGx2p67DC_ASAP7_75t_R c3592(
.ENA(net2748),
.SE(net3608),
.CLK(clk),
.GCLK(net3616)
);

NOR2x1_ASAP7_75t_R c3593(
.A(net2734),
.B(net3513),
.Y(net3617)
);

AND3x4_ASAP7_75t_R c3594(
.A(net3593),
.B(net1807),
.C(net10216),
.Y(net3618)
);

NOR2x1p5_ASAP7_75t_R c3595(
.A(net3514),
.B(net2584),
.Y(net3619)
);

NOR2x2_ASAP7_75t_R c3596(
.A(net1802),
.B(net3609),
.Y(net3620)
);

NOR2xp33_ASAP7_75t_R c3597(
.A(net3598),
.B(net9805),
.Y(net3621)
);

NOR2xp67_ASAP7_75t_R c3598(
.A(net2696),
.B(net1769),
.Y(net3622)
);

AO21x1_ASAP7_75t_R c3599(
.A1(net3620),
.A2(net3593),
.B(net836),
.Y(net3623)
);

AO21x2_ASAP7_75t_R c3600(
.A1(net3621),
.A2(net3620),
.B(net2707),
.Y(net3624)
);

OR2x2_ASAP7_75t_R c3601(
.A(net2693),
.B(net2719),
.Y(net3625)
);

OR2x4_ASAP7_75t_R c3602(
.A(net2645),
.B(net1798),
.Y(net3626)
);

AOI21x1_ASAP7_75t_R c3603(
.A1(net1775),
.A2(net2620),
.B(net9733),
.Y(net3627)
);

OR2x6_ASAP7_75t_R c3604(
.A(net3433),
.B(net2463),
.Y(net3628)
);

BUFx12_ASAP7_75t_R c3605(
.A(net10524),
.Y(net3629)
);

XNOR2x1_ASAP7_75t_R c3606(
.B(net2619),
.A(net3599),
.Y(net3630)
);

XNOR2x2_ASAP7_75t_R c3607(
.A(net2620),
.B(net839),
.Y(net3631)
);

DFFASRHQNx1_ASAP7_75t_R c3608(
.D(net3623),
.RESETN(net3596),
.SETN(net3361),
.CLK(clk),
.QN(net3632)
);

XNOR2xp5_ASAP7_75t_R c3609(
.A(net3598),
.B(net3612),
.Y(net3633)
);

AOI21xp33_ASAP7_75t_R c3610(
.A1(net3615),
.A2(net3620),
.B(net849),
.Y(net3634)
);

SDFHx1_ASAP7_75t_R c3611(
.D(net3602),
.SE(net2671),
.SI(net2615),
.CLK(clk),
.QN(net3635)
);

XOR2x1_ASAP7_75t_R c3612(
.A(net3619),
.B(net9984),
.Y(net3636)
);

AOI21xp5_ASAP7_75t_R c3613(
.A1(net3510),
.A2(net3620),
.B(net3628),
.Y(net3637)
);

FAx1_ASAP7_75t_R c3614(
.A(net3630),
.B(net3632),
.CI(net2699),
.SN(net3638)
);

XOR2x2_ASAP7_75t_R c3615(
.A(net10160),
.B(net10217),
.Y(net3639)
);

BUFx12f_ASAP7_75t_R c3616(
.A(net10483),
.Y(net3640)
);

XOR2xp5_ASAP7_75t_R c3617(
.A(net3554),
.B(net10216),
.Y(net3641)
);

MAJIxp5_ASAP7_75t_R c3618(
.A(net2699),
.B(net2681),
.C(net3620),
.Y(net3642)
);

MAJx2_ASAP7_75t_R c3619(
.A(net2693),
.B(net3616),
.C(net9871),
.Y(net3643)
);

AND2x2_ASAP7_75t_R c3620(
.A(net1787),
.B(net2689),
.Y(net3644)
);

AND2x4_ASAP7_75t_R c3621(
.A(net849),
.B(net3580),
.Y(net3645)
);

AND2x6_ASAP7_75t_R c3622(
.A(net2681),
.B(net3640),
.Y(net3646)
);

HAxp5_ASAP7_75t_R c3623(
.A(net3614),
.B(net3641),
.CON(net3648),
.SN(net3647)
);

MAJx3_ASAP7_75t_R c3624(
.A(net1782),
.B(net3612),
.C(net3611),
.Y(net3649)
);

ICGx3_ASAP7_75t_R c3625(
.ENA(net3649),
.SE(net1769),
.CLK(clk),
.GCLK(net3650)
);

NAND2x1_ASAP7_75t_R c3626(
.A(net3519),
.B(net3640),
.Y(net3651)
);

NAND3x1_ASAP7_75t_R c3627(
.A(net2615),
.B(net3643),
.C(net3640),
.Y(net3652)
);

NAND2x1p5_ASAP7_75t_R c3628(
.A(net1652),
.B(net3651),
.Y(net3653)
);

NAND2x2_ASAP7_75t_R c3629(
.A(net1625),
.B(net2711),
.Y(net3654)
);

AO31x2_ASAP7_75t_R c3630(
.A1(net3625),
.A2(net3646),
.A3(net3635),
.B(net3361),
.Y(net3655)
);

ICGx4DC_ASAP7_75t_R c3631(
.ENA(net3637),
.SE(net3648),
.CLK(clk),
.GCLK(net3656)
);

NAND2xp33_ASAP7_75t_R c3632(
.A(net738),
.B(net2752),
.Y(net3657)
);

OAI33xp33_ASAP7_75t_R c3633(
.A1(net1794),
.A2(net3657),
.A3(net3635),
.B1(net824),
.B2(net2707),
.B3(net2747),
.Y(net3658)
);

AOI211x1_ASAP7_75t_R c3634(
.A1(net3651),
.A2(net3641),
.B(net3649),
.C(net3519),
.Y(net3659)
);

AOI211xp5_ASAP7_75t_R c3635(
.A1(net3634),
.A2(net3433),
.B(net2584),
.C(net3655),
.Y(net3660)
);

AOI22x1_ASAP7_75t_R c3636(
.A1(net3610),
.A2(net3648),
.B1(net1744),
.B2(net10230),
.Y(net3661)
);

AOI22xp33_ASAP7_75t_R c3637(
.A1(net2725),
.A2(net3631),
.B1(net2703),
.B2(net1802),
.Y(net3662)
);

NAND2xp5_ASAP7_75t_R c3638(
.A(net3657),
.B(net9899),
.Y(net3663)
);

NAND3x2_ASAP7_75t_R c3639(
.B(net3605),
.C(net3627),
.A(net3641),
.Y(net3664)
);

AOI22xp5_ASAP7_75t_R c3640(
.A1(net3651),
.A2(net3655),
.B1(net2708),
.B2(net9856),
.Y(net3665)
);

BUFx16f_ASAP7_75t_R c3641(
.A(net10330),
.Y(net3666)
);

NAND3xp33_ASAP7_75t_R c3642(
.A(net3594),
.B(net2736),
.C(net3619),
.Y(net3667)
);

AOI31xp33_ASAP7_75t_R c3643(
.A1(net3653),
.A2(net2719),
.A3(net3635),
.B(net10231),
.Y(net3668)
);

AOI31xp67_ASAP7_75t_R c3644(
.A1(net2672),
.A2(net3644),
.A3(net3640),
.B(net9856),
.Y(net3669)
);

NOR3x1_ASAP7_75t_R c3645(
.A(net3513),
.B(net3654),
.C(net3628),
.Y(net3670)
);

NAND4xp25_ASAP7_75t_R c3646(
.A(net3627),
.B(net3645),
.C(net1787),
.D(net10233),
.Y(net3671)
);

NAND4xp75_ASAP7_75t_R c3647(
.A(net3612),
.B(net3485),
.C(net10231),
.D(net10232),
.Y(net3672)
);

SDFHx2_ASAP7_75t_R c3648(
.D(net2716),
.SE(net3616),
.SI(net2729),
.CLK(clk),
.QN(net3673)
);

SDFHx3_ASAP7_75t_R c3649(
.D(net3669),
.SE(net3672),
.SI(net10232),
.CLK(clk),
.QN(net3674)
);

NOR4xp25_ASAP7_75t_R c3650(
.A(net3657),
.B(net3672),
.C(net3640),
.D(net10233),
.Y(net3675)
);

NOR3x2_ASAP7_75t_R c3651(
.B(net859),
.C(net686),
.A(net9922),
.Y(net3676)
);

BUFx24_ASAP7_75t_R c3652(
.A(net9164),
.Y(net3677)
);

BUFx2_ASAP7_75t_R c3653(
.A(net959),
.Y(net3678)
);

BUFx3_ASAP7_75t_R c3654(
.A(net9164),
.Y(net3679)
);

BUFx4_ASAP7_75t_R c3655(
.A(net2757),
.Y(net3680)
);

BUFx4f_ASAP7_75t_R c3656(
.A(net1864),
.Y(net3681)
);

ICGx4_ASAP7_75t_R c3657(
.ENA(net970),
.SE(net2819),
.CLK(clk),
.GCLK(net3682)
);

NAND2xp67_ASAP7_75t_R c3658(
.A(net3677),
.B(net3678),
.Y(net3683)
);

NOR2x1_ASAP7_75t_R c3659(
.A(net1839),
.B(net2777),
.Y(net3684)
);

BUFx5_ASAP7_75t_R c3660(
.A(net2819),
.Y(net3685)
);

BUFx6f_ASAP7_75t_R c3661(
.A(net3680),
.Y(net3686)
);

NOR2x1p5_ASAP7_75t_R c3662(
.A(net3686),
.B(net980),
.Y(net3687)
);

NOR2x2_ASAP7_75t_R c3663(
.A(net913),
.B(net3686),
.Y(net3688)
);

BUFx8_ASAP7_75t_R c3664(
.A(net2763),
.Y(net3689)
);

NOR2xp33_ASAP7_75t_R c3665(
.A(net1890),
.B(net2828),
.Y(net3690)
);

CKINVDCx10_ASAP7_75t_R c3666(
.A(net30),
.Y(net3691)
);

CKINVDCx11_ASAP7_75t_R c3667(
.A(net3677),
.Y(net3692)
);

NOR2xp67_ASAP7_75t_R c3668(
.A(net3683),
.B(net3689),
.Y(net3693)
);

CKINVDCx12_ASAP7_75t_R c3669(
.A(net3691),
.Y(net3694)
);

CKINVDCx14_ASAP7_75t_R c3670(
.A(net3678),
.Y(net3695)
);

OR2x2_ASAP7_75t_R c3671(
.A(net1904),
.B(net3683),
.Y(net3696)
);

CKINVDCx16_ASAP7_75t_R c3672(
.A(net9258),
.Y(net3697)
);

CKINVDCx20_ASAP7_75t_R c3673(
.A(net9258),
.Y(net3698)
);

CKINVDCx5p33_ASAP7_75t_R c3674(
.A(net950),
.Y(net3699)
);

CKINVDCx6p67_ASAP7_75t_R c3675(
.A(net3697),
.Y(net3700)
);

OR2x4_ASAP7_75t_R c3676(
.A(net3695),
.B(net3689),
.Y(net3701)
);

ICGx5_ASAP7_75t_R c3677(
.ENA(net3693),
.SE(net3685),
.CLK(clk),
.GCLK(net3702)
);

OR2x6_ASAP7_75t_R c3678(
.A(net3702),
.B(net2777),
.Y(net3703)
);

CKINVDCx8_ASAP7_75t_R c3679(
.A(net3692),
.Y(net3704)
);

CKINVDCx9p33_ASAP7_75t_R c3680(
.A(net1864),
.Y(net3705)
);

ICGx5p33DC_ASAP7_75t_R c3681(
.ENA(net2831),
.SE(net3692),
.CLK(clk),
.GCLK(net3706)
);

XNOR2x1_ASAP7_75t_R c3682(
.B(net3703),
.A(net1892),
.Y(net3707)
);

HB1xp67_ASAP7_75t_R c3683(
.A(net9279),
.Y(net3708)
);

HB2xp67_ASAP7_75t_R c3684(
.A(net2804),
.Y(net3709)
);

ICGx6p67DC_ASAP7_75t_R c3685(
.ENA(net3708),
.SE(net3701),
.CLK(clk),
.GCLK(net3710)
);

HB3xp67_ASAP7_75t_R c3686(
.A(net1891),
.Y(net3711)
);

ICGx8DC_ASAP7_75t_R c3687(
.ENA(net2759),
.SE(net3696),
.CLK(clk),
.GCLK(net3712)
);

HB4xp67_ASAP7_75t_R c3688(
.A(net9286),
.Y(net3713)
);

INVx11_ASAP7_75t_R c3689(
.A(net3704),
.Y(net3714)
);

ICGx1_ASAP7_75t_R c3690(
.ENA(net3686),
.SE(net3693),
.CLK(clk),
.GCLK(net3715)
);

INVx13_ASAP7_75t_R c3691(
.A(net3715),
.Y(net3716)
);

INVx1_ASAP7_75t_R c3692(
.A(net3712),
.Y(net3717)
);

INVx2_ASAP7_75t_R c3693(
.A(net3717),
.Y(net3718)
);

XNOR2x2_ASAP7_75t_R c3694(
.A(net900),
.B(net3691),
.Y(net3719)
);

INVx3_ASAP7_75t_R c3695(
.A(net9286),
.Y(net3720)
);

INVx4_ASAP7_75t_R c3696(
.A(net3698),
.Y(net3721)
);

INVx5_ASAP7_75t_R c3697(
.A(net3700),
.Y(net3722)
);

INVx6_ASAP7_75t_R c3698(
.A(net9713),
.Y(net3723)
);

XNOR2xp5_ASAP7_75t_R c3699(
.A(net1884),
.B(net3705),
.Y(net3724)
);

XOR2x1_ASAP7_75t_R c3700(
.A(net3721),
.B(net2763),
.Y(net3725)
);

INVx8_ASAP7_75t_R c3701(
.A(net3715),
.Y(net3726)
);

NOR3xp33_ASAP7_75t_R c3702(
.A(net2777),
.B(net3712),
.C(net3699),
.Y(net3727)
);

XOR2x2_ASAP7_75t_R c3703(
.A(net3691),
.B(net3709),
.Y(net3728)
);

SDFHx4_ASAP7_75t_R c3704(
.D(net2812),
.SE(net3724),
.SI(net3704),
.CLK(clk),
.QN(net3729)
);

INVxp33_ASAP7_75t_R c3705(
.A(net3723),
.Y(net3730)
);

INVxp67_ASAP7_75t_R c3706(
.A(net3719),
.Y(net3731)
);

BUFx10_ASAP7_75t_R c3707(
.A(net3687),
.Y(net3732)
);

XOR2xp5_ASAP7_75t_R c3708(
.A(net3722),
.B(net3718),
.Y(net3733)
);

BUFx12_ASAP7_75t_R c3709(
.A(net9713),
.Y(net3734)
);

AO222x2_ASAP7_75t_R c3710(
.A1(net3718),
.A2(net3721),
.B1(net3703),
.B2(net3708),
.C1(net3699),
.C2(net2763),
.Y(net3735)
);

AND2x2_ASAP7_75t_R c3711(
.A(net3718),
.B(net3704),
.Y(net3736)
);

AO33x2_ASAP7_75t_R c3712(
.A1(net3689),
.A2(net3717),
.A3(net3682),
.B1(net2777),
.B2(net3701),
.B3(net3699),
.Y(net3737)
);

BUFx12f_ASAP7_75t_R c3713(
.A(net3716),
.Y(net3738)
);

AND2x4_ASAP7_75t_R c3714(
.A(net3730),
.B(net3711),
.Y(net3739)
);

BUFx16f_ASAP7_75t_R c3715(
.A(net9310),
.Y(net3740)
);

BUFx24_ASAP7_75t_R c3716(
.A(net3736),
.Y(net3741)
);

OA21x2_ASAP7_75t_R c3717(
.A1(net3740),
.A2(net3709),
.B(net3713),
.Y(net3742)
);

AND2x6_ASAP7_75t_R c3718(
.A(net3734),
.B(net3715),
.Y(net3743)
);

BUFx2_ASAP7_75t_R c3719(
.A(net9279),
.Y(net3744)
);

HAxp5_ASAP7_75t_R c3720(
.A(net3735),
.B(net2777),
.CON(net3746),
.SN(net3745)
);

NAND2x1_ASAP7_75t_R c3721(
.A(net3681),
.B(net3722),
.Y(net3747)
);

NAND2x1p5_ASAP7_75t_R c3722(
.A(net2825),
.B(net3701),
.Y(net3748)
);

OAI21x1_ASAP7_75t_R c3723(
.A1(net3724),
.A2(net2804),
.B(net2812),
.Y(net3749)
);

NAND2x2_ASAP7_75t_R c3724(
.A(net3727),
.B(net3713),
.Y(net3750)
);

ICGx2_ASAP7_75t_R c3725(
.ENA(net3719),
.SE(net3731),
.CLK(clk),
.GCLK(net3751)
);

BUFx3_ASAP7_75t_R c3726(
.A(net3732),
.Y(net3752)
);

BUFx4_ASAP7_75t_R c3727(
.A(net3729),
.Y(net3753)
);

NAND2xp33_ASAP7_75t_R c3728(
.A(net3691),
.B(net9857),
.Y(net3754)
);

OAI21xp33_ASAP7_75t_R c3729(
.A1(net3738),
.A2(net3714),
.B(net2792),
.Y(net3755)
);

NAND2xp5_ASAP7_75t_R c3730(
.A(net3742),
.B(net3745),
.Y(net3756)
);

NAND2xp67_ASAP7_75t_R c3731(
.A(net3744),
.B(net3752),
.Y(net3757)
);

OAI21xp5_ASAP7_75t_R c3732(
.A1(net3757),
.A2(net3735),
.B(net3729),
.Y(net3758)
);

NOR2x1_ASAP7_75t_R c3733(
.A(net3750),
.B(net9857),
.Y(net3759)
);

NOR2x1p5_ASAP7_75t_R c3734(
.A(net3756),
.B(net3747),
.Y(net3760)
);

BUFx4f_ASAP7_75t_R c3735(
.A(net2897),
.Y(net3761)
);

NOR2x2_ASAP7_75t_R c3736(
.A(net2919),
.B(net3731),
.Y(net3762)
);

BUFx5_ASAP7_75t_R c3737(
.A(net1962),
.Y(net3763)
);

NOR2xp33_ASAP7_75t_R c3738(
.A(net2900),
.B(net1962),
.Y(net3764)
);

BUFx6f_ASAP7_75t_R c3739(
.A(net2867),
.Y(net3765)
);

BUFx8_ASAP7_75t_R c3740(
.A(net10497),
.Y(net3766)
);

OR3x1_ASAP7_75t_R c3741(
.A(net2811),
.B(net2899),
.C(net10220),
.Y(net3767)
);

NOR2xp67_ASAP7_75t_R c3742(
.A(net1948),
.B(net900),
.Y(net3768)
);

OR3x2_ASAP7_75t_R c3743(
.A(net3743),
.B(net2900),
.C(net1948),
.Y(net3769)
);

CKINVDCx10_ASAP7_75t_R c3744(
.A(net3754),
.Y(net3770)
);

CKINVDCx11_ASAP7_75t_R c3745(
.A(net9142),
.Y(net3771)
);

ICGx2p67DC_ASAP7_75t_R c3746(
.ENA(net3711),
.SE(net1848),
.CLK(clk),
.GCLK(net3772)
);

ICGx3_ASAP7_75t_R c3747(
.ENA(net3769),
.SE(net2882),
.CLK(clk),
.GCLK(net3773)
);

OR2x2_ASAP7_75t_R c3748(
.A(net2870),
.B(net3711),
.Y(net3774)
);

OR2x4_ASAP7_75t_R c3749(
.A(net3770),
.B(net2829),
.Y(net3775)
);

OR2x6_ASAP7_75t_R c3750(
.A(net3720),
.B(net2823),
.Y(net3776)
);

XNOR2x1_ASAP7_75t_R c3751(
.B(net3763),
.A(net2867),
.Y(net3777)
);

CKINVDCx12_ASAP7_75t_R c3752(
.A(net10235),
.Y(net3778)
);

CKINVDCx14_ASAP7_75t_R c3753(
.A(net9729),
.Y(net3779)
);

CKINVDCx16_ASAP7_75t_R c3754(
.A(net10189),
.Y(net3780)
);

OR3x4_ASAP7_75t_R c3755(
.A(net1991),
.B(net2870),
.C(net10187),
.Y(net3781)
);

CKINVDCx20_ASAP7_75t_R c3756(
.A(net9954),
.Y(net3782)
);

AND3x1_ASAP7_75t_R c3757(
.A(net3773),
.B(net3761),
.C(net3758),
.Y(net3783)
);

AND3x2_ASAP7_75t_R c3758(
.A(net2882),
.B(net2896),
.C(net3776),
.Y(net3784)
);

CKINVDCx5p33_ASAP7_75t_R c3759(
.A(net3750),
.Y(net3785)
);

XNOR2x2_ASAP7_75t_R c3760(
.A(net3761),
.B(net9758),
.Y(net3786)
);

CKINVDCx6p67_ASAP7_75t_R c3761(
.A(net2848),
.Y(net3787)
);

XNOR2xp5_ASAP7_75t_R c3762(
.A(net1970),
.B(net3776),
.Y(net3788)
);

CKINVDCx8_ASAP7_75t_R c3763(
.A(net2896),
.Y(net3789)
);

CKINVDCx9p33_ASAP7_75t_R c3764(
.A(net3752),
.Y(net3790)
);

XOR2x1_ASAP7_75t_R c3765(
.A(net3679),
.B(net3772),
.Y(net3791)
);

HB1xp67_ASAP7_75t_R c3766(
.A(net1911),
.Y(net3792)
);

HB2xp67_ASAP7_75t_R c3767(
.A(net3785),
.Y(net3793)
);

XOR2x2_ASAP7_75t_R c3768(
.A(net3783),
.B(net9935),
.Y(net3794)
);

AND3x4_ASAP7_75t_R c3769(
.A(net2855),
.B(net3777),
.C(net2896),
.Y(net3795)
);

XOR2xp5_ASAP7_75t_R c3770(
.A(net3784),
.B(net3794),
.Y(net3796)
);

AND2x2_ASAP7_75t_R c3771(
.A(net3787),
.B(net3750),
.Y(net3797)
);

HB3xp67_ASAP7_75t_R c3772(
.A(net3782),
.Y(net3798)
);

AND2x4_ASAP7_75t_R c3773(
.A(net2884),
.B(net2896),
.Y(net3799)
);

AND2x6_ASAP7_75t_R c3774(
.A(net3794),
.B(net3799),
.Y(net3800)
);

HB4xp67_ASAP7_75t_R c3775(
.A(net3791),
.Y(net3801)
);

HAxp5_ASAP7_75t_R c3776(
.A(net3798),
.B(net3682),
.CON(net3803),
.SN(net3802)
);

INVx11_ASAP7_75t_R c3777(
.A(net10163),
.Y(net3804)
);

NOR4xp75_ASAP7_75t_R c3778(
.A(net3799),
.B(net3739),
.C(net2810),
.D(net3758),
.Y(net3805)
);

NAND2x1_ASAP7_75t_R c3779(
.A(net980),
.B(net3784),
.Y(net3806)
);

AO21x1_ASAP7_75t_R c3780(
.A1(net1848),
.A2(net3680),
.B(net1856),
.Y(net3807)
);

INVx13_ASAP7_75t_R c3781(
.A(net3803),
.Y(net3808)
);

INVx1_ASAP7_75t_R c3782(
.A(net3797),
.Y(net3809)
);

ICGx4DC_ASAP7_75t_R c3783(
.ENA(net3769),
.SE(net2848),
.CLK(clk),
.GCLK(net3810)
);

INVx2_ASAP7_75t_R c3784(
.A(net9142),
.Y(net3811)
);

NAND2x1p5_ASAP7_75t_R c3785(
.A(net2823),
.B(net9786),
.Y(net3812)
);

NAND2x2_ASAP7_75t_R c3786(
.A(net79),
.B(net3805),
.Y(net3813)
);

INVx3_ASAP7_75t_R c3787(
.A(net10542),
.Y(net3814)
);

INVx4_ASAP7_75t_R c3788(
.A(net3771),
.Y(net3815)
);

INVx5_ASAP7_75t_R c3789(
.A(net3814),
.Y(net3816)
);

NAND2xp33_ASAP7_75t_R c3790(
.A(net3801),
.B(net3794),
.Y(net3817)
);

O2A1O1Ixp33_ASAP7_75t_R c3791(
.A1(net1839),
.A2(net3812),
.B(net2866),
.C(net3772),
.Y(net3818)
);

NAND2xp5_ASAP7_75t_R c3792(
.A(net3811),
.B(net9729),
.Y(net3819)
);

AO21x2_ASAP7_75t_R c3793(
.A1(net2847),
.A2(net2848),
.B(net10236),
.Y(net3820)
);

NAND2xp67_ASAP7_75t_R c3794(
.A(net2757),
.B(net3699),
.Y(net3821)
);

AOI21x1_ASAP7_75t_R c3795(
.A1(net3806),
.A2(net3815),
.B(net10235),
.Y(net3822)
);

O2A1O1Ixp5_ASAP7_75t_R c3796(
.A1(net3812),
.A2(net3814),
.B(net3805),
.C(net3701),
.Y(net3823)
);

INVx6_ASAP7_75t_R c3797(
.A(net10575),
.Y(net3824)
);

NOR2x1_ASAP7_75t_R c3798(
.A(net3761),
.B(net3794),
.Y(net3825)
);

AOI21xp33_ASAP7_75t_R c3799(
.A1(net3779),
.A2(net3810),
.B(net3777),
.Y(net3826)
);

NOR2x1p5_ASAP7_75t_R c3800(
.A(net3780),
.B(net3791),
.Y(net3827)
);

AOI222xp33_ASAP7_75t_R c3801(
.A1(net3816),
.A2(net3791),
.B1(net3781),
.B2(net3789),
.C1(net1971),
.C2(net2918),
.Y(net3828)
);

INVx8_ASAP7_75t_R c3802(
.A(net10496),
.Y(net3829)
);

AOI21xp5_ASAP7_75t_R c3803(
.A1(net3789),
.A2(net9786),
.B(net10220),
.Y(net3830)
);

ICGx4_ASAP7_75t_R c3804(
.ENA(net3796),
.SE(net3802),
.CLK(clk),
.GCLK(net3831)
);

NOR2x2_ASAP7_75t_R c3805(
.A(net3819),
.B(net3773),
.Y(net3832)
);

NOR2xp33_ASAP7_75t_R c3806(
.A(net3829),
.B(net10237),
.Y(net3833)
);

NOR2xp67_ASAP7_75t_R c3807(
.A(net2865),
.B(net2897),
.Y(net3834)
);

OR2x2_ASAP7_75t_R c3808(
.A(net3822),
.B(net3766),
.Y(net3835)
);

INVxp33_ASAP7_75t_R c3809(
.A(net9825),
.Y(net3836)
);

OR2x4_ASAP7_75t_R c3810(
.A(net959),
.B(net3789),
.Y(net3837)
);

OR2x6_ASAP7_75t_R c3811(
.A(net3837),
.B(net3771),
.Y(net3838)
);

FAx1_ASAP7_75t_R c3812(
.A(net3833),
.B(net3831),
.CI(net3805),
.SN(net3840),
.CON(net3839)
);

MAJIxp5_ASAP7_75t_R c3813(
.A(net3820),
.B(net3752),
.C(net3835),
.Y(net3841)
);

MAJx2_ASAP7_75t_R c3814(
.A(net3824),
.B(net3835),
.C(net3839),
.Y(net3842)
);

MAJx3_ASAP7_75t_R c3815(
.A(net2913),
.B(net3839),
.C(net9745),
.Y(net3843)
);

XNOR2x1_ASAP7_75t_R c3816(
.B(net3786),
.A(net9978),
.Y(net3844)
);

NAND3x1_ASAP7_75t_R c3817(
.A(net3831),
.B(net3810),
.C(net9978),
.Y(net3845)
);

INVxp67_ASAP7_75t_R c3818(
.A(net9257),
.Y(net3846)
);

XNOR2x2_ASAP7_75t_R c3819(
.A(net2971),
.B(net2052),
.Y(net3847)
);

XNOR2xp5_ASAP7_75t_R c3820(
.A(net2914),
.B(net2996),
.Y(net3848)
);

XOR2x1_ASAP7_75t_R c3821(
.A(net1118),
.B(net2045),
.Y(net3849)
);

XOR2x2_ASAP7_75t_R c3822(
.A(net2953),
.B(net3840),
.Y(net3850)
);

XOR2xp5_ASAP7_75t_R c3823(
.A(net2899),
.B(net10047),
.Y(net3851)
);

AND2x2_ASAP7_75t_R c3824(
.A(net1119),
.B(net2918),
.Y(net3852)
);

AND2x4_ASAP7_75t_R c3825(
.A(net2970),
.B(net1089),
.Y(net3853)
);

BUFx10_ASAP7_75t_R c3826(
.A(net3753),
.Y(net3854)
);

AND2x6_ASAP7_75t_R c3827(
.A(net1137),
.B(net3831),
.Y(net3855)
);

BUFx12_ASAP7_75t_R c3828(
.A(net3840),
.Y(net3856)
);

HAxp5_ASAP7_75t_R c3829(
.A(net1089),
.B(net3804),
.CON(net3858),
.SN(net3857)
);

NAND2x1_ASAP7_75t_R c3830(
.A(net3858),
.B(net2842),
.Y(net3859)
);

NAND2x1p5_ASAP7_75t_R c3831(
.A(net1980),
.B(net2036),
.Y(net3860)
);

BUFx12f_ASAP7_75t_R c3832(
.A(net9693),
.Y(net3861)
);

BUFx16f_ASAP7_75t_R c3833(
.A(net9149),
.Y(net3862)
);

BUFx24_ASAP7_75t_R c3834(
.A(net3860),
.Y(net3863)
);

BUFx2_ASAP7_75t_R c3835(
.A(net10479),
.Y(net3864)
);

NAND2x2_ASAP7_75t_R c3836(
.A(net3832),
.B(net3835),
.Y(net3865)
);

BUFx3_ASAP7_75t_R c3837(
.A(net10136),
.Y(net3866)
);

NAND2xp33_ASAP7_75t_R c3838(
.A(net3805),
.B(net2842),
.Y(net3867)
);

NAND2xp5_ASAP7_75t_R c3839(
.A(net3851),
.B(net3741),
.Y(net3868)
);

BUFx4_ASAP7_75t_R c3840(
.A(net10016),
.Y(net3869)
);

BUFx4f_ASAP7_75t_R c3841(
.A(net9149),
.Y(net3870)
);

NAND2xp67_ASAP7_75t_R c3842(
.A(net1833),
.B(net9758),
.Y(net3871)
);

ICGx5_ASAP7_75t_R c3843(
.ENA(net3831),
.SE(net3835),
.CLK(clk),
.GCLK(net3872)
);

BUFx5_ASAP7_75t_R c3844(
.A(net9267),
.Y(net3873)
);

NOR2x1_ASAP7_75t_R c3845(
.A(net3871),
.B(net10113),
.Y(net3874)
);

NOR2x1p5_ASAP7_75t_R c3846(
.A(net3869),
.B(net3707),
.Y(net3875)
);

BUFx6f_ASAP7_75t_R c3847(
.A(net9980),
.Y(net3876)
);

NOR2x2_ASAP7_75t_R c3848(
.A(net2927),
.B(net3872),
.Y(net3877)
);

ICGx5p33DC_ASAP7_75t_R c3849(
.ENA(net3875),
.SE(net2999),
.CLK(clk),
.GCLK(net3878)
);

NAND3x2_ASAP7_75t_R c3850(
.B(net3758),
.C(net3741),
.A(net3766),
.Y(net3879)
);

NOR2xp33_ASAP7_75t_R c3851(
.A(net3874),
.B(net3863),
.Y(net3880)
);

SDFLx1_ASAP7_75t_R c3852(
.D(net1971),
.SE(net3699),
.SI(net2918),
.CLK(clk),
.QN(net3881)
);

NAND3xp33_ASAP7_75t_R c3853(
.A(net3876),
.B(net3879),
.C(net3871),
.Y(net3882)
);

BUFx8_ASAP7_75t_R c3854(
.A(net3847),
.Y(net3883)
);

NOR2xp67_ASAP7_75t_R c3855(
.A(net3864),
.B(net3867),
.Y(net3884)
);

NOR3x1_ASAP7_75t_R c3856(
.A(net3866),
.B(net3854),
.C(net3783),
.Y(net3885)
);

OR2x2_ASAP7_75t_R c3857(
.A(net2014),
.B(net3849),
.Y(net3886)
);

OR2x4_ASAP7_75t_R c3858(
.A(net3858),
.B(net3881),
.Y(net3887)
);

CKINVDCx10_ASAP7_75t_R c3859(
.A(net3885),
.Y(net3888)
);

NOR3x2_ASAP7_75t_R c3860(
.B(net3861),
.C(net3868),
.A(net3870),
.Y(net3889)
);

NOR3xp33_ASAP7_75t_R c3861(
.A(net3862),
.B(net3849),
.C(net3778),
.Y(net3890)
);

OR2x6_ASAP7_75t_R c3862(
.A(net3811),
.B(net3790),
.Y(net3891)
);

CKINVDCx11_ASAP7_75t_R c3863(
.A(net9980),
.Y(net3892)
);

CKINVDCx12_ASAP7_75t_R c3864(
.A(net3866),
.Y(net3893)
);

CKINVDCx14_ASAP7_75t_R c3865(
.A(net9969),
.Y(net3894)
);

ICGx6p67DC_ASAP7_75t_R c3866(
.ENA(net3888),
.SE(net2829),
.CLK(clk),
.GCLK(net3895)
);

XNOR2x1_ASAP7_75t_R c3867(
.B(net3882),
.A(net3861),
.Y(net3896)
);

XNOR2x2_ASAP7_75t_R c3868(
.A(net3849),
.B(net3892),
.Y(net3897)
);

XNOR2xp5_ASAP7_75t_R c3869(
.A(net3778),
.B(net10096),
.Y(net3898)
);

CKINVDCx16_ASAP7_75t_R c3870(
.A(net9992),
.Y(net3899)
);

XOR2x1_ASAP7_75t_R c3871(
.A(net3897),
.B(net3876),
.Y(net3900)
);

CKINVDCx20_ASAP7_75t_R c3872(
.A(net10088),
.Y(net3901)
);

CKINVDCx5p33_ASAP7_75t_R c3873(
.A(net10096),
.Y(net3902)
);

CKINVDCx6p67_ASAP7_75t_R c3874(
.A(net10136),
.Y(net3903)
);

OA21x2_ASAP7_75t_R c3875(
.A1(net3741),
.A2(net3886),
.B(net3903),
.Y(net3904)
);

XOR2x2_ASAP7_75t_R c3876(
.A(net3891),
.B(net3741),
.Y(net3905)
);

OAI21x1_ASAP7_75t_R c3877(
.A1(net3902),
.A2(net2954),
.B(net3892),
.Y(net3906)
);

XOR2xp5_ASAP7_75t_R c3878(
.A(net3804),
.B(net10016),
.Y(net3907)
);

OAI21xp33_ASAP7_75t_R c3879(
.A1(net2811),
.A2(net3813),
.B(net3893),
.Y(net3908)
);

AND5x1_ASAP7_75t_R c3880(
.A(net3844),
.B(net3902),
.C(net3768),
.D(net3856),
.E(net3872),
.Y(net3909)
);

AND2x2_ASAP7_75t_R c3881(
.A(net3898),
.B(net3758),
.Y(net3910)
);

OAI21xp5_ASAP7_75t_R c3882(
.A1(net3910),
.A2(net2036),
.B(net2970),
.Y(net3911)
);

OR3x1_ASAP7_75t_R c3883(
.A(net2956),
.B(net3861),
.C(net3893),
.Y(net3912)
);

CKINVDCx8_ASAP7_75t_R c3884(
.A(net10567),
.Y(net3913)
);

AND2x4_ASAP7_75t_R c3885(
.A(net3883),
.B(net3857),
.Y(net3914)
);

OR3x2_ASAP7_75t_R c3886(
.A(net3913),
.B(net3910),
.C(net1138),
.Y(net3915)
);

AND2x6_ASAP7_75t_R c3887(
.A(net3907),
.B(net3881),
.Y(net3916)
);

OR3x4_ASAP7_75t_R c3888(
.A(net3881),
.B(net2899),
.C(net3874),
.Y(net3917)
);

AOI321xp33_ASAP7_75t_R c3889(
.A1(net3850),
.A2(net2942),
.A3(net3893),
.B1(net2991),
.B2(net2918),
.C(net10138),
.Y(net3918)
);

SDFLx2_ASAP7_75t_R c3890(
.D(net2999),
.SE(net3894),
.SI(net10237),
.CLK(clk),
.QN(net3919)
);

SDFLx3_ASAP7_75t_R c3891(
.D(net3915),
.SE(net3862),
.SI(net3850),
.CLK(clk),
.QN(net3920)
);

CKINVDCx9p33_ASAP7_75t_R c3892(
.A(net10529),
.Y(net3921)
);

AND3x1_ASAP7_75t_R c3893(
.A(net3880),
.B(net2811),
.C(net3917),
.Y(net3922)
);

HAxp5_ASAP7_75t_R c3894(
.A(net3921),
.B(net10138),
.CON(net3924),
.SN(net3923)
);

AND5x2_ASAP7_75t_R c3895(
.A(net3894),
.B(net3893),
.C(net3875),
.D(net3846),
.E(net2045),
.Y(net3925)
);

AND3x2_ASAP7_75t_R c3896(
.A(net2934),
.B(net3923),
.C(net10238),
.Y(net3926)
);

AO221x1_ASAP7_75t_R c3897(
.A1(net3879),
.A2(net3917),
.B1(net3924),
.B2(net3872),
.C(net3772),
.Y(net3927)
);

OA211x2_ASAP7_75t_R c3898(
.A1(net3889),
.A2(net3890),
.B(net3805),
.C(net10238),
.Y(net3928)
);

NAND2x1_ASAP7_75t_R c3899(
.A(net3916),
.B(net10238),
.Y(net3929)
);

AND3x4_ASAP7_75t_R c3900(
.A(net3919),
.B(net3929),
.C(net9807),
.Y(net3930)
);

NAND2x1p5_ASAP7_75t_R c3901(
.A(net2989),
.B(net3930),
.Y(net3931)
);

NAND2x2_ASAP7_75t_R c3902(
.A(net3905),
.B(net10236),
.Y(net3932)
);

HB1xp67_ASAP7_75t_R c3903(
.A(net9973),
.Y(net3933)
);

HB2xp67_ASAP7_75t_R c3904(
.A(net10510),
.Y(net3934)
);

NAND2xp33_ASAP7_75t_R c3905(
.A(net2036),
.B(net3086),
.Y(net3935)
);

HB3xp67_ASAP7_75t_R c3906(
.A(net3870),
.Y(net3936)
);

NAND2xp5_ASAP7_75t_R c3907(
.A(net87),
.B(net1933),
.Y(net3937)
);

NAND2xp67_ASAP7_75t_R c3908(
.A(net1077),
.B(net3895),
.Y(net3938)
);

HB4xp67_ASAP7_75t_R c3909(
.A(net10158),
.Y(net3939)
);

NOR2x1_ASAP7_75t_R c3910(
.A(net2997),
.B(net3013),
.Y(net3940)
);

NOR2x1p5_ASAP7_75t_R c3911(
.A(net1861),
.B(net10236),
.Y(net3941)
);

NOR2x2_ASAP7_75t_R c3912(
.A(net1933),
.B(net3073),
.Y(net3942)
);

INVx11_ASAP7_75t_R c3913(
.A(net3932),
.Y(net3943)
);

INVx13_ASAP7_75t_R c3914(
.A(net10553),
.Y(net3944)
);

NOR2xp33_ASAP7_75t_R c3915(
.A(net3089),
.B(net2984),
.Y(net3945)
);

NOR2xp67_ASAP7_75t_R c3916(
.A(net3853),
.B(net2962),
.Y(net3946)
);

INVx1_ASAP7_75t_R c3917(
.A(net10066),
.Y(net3947)
);

OR2x2_ASAP7_75t_R c3918(
.A(net3024),
.B(net3707),
.Y(net3948)
);

OR2x4_ASAP7_75t_R c3919(
.A(net2918),
.B(net3867),
.Y(net3949)
);

OR2x6_ASAP7_75t_R c3920(
.A(net1991),
.B(net3920),
.Y(net3950)
);

AO21x1_ASAP7_75t_R c3921(
.A1(net2991),
.A2(net1991),
.B(net3783),
.Y(net3951)
);

AO21x2_ASAP7_75t_R c3922(
.A1(net3934),
.A2(net3710),
.B(net2153),
.Y(net3952)
);

AOI33xp33_ASAP7_75t_R c3923(
.A1(net2921),
.A2(net3942),
.A3(net1077),
.B1(net1991),
.B2(net3950),
.B3(net3066),
.Y(net3953)
);

ICGx8DC_ASAP7_75t_R c3924(
.ENA(net2938),
.SE(net3943),
.CLK(clk),
.GCLK(net3954)
);

XNOR2x1_ASAP7_75t_R c3925(
.B(net3937),
.A(net3947),
.Y(net3955)
);

XNOR2x2_ASAP7_75t_R c3926(
.A(net3048),
.B(net3950),
.Y(net3956)
);

XNOR2xp5_ASAP7_75t_R c3927(
.A(net3846),
.B(net9741),
.Y(net3957)
);

XOR2x1_ASAP7_75t_R c3928(
.A(net3954),
.B(net3710),
.Y(net3958)
);

XOR2x2_ASAP7_75t_R c3929(
.A(net3944),
.B(net3782),
.Y(net3959)
);

XOR2xp5_ASAP7_75t_R c3930(
.A(net3959),
.B(net10239),
.Y(net3960)
);

AOI21x1_ASAP7_75t_R c3931(
.A1(net3954),
.A2(net2842),
.B(net3950),
.Y(net3961)
);

AND2x2_ASAP7_75t_R c3932(
.A(net3945),
.B(net3867),
.Y(net3962)
);

AOI21xp33_ASAP7_75t_R c3933(
.A1(net3960),
.A2(net10236),
.B(net10239),
.Y(net3963)
);

AOI21xp5_ASAP7_75t_R c3934(
.A1(net3001),
.A2(net1915),
.B(net3963),
.Y(net3964)
);

INVx2_ASAP7_75t_R c3935(
.A(net10079),
.Y(net3965)
);

INVx3_ASAP7_75t_R c3936(
.A(net2121),
.Y(net3966)
);

AND2x4_ASAP7_75t_R c3937(
.A(net3931),
.B(net2997),
.Y(net3967)
);

AND2x6_ASAP7_75t_R c3938(
.A(net3958),
.B(net3957),
.Y(net3968)
);

HAxp5_ASAP7_75t_R c3939(
.A(net2891),
.B(net2899),
.CON(net3970),
.SN(net3969)
);

FAx1_ASAP7_75t_R c3940(
.A(net3887),
.B(net1163),
.CI(net3892),
.SN(net3971)
);

INVx4_ASAP7_75t_R c3941(
.A(net10163),
.Y(net3972)
);

NAND2x1_ASAP7_75t_R c3942(
.A(net3966),
.B(net1059),
.Y(net3973)
);

NAND2x1p5_ASAP7_75t_R c3943(
.A(net3948),
.B(net10239),
.Y(net3974)
);

INVx5_ASAP7_75t_R c3944(
.A(net10554),
.Y(net3975)
);

INVx6_ASAP7_75t_R c3945(
.A(net10066),
.Y(net3976)
);

NAND2x2_ASAP7_75t_R c3946(
.A(net3975),
.B(net3039),
.Y(net3977)
);

NAND2xp33_ASAP7_75t_R c3947(
.A(net3976),
.B(net3963),
.Y(net3978)
);

NAND2xp5_ASAP7_75t_R c3948(
.A(net3947),
.B(net2090),
.Y(net3979)
);

NAND2xp67_ASAP7_75t_R c3949(
.A(net3968),
.B(net3978),
.Y(net3980)
);

NOR2x1_ASAP7_75t_R c3950(
.A(net3978),
.B(net3958),
.Y(net3981)
);

INVx8_ASAP7_75t_R c3951(
.A(net10019),
.Y(net3982)
);

NOR2x1p5_ASAP7_75t_R c3952(
.A(net3033),
.B(net3965),
.Y(net3983)
);

NOR2x2_ASAP7_75t_R c3953(
.A(net3899),
.B(net3838),
.Y(net3984)
);

SDFLx4_ASAP7_75t_R c3954(
.D(net3981),
.SE(net3950),
.SI(net3049),
.CLK(clk),
.QN(net3985)
);

NOR2xp33_ASAP7_75t_R c3955(
.A(net3013),
.B(net3985),
.Y(net3986)
);

NOR2xp67_ASAP7_75t_R c3956(
.A(net3082),
.B(net10095),
.Y(net3987)
);

OR2x2_ASAP7_75t_R c3957(
.A(net3982),
.B(net3870),
.Y(net3988)
);

MAJIxp5_ASAP7_75t_R c3958(
.A(net3980),
.B(net3979),
.C(net3954),
.Y(net3989)
);

INVxp33_ASAP7_75t_R c3959(
.A(net9954),
.Y(net3990)
);

INVxp67_ASAP7_75t_R c3960(
.A(net10070),
.Y(net3991)
);

OR2x4_ASAP7_75t_R c3961(
.A(net3979),
.B(net3867),
.Y(net3992)
);

BUFx10_ASAP7_75t_R c3962(
.A(net10091),
.Y(net3993)
);

OR2x6_ASAP7_75t_R c3963(
.A(net3974),
.B(net3760),
.Y(net3994)
);

MAJx2_ASAP7_75t_R c3964(
.A(net3993),
.B(net3933),
.C(net2095),
.Y(net3995)
);

XNOR2x1_ASAP7_75t_R c3965(
.B(net3082),
.A(net3976),
.Y(net3996)
);

XNOR2x2_ASAP7_75t_R c3966(
.A(net2899),
.B(net3991),
.Y(net3997)
);

MAJx3_ASAP7_75t_R c3967(
.A(net3986),
.B(net3958),
.C(net3996),
.Y(net3998)
);

NAND3x1_ASAP7_75t_R c3968(
.A(net3972),
.B(net3981),
.C(net3976),
.Y(net3999)
);

XNOR2xp5_ASAP7_75t_R c3969(
.A(net3965),
.B(net3988),
.Y(net4000)
);

XOR2x1_ASAP7_75t_R c3970(
.A(net3851),
.B(net3980),
.Y(net4001)
);

XOR2x2_ASAP7_75t_R c3971(
.A(net3872),
.B(net9806),
.Y(net4002)
);

BUFx12_ASAP7_75t_R c3972(
.A(net10079),
.Y(net4003)
);

NAND3x2_ASAP7_75t_R c3973(
.B(net3999),
.C(net2045),
.A(net4002),
.Y(net4004)
);

NAND3xp33_ASAP7_75t_R c3974(
.A(net3935),
.B(net1211),
.C(net3996),
.Y(net4005)
);

OA222x2_ASAP7_75t_R c3975(
.A1(net3940),
.A2(net2149),
.B1(net3980),
.B2(net3942),
.C1(net3941),
.C2(net3950),
.Y(net4006)
);

XOR2xp5_ASAP7_75t_R c3976(
.A(net3967),
.B(net3980),
.Y(net4007)
);

NOR3x1_ASAP7_75t_R c3977(
.A(net4004),
.B(net3922),
.C(net3992),
.Y(net4008)
);

BUFx12f_ASAP7_75t_R c3978(
.A(net10079),
.Y(net4009)
);

NOR3x2_ASAP7_75t_R c3979(
.B(net3966),
.C(net4009),
.A(net10023),
.Y(net4010)
);

BUFx16f_ASAP7_75t_R c3980(
.A(net10399),
.Y(net4011)
);

NOR3xp33_ASAP7_75t_R c3981(
.A(net270),
.B(net3999),
.C(net3996),
.Y(net4012)
);

BUFx24_ASAP7_75t_R c3982(
.A(net10158),
.Y(net4013)
);

OA21x2_ASAP7_75t_R c3983(
.A1(net3991),
.A2(net4003),
.B(net9860),
.Y(net4014)
);

AND2x2_ASAP7_75t_R c3984(
.A(net3039),
.B(net3783),
.Y(net4015)
);

BUFx2_ASAP7_75t_R c3985(
.A(net3170),
.Y(net4016)
);

BUFx3_ASAP7_75t_R c3986(
.A(net9967),
.Y(net4017)
);

AO221x2_ASAP7_75t_R c3987(
.A1(net3985),
.A2(net4016),
.B1(net3895),
.B2(net3943),
.C(net1160),
.Y(net4018)
);

BUFx4_ASAP7_75t_R c3988(
.A(net10562),
.Y(net4019)
);

AND2x4_ASAP7_75t_R c3989(
.A(net2034),
.B(net3838),
.Y(net4020)
);

OAI21x1_ASAP7_75t_R c3990(
.A1(net3153),
.A2(net3708),
.B(net3151),
.Y(net4021)
);

AND2x6_ASAP7_75t_R c3991(
.A(net3929),
.B(net2164),
.Y(net4022)
);

BUFx4f_ASAP7_75t_R c3992(
.A(net10425),
.Y(net4023)
);

HAxp5_ASAP7_75t_R c3993(
.A(net4000),
.B(net3085),
.CON(net4024)
);

BUFx5_ASAP7_75t_R c3994(
.A(net3156),
.Y(net4025)
);

NAND2x1_ASAP7_75t_R c3995(
.A(net3920),
.B(net4017),
.Y(net4026)
);

BUFx6f_ASAP7_75t_R c3996(
.A(net4025),
.Y(net4027)
);

NAND2x1p5_ASAP7_75t_R c3997(
.A(net4015),
.B(net3846),
.Y(net4028)
);

NAND2x2_ASAP7_75t_R c3998(
.A(net3119),
.B(net1238),
.Y(net4029)
);

OAI21xp33_ASAP7_75t_R c3999(
.A1(net4020),
.A2(net3139),
.B(net4015),
.Y(net4030)
);

BUFx8_ASAP7_75t_R c4000(
.A(net3073),
.Y(net4031)
);

CKINVDCx10_ASAP7_75t_R c4001(
.A(net9745),
.Y(net4032)
);

CKINVDCx11_ASAP7_75t_R c4002(
.A(net10106),
.Y(net4033)
);

CKINVDCx12_ASAP7_75t_R c4003(
.A(net3957),
.Y(net4034)
);

CKINVDCx14_ASAP7_75t_R c4004(
.A(net2183),
.Y(net4035)
);

NAND2xp33_ASAP7_75t_R c4005(
.A(net1280),
.B(net2204),
.Y(net4036)
);

NAND2xp5_ASAP7_75t_R c4006(
.A(net3783),
.B(net3992),
.Y(net4037)
);

CKINVDCx16_ASAP7_75t_R c4007(
.A(net3868),
.Y(net4038)
);

OAI21xp5_ASAP7_75t_R c4008(
.A1(net4029),
.A2(net3170),
.B(net9709),
.Y(net4039)
);

NAND2xp67_ASAP7_75t_R c4009(
.A(net3096),
.B(net2045),
.Y(net4040)
);

NOR2x1_ASAP7_75t_R c4010(
.A(net3923),
.B(net9900),
.Y(net4041)
);

CKINVDCx20_ASAP7_75t_R c4011(
.A(net3120),
.Y(net4042)
);

CKINVDCx5p33_ASAP7_75t_R c4012(
.A(net10106),
.Y(net4043)
);

OR3x1_ASAP7_75t_R c4013(
.A(net3838),
.B(net3137),
.C(net4036),
.Y(net4044)
);

CKINVDCx6p67_ASAP7_75t_R c4014(
.A(net9864),
.Y(net4045)
);

NOR2x1p5_ASAP7_75t_R c4015(
.A(net4042),
.B(net3153),
.Y(net4046)
);

NOR2x2_ASAP7_75t_R c4016(
.A(net3933),
.B(net3150),
.Y(net4047)
);

CKINVDCx8_ASAP7_75t_R c4017(
.A(net9982),
.Y(net4048)
);

OR3x2_ASAP7_75t_R c4018(
.A(net3991),
.B(net2164),
.C(net10038),
.Y(net4049)
);

CKINVDCx9p33_ASAP7_75t_R c4019(
.A(net3137),
.Y(net4050)
);

NOR2xp33_ASAP7_75t_R c4020(
.A(net4023),
.B(net4036),
.Y(net4051)
);

HB1xp67_ASAP7_75t_R c4021(
.A(net4048),
.Y(net4052)
);

NOR2xp67_ASAP7_75t_R c4022(
.A(net2942),
.B(net10023),
.Y(net4053)
);

OR3x4_ASAP7_75t_R c4023(
.A(net3151),
.B(net4052),
.C(net3092),
.Y(net4054)
);

HB2xp67_ASAP7_75t_R c4024(
.A(net10444),
.Y(net4055)
);

OR2x2_ASAP7_75t_R c4025(
.A(net3845),
.B(net4042),
.Y(net4056)
);

OR2x4_ASAP7_75t_R c4026(
.A(net4035),
.B(net4047),
.Y(net4057)
);

HB3xp67_ASAP7_75t_R c4027(
.A(net4057),
.Y(net4058)
);

HB4xp67_ASAP7_75t_R c4028(
.A(net10096),
.Y(net4059)
);

OR2x6_ASAP7_75t_R c4029(
.A(net3135),
.B(net3132),
.Y(net4060)
);

XNOR2x1_ASAP7_75t_R c4030(
.B(net4034),
.A(net4017),
.Y(net4061)
);

XNOR2x2_ASAP7_75t_R c4031(
.A(net4053),
.B(net4056),
.Y(net4062)
);

INVx11_ASAP7_75t_R c4032(
.A(net10539),
.Y(net4063)
);

XNOR2xp5_ASAP7_75t_R c4033(
.A(net4011),
.B(net4054),
.Y(net4064)
);

XOR2x1_ASAP7_75t_R c4034(
.A(net3707),
.B(net4059),
.Y(net4065)
);

DFFASRHQNx1_ASAP7_75t_R c4035(
.D(net4028),
.RESETN(net3941),
.SETN(net4036),
.CLK(clk),
.QN(net4066)
);

XOR2x2_ASAP7_75t_R c4036(
.A(net4013),
.B(net4059),
.Y(net4067)
);

AND3x1_ASAP7_75t_R c4037(
.A(net3924),
.B(net3895),
.C(net4035),
.Y(net4068)
);

INVx13_ASAP7_75t_R c4038(
.A(net10481),
.Y(net4069)
);

XOR2xp5_ASAP7_75t_R c4039(
.A(net4050),
.B(net3939),
.Y(net4070)
);

SDFHx1_ASAP7_75t_R c4040(
.D(net4066),
.SE(net3859),
.SI(net9741),
.CLK(clk),
.QN(net4071)
);

AND3x2_ASAP7_75t_R c4041(
.A(net4029),
.B(net2235),
.C(net4066),
.Y(net4072)
);

AND2x2_ASAP7_75t_R c4042(
.A(net4060),
.B(net4061),
.Y(net4073)
);

AND2x4_ASAP7_75t_R c4043(
.A(net4052),
.B(net4064),
.Y(net4074)
);

AND2x6_ASAP7_75t_R c4044(
.A(net3867),
.B(net4054),
.Y(net4075)
);

ICGx1_ASAP7_75t_R c4045(
.ENA(net4036),
.SE(net4075),
.CLK(clk),
.GCLK(net4076)
);

AND3x4_ASAP7_75t_R c4046(
.A(net4076),
.B(net4042),
.C(net10089),
.Y(net4077)
);

INVx1_ASAP7_75t_R c4047(
.A(net10425),
.Y(net4078)
);

OA22x2_ASAP7_75t_R c4048(
.A1(net4078),
.A2(net4073),
.B1(net4055),
.B2(net4059),
.Y(net4079)
);

AO21x1_ASAP7_75t_R c4049(
.A1(net4079),
.A2(net4045),
.B(net4077),
.Y(net4080)
);

AO21x2_ASAP7_75t_R c4050(
.A1(net4022),
.A2(net4076),
.B(net10089),
.Y(net4081)
);

HAxp5_ASAP7_75t_R c4051(
.A(net3073),
.B(net10038),
.CON(net4083),
.SN(net4082)
);

NAND2x1_ASAP7_75t_R c4052(
.A(net3091),
.B(net2183),
.Y(net4084)
);

AOI21x1_ASAP7_75t_R c4053(
.A1(net3997),
.A2(net4075),
.B(net4036),
.Y(net4085)
);

NAND2x1p5_ASAP7_75t_R c4054(
.A(net3000),
.B(net4045),
.Y(net4086)
);

SDFHx2_ASAP7_75t_R c4055(
.D(net3950),
.SE(net4086),
.SI(net4076),
.CLK(clk),
.QN(net4087)
);

AOI21xp33_ASAP7_75t_R c4056(
.A1(net3139),
.A2(net4077),
.B(net4055),
.Y(net4088)
);

AOI21xp5_ASAP7_75t_R c4057(
.A1(net4074),
.A2(net4071),
.B(net4055),
.Y(net4089)
);

OA31x2_ASAP7_75t_R c4058(
.A1(net4076),
.A2(net3977),
.A3(net3951),
.B1(net9777),
.Y(net4090)
);

FAx1_ASAP7_75t_R c4059(
.A(net4089),
.B(net4059),
.CI(net4082),
.SN(net4092),
.CON(net4091)
);

MAJIxp5_ASAP7_75t_R c4060(
.A(net4069),
.B(net3003),
.C(net10240),
.Y(net4093)
);

MAJx2_ASAP7_75t_R c4061(
.A(net4087),
.B(net4092),
.C(net3951),
.Y(net4094)
);

MAJx3_ASAP7_75t_R c4062(
.A(net4070),
.B(net4061),
.C(net4091),
.Y(net4095)
);

SDFHx3_ASAP7_75t_R c4063(
.D(net4092),
.SE(net4088),
.SI(net4082),
.CLK(clk),
.QN(net4096)
);

OA33x2_ASAP7_75t_R c4064(
.A1(net4093),
.A2(net3951),
.A3(net4087),
.B1(net4086),
.B2(net4045),
.B3(net4027),
.Y(net4097)
);

NAND3x1_ASAP7_75t_R c4065(
.A(net4039),
.B(net4071),
.C(net9900),
.Y(net4098)
);

SDFHx4_ASAP7_75t_R c4066(
.D(net3951),
.SE(net4052),
.SI(net10130),
.CLK(clk),
.QN(net4099)
);

OAI222xp33_ASAP7_75t_R c4067(
.A1(net4163),
.A2(net3177),
.B1(net3234),
.B2(net4179),
.C1(net3163),
.C2(net2167),
.Y(net4100)
);

NAND2x2_ASAP7_75t_R c4068(
.A(net4161),
.B(net4179),
.Y(net4101)
);

NAND2xp33_ASAP7_75t_R c4069(
.A(net4178),
.B(net4177),
.Y(net4102)
);

NAND2xp5_ASAP7_75t_R c4070(
.A(net4156),
.B(net4136),
.Y(net4103)
);

SDFLx1_ASAP7_75t_R c4071(
.D(net4152),
.SE(net3234),
.SI(net3229),
.CLK(clk),
.QN(net4104)
);

OAI211xp5_ASAP7_75t_R c4072(
.A1(net2153),
.A2(net4177),
.B(net4138),
.C(net3941),
.Y(net4105)
);

NAND3x2_ASAP7_75t_R c4073(
.B(net4088),
.C(net4103),
.A(net4130),
.Y(net4106)
);

NAND2xp67_ASAP7_75t_R c4074(
.A(net4181),
.B(net4136),
.Y(net4107)
);

NOR2x1_ASAP7_75t_R c4075(
.A(net4175),
.B(net4146),
.Y(net4108)
);

NOR2x1p5_ASAP7_75t_R c4076(
.A(net4103),
.B(net3203),
.Y(net4109)
);

NAND3xp33_ASAP7_75t_R c4077(
.A(net4183),
.B(net4109),
.C(net4108),
.Y(net4110)
);

NOR3x1_ASAP7_75t_R c4078(
.A(net4174),
.B(net4067),
.C(net10084),
.Y(net4111)
);

NOR2x2_ASAP7_75t_R c4079(
.A(net4160),
.B(net4031),
.Y(net4112)
);

NOR2xp33_ASAP7_75t_R c4080(
.A(net4133),
.B(net4073),
.Y(net4113)
);

NOR2xp67_ASAP7_75t_R c4081(
.A(net4105),
.B(net4179),
.Y(net4114)
);

OR2x2_ASAP7_75t_R c4082(
.A(net4102),
.B(net4175),
.Y(net4115)
);

OR2x4_ASAP7_75t_R c4083(
.A(net4146),
.B(net4109),
.Y(net4116)
);

INVx2_ASAP7_75t_R c4084(
.A(net4130),
.Y(net4117)
);

ICGx2_ASAP7_75t_R c4085(
.ENA(net4114),
.SE(net3218),
.CLK(clk),
.GCLK(net4118)
);

NOR3x2_ASAP7_75t_R c4086(
.B(net3229),
.C(net4105),
.A(net4081),
.Y(net4119)
);

NOR3xp33_ASAP7_75t_R c4087(
.A(net4118),
.B(net4130),
.C(net4171),
.Y(net4120)
);

OA21x2_ASAP7_75t_R c4088(
.A1(net4164),
.A2(net4154),
.B(net4116),
.Y(net4121)
);

INVx3_ASAP7_75t_R c4089(
.A(net4144),
.Y(net4122)
);

OR2x6_ASAP7_75t_R c4090(
.A(net4111),
.B(net3155),
.Y(net4123)
);

OAI321xp33_ASAP7_75t_R c4091(
.A1(net4068),
.A2(net4104),
.A3(net3228),
.B1(net4077),
.B2(net4054),
.C(net3246),
.Y(net4124)
);

OAI21x1_ASAP7_75t_R c4092(
.A1(net2265),
.A2(net4118),
.B(net4123),
.Y(net4125)
);

OAI21xp33_ASAP7_75t_R c4093(
.A1(net4120),
.A2(net4145),
.B(net10084),
.Y(net4126)
);

OAI21xp5_ASAP7_75t_R c4094(
.A1(net4115),
.A2(net4120),
.B(net4124),
.Y(net4127)
);

OR3x1_ASAP7_75t_R c4095(
.A(net4115),
.B(net4040),
.C(net10073),
.Y(net4128)
);

XNOR2x1_ASAP7_75t_R c4096(
.B(net4109),
.A(net10073),
.Y(net4129)
);

SDFLx2_ASAP7_75t_R c4097(
.D(net3817),
.SE(net3245),
.SI(net9709),
.CLK(clk),
.QN(net4130)
);

XNOR2x2_ASAP7_75t_R c4098(
.A(net1833),
.B(net4077),
.Y(net4131)
);

XNOR2xp5_ASAP7_75t_R c4099(
.A(net3895),
.B(net4054),
.Y(net4132)
);

INVx4_ASAP7_75t_R c4100(
.A(net4132),
.Y(net4133)
);

INVx5_ASAP7_75t_R c4101(
.A(net9933),
.Y(net4134)
);

INVx6_ASAP7_75t_R c4102(
.A(net2167),
.Y(net4135)
);

INVx8_ASAP7_75t_R c4103(
.A(net9136),
.Y(net4136)
);

INVxp33_ASAP7_75t_R c4104(
.A(net9136),
.Y(net4137)
);

INVxp67_ASAP7_75t_R c4105(
.A(net10132),
.Y(net4138)
);

XOR2x1_ASAP7_75t_R c4106(
.A(net3204),
.B(net1196),
.Y(net4139)
);

BUFx10_ASAP7_75t_R c4107(
.A(net3245),
.Y(net4140)
);

BUFx12_ASAP7_75t_R c4108(
.A(net9218),
.Y(net4141)
);

BUFx12f_ASAP7_75t_R c4109(
.A(net9966),
.Y(net4142)
);

XOR2x2_ASAP7_75t_R c4110(
.A(net4041),
.B(net4054),
.Y(net4143)
);

BUFx16f_ASAP7_75t_R c4111(
.A(net4067),
.Y(net4144)
);

XOR2xp5_ASAP7_75t_R c4112(
.A(net3211),
.B(net3227),
.Y(net4145)
);

AND2x2_ASAP7_75t_R c4113(
.A(net4096),
.B(net1348),
.Y(net4146)
);

AND2x4_ASAP7_75t_R c4114(
.A(net3254),
.B(net4134),
.Y(net4147)
);

OR3x2_ASAP7_75t_R c4115(
.A(net3157),
.B(net4066),
.C(net3772),
.Y(net4148)
);

AND2x6_ASAP7_75t_R c4116(
.A(net4145),
.B(net4096),
.Y(net4149)
);

BUFx24_ASAP7_75t_R c4117(
.A(net3177),
.Y(net4150)
);

HAxp5_ASAP7_75t_R c4118(
.A(net4063),
.B(net4027),
.CON(net4152),
.SN(net4151)
);

BUFx2_ASAP7_75t_R c4119(
.A(net2264),
.Y(net4153)
);

ICGx2p67DC_ASAP7_75t_R c4120(
.ENA(net4152),
.SE(net4080),
.CLK(clk),
.GCLK(net4154)
);

OR3x4_ASAP7_75t_R c4121(
.A(net350),
.B(net4144),
.C(net3872),
.Y(net4155)
);

NAND2x1_ASAP7_75t_R c4122(
.A(net4154),
.B(net3941),
.Y(net4156)
);

AND3x1_ASAP7_75t_R c4123(
.A(net4084),
.B(net4151),
.C(net3254),
.Y(net4157)
);

AND3x2_ASAP7_75t_R c4124(
.A(net3155),
.B(net4061),
.C(net2264),
.Y(net4158)
);

NAND2x1p5_ASAP7_75t_R c4125(
.A(net4144),
.B(net2264),
.Y(net4159)
);

BUFx3_ASAP7_75t_R c4126(
.A(net10504),
.Y(net4160)
);

OAI22x1_ASAP7_75t_R c4127(
.A1(net4142),
.A2(net3254),
.B1(net4158),
.B2(net2214),
.Y(net4161)
);

NAND2x2_ASAP7_75t_R c4128(
.A(net4135),
.B(net3157),
.Y(net4162)
);

NAND2xp33_ASAP7_75t_R c4129(
.A(net4161),
.B(net2292),
.Y(net4163)
);

NAND2xp5_ASAP7_75t_R c4130(
.A(net4061),
.B(net4096),
.Y(net4164)
);

BUFx4_ASAP7_75t_R c4131(
.A(net4159),
.Y(net4165)
);

BUFx4f_ASAP7_75t_R c4132(
.A(net4136),
.Y(net4166)
);

NAND2xp67_ASAP7_75t_R c4133(
.A(net3772),
.B(net3211),
.Y(net4167)
);

NOR2x1_ASAP7_75t_R c4134(
.A(net4066),
.B(net4153),
.Y(net4168)
);

NOR2x1p5_ASAP7_75t_R c4135(
.A(net4159),
.B(net4150),
.Y(net4169)
);

BUFx5_ASAP7_75t_R c4136(
.A(net10552),
.Y(net4170)
);

NOR2x2_ASAP7_75t_R c4137(
.A(net4156),
.B(net10195),
.Y(net4171)
);

BUFx6f_ASAP7_75t_R c4138(
.A(net10071),
.Y(net4172)
);

BUFx8_ASAP7_75t_R c4139(
.A(net9967),
.Y(net4173)
);

SDFLx3_ASAP7_75t_R c4140(
.D(net4131),
.SE(net3176),
.SI(net2214),
.CLK(clk),
.QN(net4174)
);

CKINVDCx10_ASAP7_75t_R c4141(
.A(net3203),
.Y(net4175)
);

CKINVDCx11_ASAP7_75t_R c4142(
.A(net10395),
.Y(net4176)
);

SDFLx4_ASAP7_75t_R c4143(
.D(net1371),
.SE(net4169),
.SI(net3192),
.CLK(clk),
.QN(net4177)
);

NOR2xp33_ASAP7_75t_R c4144(
.A(net4054),
.B(net4143),
.Y(net4178)
);

NOR2xp67_ASAP7_75t_R c4145(
.A(net4169),
.B(net9868),
.Y(net4179)
);

OR2x2_ASAP7_75t_R c4146(
.A(net3186),
.B(net2214),
.Y(net4180)
);

OR2x4_ASAP7_75t_R c4147(
.A(net4143),
.B(net3086),
.Y(net4181)
);

OR2x6_ASAP7_75t_R c4148(
.A(net4172),
.B(net446),
.Y(net4182)
);

CKINVDCx12_ASAP7_75t_R c4149(
.A(net10517),
.Y(net4183)
);

CKINVDCx14_ASAP7_75t_R c4150(
.A(net10491),
.Y(net4184)
);

AND3x4_ASAP7_75t_R c4151(
.A(net3878),
.B(net3228),
.C(net9813),
.Y(net4185)
);

CKINVDCx16_ASAP7_75t_R c4152(
.A(net10017),
.Y(net4186)
);

XNOR2x1_ASAP7_75t_R c4153(
.B(net3329),
.A(net3339),
.Y(net4187)
);

XNOR2x2_ASAP7_75t_R c4154(
.A(net3275),
.B(net4182),
.Y(net4188)
);

CKINVDCx20_ASAP7_75t_R c4155(
.A(net4083),
.Y(net4189)
);

XNOR2xp5_ASAP7_75t_R c4156(
.A(net3318),
.B(net4169),
.Y(net4190)
);

XOR2x1_ASAP7_75t_R c4157(
.A(net4108),
.B(net4095),
.Y(net4191)
);

CKINVDCx5p33_ASAP7_75t_R c4158(
.A(net4153),
.Y(net4192)
);

XOR2x2_ASAP7_75t_R c4159(
.A(net3235),
.B(net4107),
.Y(net4193)
);

CKINVDCx6p67_ASAP7_75t_R c4160(
.A(net4077),
.Y(net4194)
);

CKINVDCx8_ASAP7_75t_R c4161(
.A(net4123),
.Y(net4195)
);

AO21x1_ASAP7_75t_R c4162(
.A1(net4186),
.A2(net3339),
.B(net4166),
.Y(net4196)
);

XOR2xp5_ASAP7_75t_R c4163(
.A(net3340),
.B(net3218),
.Y(net4197)
);

CKINVDCx9p33_ASAP7_75t_R c4164(
.A(net10038),
.Y(net4198)
);

AO21x2_ASAP7_75t_R c4165(
.A1(net4197),
.A2(net4124),
.B(net4083),
.Y(net4199)
);

AOI21x1_ASAP7_75t_R c4166(
.A1(net3280),
.A2(net4165),
.B(net1446),
.Y(net4200)
);

AND2x2_ASAP7_75t_R c4167(
.A(net3277),
.B(net2399),
.Y(net4201)
);

AND2x4_ASAP7_75t_R c4168(
.A(net4196),
.B(net4134),
.Y(net4202)
);

AND2x6_ASAP7_75t_R c4169(
.A(net4191),
.B(net2345),
.Y(net4203)
);

HAxp5_ASAP7_75t_R c4170(
.A(net4165),
.B(net4197),
.CON(net4204)
);

HB1xp67_ASAP7_75t_R c4171(
.A(net445),
.Y(net4205)
);

HB2xp67_ASAP7_75t_R c4172(
.A(net10512),
.Y(net4206)
);

NAND2x1_ASAP7_75t_R c4173(
.A(net4107),
.B(net4198),
.Y(net4207)
);

NAND2x1p5_ASAP7_75t_R c4174(
.A(net4169),
.B(net4170),
.Y(net4208)
);

HB3xp67_ASAP7_75t_R c4175(
.A(net3274),
.Y(net4209)
);

HB4xp67_ASAP7_75t_R c4176(
.A(net4141),
.Y(net4210)
);

INVx11_ASAP7_75t_R c4177(
.A(net10510),
.Y(net4211)
);

INVx13_ASAP7_75t_R c4178(
.A(net4201),
.Y(net4212)
);

INVx1_ASAP7_75t_R c4179(
.A(net10390),
.Y(net4213)
);

INVx2_ASAP7_75t_R c4180(
.A(net4129),
.Y(net4214)
);

NAND2x2_ASAP7_75t_R c4181(
.A(net4211),
.B(net4027),
.Y(net4215)
);

NAND2xp33_ASAP7_75t_R c4182(
.A(net3228),
.B(net4027),
.Y(net4216)
);

NAND2xp5_ASAP7_75t_R c4183(
.A(net4208),
.B(net4214),
.Y(net4217)
);

INVx3_ASAP7_75t_R c4184(
.A(net4205),
.Y(net4218)
);

AOI21xp33_ASAP7_75t_R c4185(
.A1(net2359),
.A2(net1462),
.B(net4214),
.Y(net4219)
);

NAND2xp67_ASAP7_75t_R c4186(
.A(net4189),
.B(net4195),
.Y(net4220)
);

DFFASRHQNx1_ASAP7_75t_R c4187(
.D(net3296),
.RESETN(net4197),
.SETN(net353),
.CLK(clk),
.QN(net4221)
);

INVx4_ASAP7_75t_R c4188(
.A(net4190),
.Y(net4222)
);

NOR2x1_ASAP7_75t_R c4189(
.A(net2413),
.B(net3339),
.Y(net4223)
);

AOI21xp5_ASAP7_75t_R c4190(
.A1(net3231),
.A2(net4153),
.B(net3269),
.Y(net4224)
);

FAx1_ASAP7_75t_R c4191(
.A(net4220),
.B(net3297),
.CI(net3280),
.SN(net4226),
.CON(net4225)
);

SDFHx1_ASAP7_75t_R c4192(
.D(net2253),
.SE(net4203),
.SI(net4188),
.CLK(clk),
.QN(net4227)
);

NOR2x1p5_ASAP7_75t_R c4193(
.A(net4221),
.B(net4108),
.Y(net4228)
);

NOR2x2_ASAP7_75t_R c4194(
.A(net4224),
.B(net4222),
.Y(net4229)
);

NOR2xp33_ASAP7_75t_R c4195(
.A(net4225),
.B(net10156),
.Y(net4230)
);

MAJIxp5_ASAP7_75t_R c4196(
.A(net4205),
.B(net4225),
.C(net9899),
.Y(net4231)
);

INVx5_ASAP7_75t_R c4197(
.A(net10549),
.Y(net4232)
);

INVx6_ASAP7_75t_R c4198(
.A(net10361),
.Y(net4233)
);

INVx8_ASAP7_75t_R c4199(
.A(net4226),
.Y(net4234)
);

MAJx2_ASAP7_75t_R c4200(
.A(net4216),
.B(net4206),
.C(net4083),
.Y(net4235)
);

NOR2xp67_ASAP7_75t_R c4201(
.A(net4227),
.B(net4213),
.Y(net4236)
);

OR2x2_ASAP7_75t_R c4202(
.A(net3327),
.B(net10161),
.Y(net4237)
);

INVxp33_ASAP7_75t_R c4203(
.A(net10445),
.Y(net4238)
);

MAJx3_ASAP7_75t_R c4204(
.A(net4212),
.B(net4002),
.C(net4081),
.Y(net4239)
);

NAND3x1_ASAP7_75t_R c4205(
.A(net4237),
.B(net4226),
.C(net4221),
.Y(net4240)
);

OR2x4_ASAP7_75t_R c4206(
.A(net4238),
.B(net4220),
.Y(net4241)
);

NAND3x2_ASAP7_75t_R c4207(
.B(net4119),
.C(net4184),
.A(net3235),
.Y(net4242)
);

OR2x6_ASAP7_75t_R c4208(
.A(net4239),
.B(net4198),
.Y(net4243)
);

XNOR2x1_ASAP7_75t_R c4209(
.B(net4192),
.A(net4226),
.Y(net4244)
);

SDFHx2_ASAP7_75t_R c4210(
.D(net3092),
.SE(net4238),
.SI(net2393),
.CLK(clk),
.QN(net4245)
);

XNOR2x2_ASAP7_75t_R c4211(
.A(net4215),
.B(net4227),
.Y(net4246)
);

XNOR2xp5_ASAP7_75t_R c4212(
.A(net4222),
.B(net10067),
.Y(net4247)
);

INVxp67_ASAP7_75t_R c4213(
.A(net10157),
.Y(net4248)
);

BUFx10_ASAP7_75t_R c4214(
.A(net10017),
.Y(net4249)
);

AO32x1_ASAP7_75t_R c4215(
.A1(net1355),
.A2(net4227),
.A3(net4246),
.B1(net3092),
.B2(net2337),
.Y(net4250)
);

SDFHx3_ASAP7_75t_R c4216(
.D(net4184),
.SE(net3163),
.SI(net2235),
.CLK(clk),
.QN(net4251)
);

XOR2x1_ASAP7_75t_R c4217(
.A(net4232),
.B(net4233),
.Y(net4252)
);

NAND3xp33_ASAP7_75t_R c4218(
.A(net4233),
.B(net4220),
.C(net4252),
.Y(net4253)
);

NOR3x1_ASAP7_75t_R c4219(
.A(net4194),
.B(net4243),
.C(net4241),
.Y(net4254)
);

XOR2x2_ASAP7_75t_R c4220(
.A(net4193),
.B(net4243),
.Y(net4255)
);

XOR2xp5_ASAP7_75t_R c4221(
.A(net4240),
.B(net4255),
.Y(net4256)
);

NOR3x2_ASAP7_75t_R c4222(
.B(net4248),
.C(net4221),
.A(net4223),
.Y(net4257)
);

NOR3xp33_ASAP7_75t_R c4223(
.A(net3297),
.B(net4238),
.C(net4245),
.Y(net4258)
);

AND2x2_ASAP7_75t_R c4224(
.A(net4253),
.B(net4258),
.Y(net4259)
);

OA21x2_ASAP7_75t_R c4225(
.A1(net4213),
.A2(net4259),
.B(net3092),
.Y(net4260)
);

OAI21x1_ASAP7_75t_R c4226(
.A1(net4244),
.A2(net4255),
.B(net10103),
.Y(net4261)
);

AND2x4_ASAP7_75t_R c4227(
.A(net4259),
.B(net4244),
.Y(net4262)
);

OAI21xp33_ASAP7_75t_R c4228(
.A1(net4245),
.A2(net4262),
.B(net4257),
.Y(net4263)
);

AND2x6_ASAP7_75t_R c4229(
.A(net4205),
.B(net10165),
.Y(net4264)
);

OAI21xp5_ASAP7_75t_R c4230(
.A1(net4263),
.A2(net4259),
.B(net4252),
.Y(net4265)
);

SDFHx4_ASAP7_75t_R c4231(
.D(net4086),
.SE(net4258),
.SI(net4260),
.CLK(clk),
.QN(net4266)
);

OR3x1_ASAP7_75t_R c4232(
.A(net4261),
.B(net4266),
.C(net4264),
.Y(net4267)
);

OR3x2_ASAP7_75t_R c4233(
.A(net4260),
.B(net4095),
.C(net1446),
.Y(net4268)
);

BUFx12_ASAP7_75t_R c4234(
.A(net4241),
.Y(net4269)
);

OR3x4_ASAP7_75t_R c4235(
.A(net4073),
.B(net3366),
.C(net3421),
.Y(net4270)
);

BUFx12f_ASAP7_75t_R c4236(
.A(net3409),
.Y(net4271)
);

BUFx16f_ASAP7_75t_R c4237(
.A(net3327),
.Y(net4272)
);

HAxp5_ASAP7_75t_R c4238(
.A(net4228),
.B(net10241),
.CON(net4274),
.SN(net4273)
);

NAND2x1_ASAP7_75t_R c4239(
.A(net4258),
.B(net4256),
.Y(net4275)
);

NAND2x1p5_ASAP7_75t_R c4240(
.A(net3366),
.B(net10226),
.Y(net4276)
);

AND3x1_ASAP7_75t_R c4241(
.A(net2421),
.B(net4229),
.C(net624),
.Y(net4277)
);

NAND2x2_ASAP7_75t_R c4242(
.A(net3418),
.B(net4241),
.Y(net4278)
);

BUFx24_ASAP7_75t_R c4243(
.A(net4278),
.Y(net4279)
);

AND3x2_ASAP7_75t_R c4244(
.A(net624),
.B(net3418),
.C(net2499),
.Y(net4280)
);

NAND2xp33_ASAP7_75t_R c4245(
.A(net3278),
.B(net3366),
.Y(net4281)
);

BUFx2_ASAP7_75t_R c4246(
.A(net10150),
.Y(net4282)
);

NAND2xp5_ASAP7_75t_R c4247(
.A(net2259),
.B(net4200),
.Y(net4283)
);

AO32x2_ASAP7_75t_R c4248(
.A1(net4230),
.A2(net3362),
.A3(net2498),
.B1(net3412),
.B2(net10241),
.Y(net4284)
);

NAND2xp67_ASAP7_75t_R c4249(
.A(net561),
.B(net4158),
.Y(net4285)
);

NOR2x1_ASAP7_75t_R c4250(
.A(net2404),
.B(net4260),
.Y(net4286)
);

NOR2x1p5_ASAP7_75t_R c4251(
.A(net4200),
.B(net3373),
.Y(net4287)
);

BUFx3_ASAP7_75t_R c4252(
.A(net3291),
.Y(net4288)
);

NOR2x2_ASAP7_75t_R c4253(
.A(net3163),
.B(net4200),
.Y(net4289)
);

BUFx4_ASAP7_75t_R c4254(
.A(net3385),
.Y(net4290)
);

NOR2xp33_ASAP7_75t_R c4255(
.A(net1446),
.B(net10241),
.Y(net4291)
);

AOI221x1_ASAP7_75t_R c4256(
.A1(net4271),
.A2(net4268),
.B1(net3327),
.B2(net3163),
.C(net3412),
.Y(net4292)
);

NOR2xp67_ASAP7_75t_R c4257(
.A(net4282),
.B(net3416),
.Y(net4293)
);

OR2x2_ASAP7_75t_R c4258(
.A(net2437),
.B(net3412),
.Y(net4294)
);

OAI22xp33_ASAP7_75t_R c4259(
.A1(net1571),
.A2(net3403),
.B1(net3214),
.B2(net2463),
.Y(net4295)
);

BUFx4f_ASAP7_75t_R c4260(
.A(net4276),
.Y(net4296)
);

OR2x4_ASAP7_75t_R c4261(
.A(net4279),
.B(net4269),
.Y(net4297)
);

BUFx5_ASAP7_75t_R c4262(
.A(net10478),
.Y(net4298)
);

BUFx6f_ASAP7_75t_R c4263(
.A(net4255),
.Y(net4299)
);

BUFx8_ASAP7_75t_R c4264(
.A(net4150),
.Y(net4300)
);

OR2x6_ASAP7_75t_R c4265(
.A(net4235),
.B(net4274),
.Y(net4301)
);

XNOR2x1_ASAP7_75t_R c4266(
.B(net4285),
.A(net4081),
.Y(net4302)
);

CKINVDCx10_ASAP7_75t_R c4267(
.A(net10213),
.Y(net4303)
);

CKINVDCx11_ASAP7_75t_R c4268(
.A(net10470),
.Y(net4304)
);

XNOR2x2_ASAP7_75t_R c4269(
.A(net4304),
.B(net10113),
.Y(net4305)
);

XNOR2xp5_ASAP7_75t_R c4270(
.A(net4297),
.B(net3385),
.Y(net4306)
);

CKINVDCx12_ASAP7_75t_R c4271(
.A(net10518),
.Y(net4307)
);

XOR2x1_ASAP7_75t_R c4272(
.A(net4223),
.B(net4252),
.Y(net4308)
);

XOR2x2_ASAP7_75t_R c4273(
.A(net4291),
.B(net4308),
.Y(net4309)
);

XOR2xp5_ASAP7_75t_R c4274(
.A(net3362),
.B(net4308),
.Y(net4310)
);

AND2x2_ASAP7_75t_R c4275(
.A(net3345),
.B(net4297),
.Y(net4311)
);

AND2x4_ASAP7_75t_R c4276(
.A(net4303),
.B(net4294),
.Y(net4312)
);

AND2x6_ASAP7_75t_R c4277(
.A(net4269),
.B(net325),
.Y(net4313)
);

CKINVDCx14_ASAP7_75t_R c4278(
.A(net4280),
.Y(net4314)
);

CKINVDCx16_ASAP7_75t_R c4279(
.A(net4304),
.Y(net4315)
);

OAI22xp5_ASAP7_75t_R c4280(
.A1(net4306),
.A2(net272),
.B1(net4269),
.B2(net3412),
.Y(net4316)
);

CKINVDCx20_ASAP7_75t_R c4281(
.A(net4296),
.Y(net4317)
);

CKINVDCx5p33_ASAP7_75t_R c4282(
.A(net10137),
.Y(net4318)
);

HAxp5_ASAP7_75t_R c4283(
.A(net4290),
.B(net10113),
.CON(net4319)
);

NAND2x1_ASAP7_75t_R c4284(
.A(net4319),
.B(net2262),
.Y(net4320)
);

CKINVDCx6p67_ASAP7_75t_R c4285(
.A(net9985),
.Y(net4321)
);

AND3x4_ASAP7_75t_R c4286(
.A(net4274),
.B(net4236),
.C(net4223),
.Y(net4322)
);

CKINVDCx8_ASAP7_75t_R c4287(
.A(net4300),
.Y(net4323)
);

NAND2x1p5_ASAP7_75t_R c4288(
.A(net1462),
.B(net4297),
.Y(net4324)
);

CKINVDCx9p33_ASAP7_75t_R c4289(
.A(net4299),
.Y(net4325)
);

HB1xp67_ASAP7_75t_R c4290(
.A(net10076),
.Y(net4326)
);

OAI31xp33_ASAP7_75t_R c4291(
.A1(net4266),
.A2(net4309),
.A3(net4324),
.B(net10156),
.Y(net4327)
);

HB2xp67_ASAP7_75t_R c4292(
.A(net10045),
.Y(net4328)
);

NAND2x2_ASAP7_75t_R c4293(
.A(net4326),
.B(net4214),
.Y(net4329)
);

NAND2xp33_ASAP7_75t_R c4294(
.A(net4314),
.B(net3941),
.Y(net4330)
);

AOI221xp5_ASAP7_75t_R c4295(
.A1(net4320),
.A2(net3163),
.B1(net4328),
.B2(net3404),
.C(net3412),
.Y(net4331)
);

NAND2xp5_ASAP7_75t_R c4296(
.A(net4273),
.B(net9735),
.Y(net4332)
);

OAI31xp67_ASAP7_75t_R c4297(
.A1(net4318),
.A2(net3409),
.A3(net4256),
.B(net3272),
.Y(net4333)
);

AO21x1_ASAP7_75t_R c4298(
.A1(net4323),
.A2(net3419),
.B(net3239),
.Y(net4334)
);

HB3xp67_ASAP7_75t_R c4299(
.A(net10478),
.Y(net4335)
);

HB4xp67_ASAP7_75t_R c4300(
.A(net10535),
.Y(net4336)
);

INVx11_ASAP7_75t_R c4301(
.A(net10150),
.Y(net4337)
);

OR4x1_ASAP7_75t_R c4302(
.A(net4277),
.B(net4325),
.C(net4328),
.D(net4307),
.Y(net4338)
);

NAND2xp67_ASAP7_75t_R c4303(
.A(net9855),
.B(net10243),
.Y(net4339)
);

INVx13_ASAP7_75t_R c4304(
.A(net10137),
.Y(net4340)
);

AO21x2_ASAP7_75t_R c4305(
.A1(net4284),
.A2(net4340),
.B(net3163),
.Y(net4341)
);

OR4x2_ASAP7_75t_R c4306(
.A(net4341),
.B(net4307),
.C(net4294),
.D(net10242),
.Y(net4342)
);

INVx1_ASAP7_75t_R c4307(
.A(net10528),
.Y(net4343)
);

AOI21x1_ASAP7_75t_R c4308(
.A1(net4343),
.A2(net4340),
.B(net10243),
.Y(net4344)
);

NOR2x1_ASAP7_75t_R c4309(
.A(net4313),
.B(net10100),
.Y(net4345)
);

AOI311xp33_ASAP7_75t_R c4310(
.A1(net4328),
.A2(net4332),
.A3(net4304),
.B(net4047),
.C(net4310),
.Y(net4346)
);

NOR2x1p5_ASAP7_75t_R c4311(
.A(net4340),
.B(net9945),
.Y(net4347)
);

INVx2_ASAP7_75t_R c4312(
.A(net10461),
.Y(net4348)
);

NOR2x2_ASAP7_75t_R c4313(
.A(net4345),
.B(net4347),
.Y(net4349)
);

A2O1A1Ixp33_ASAP7_75t_R c4314(
.A1(net4348),
.A2(net4347),
.B(net4332),
.C(net4309),
.Y(net4350)
);

NOR2xp33_ASAP7_75t_R c4315(
.A(net4328),
.B(net10124),
.Y(net4351)
);

ICGx3_ASAP7_75t_R c4316(
.ENA(net1650),
.SE(net10228),
.CLK(clk),
.GCLK(net4352)
);

NOR2xp67_ASAP7_75t_R c4317(
.A(net4234),
.B(net4294),
.Y(net4353)
);

AOI21xp33_ASAP7_75t_R c4318(
.A1(net3475),
.A2(net624),
.B(net4294),
.Y(net4354)
);

INVx3_ASAP7_75t_R c4319(
.A(net2963),
.Y(net4355)
);

INVx4_ASAP7_75t_R c4320(
.A(net9137),
.Y(net4356)
);

INVx5_ASAP7_75t_R c4321(
.A(net10172),
.Y(net4357)
);

INVx6_ASAP7_75t_R c4322(
.A(net4335),
.Y(net4358)
);

AOI21xp5_ASAP7_75t_R c4323(
.A1(net3496),
.A2(net4355),
.B(net4289),
.Y(net4359)
);

INVx8_ASAP7_75t_R c4324(
.A(net4346),
.Y(net4360)
);

INVxp33_ASAP7_75t_R c4325(
.A(net2549),
.Y(net4361)
);

INVxp67_ASAP7_75t_R c4326(
.A(net10162),
.Y(net4362)
);

BUFx10_ASAP7_75t_R c4327(
.A(net9231),
.Y(net4363)
);

BUFx12_ASAP7_75t_R c4328(
.A(net3467),
.Y(net4364)
);

OR2x2_ASAP7_75t_R c4329(
.A(net4363),
.B(net9696),
.Y(net4365)
);

OR2x4_ASAP7_75t_R c4330(
.A(net4352),
.B(net4353),
.Y(net4366)
);

BUFx12f_ASAP7_75t_R c4331(
.A(net9231),
.Y(net4367)
);

BUFx16f_ASAP7_75t_R c4332(
.A(net10241),
.Y(net4368)
);

BUFx24_ASAP7_75t_R c4333(
.A(net9230),
.Y(net4369)
);

BUFx2_ASAP7_75t_R c4334(
.A(net4364),
.Y(net4370)
);

BUFx3_ASAP7_75t_R c4335(
.A(net9230),
.Y(net4371)
);

BUFx4_ASAP7_75t_R c4336(
.A(net3403),
.Y(net4372)
);

BUFx4f_ASAP7_75t_R c4337(
.A(net9223),
.Y(net4373)
);

BUFx5_ASAP7_75t_R c4338(
.A(net10152),
.Y(net4374)
);

BUFx6f_ASAP7_75t_R c4339(
.A(net4361),
.Y(net4375)
);

AND4x1_ASAP7_75t_R c4340(
.A(net3452),
.B(net4236),
.C(net4291),
.D(net4363),
.Y(net4376)
);

OR2x6_ASAP7_75t_R c4341(
.A(net1651),
.B(net4335),
.Y(net4377)
);

BUFx8_ASAP7_75t_R c4342(
.A(net4256),
.Y(net4378)
);

CKINVDCx10_ASAP7_75t_R c4343(
.A(net2529),
.Y(net4379)
);

CKINVDCx11_ASAP7_75t_R c4344(
.A(net4266),
.Y(net4380)
);

XNOR2x1_ASAP7_75t_R c4345(
.B(net3477),
.A(net3450),
.Y(net4381)
);

CKINVDCx12_ASAP7_75t_R c4346(
.A(net9195),
.Y(net4382)
);

XNOR2x2_ASAP7_75t_R c4347(
.A(net4363),
.B(net9795),
.Y(net4383)
);

CKINVDCx14_ASAP7_75t_R c4348(
.A(net4095),
.Y(net4384)
);

FAx1_ASAP7_75t_R c4349(
.A(net4365),
.B(net4307),
.CI(net4291),
.SN(net4386),
.CON(net4385)
);

MAJIxp5_ASAP7_75t_R c4350(
.A(net662),
.B(net4373),
.C(net4268),
.Y(net4387)
);

MAJx2_ASAP7_75t_R c4351(
.A(net4374),
.B(net3450),
.C(net4384),
.Y(net4388)
);

CKINVDCx16_ASAP7_75t_R c4352(
.A(net9195),
.Y(net4389)
);

XNOR2xp5_ASAP7_75t_R c4353(
.A(net4294),
.B(net4355),
.Y(net4390)
);

CKINVDCx20_ASAP7_75t_R c4354(
.A(net3455),
.Y(net4391)
);

CKINVDCx5p33_ASAP7_75t_R c4355(
.A(net10554),
.Y(net4392)
);

CKINVDCx6p67_ASAP7_75t_R c4356(
.A(net10381),
.Y(net4393)
);

CKINVDCx8_ASAP7_75t_R c4357(
.A(net10107),
.Y(net4394)
);

XOR2x1_ASAP7_75t_R c4358(
.A(net2566),
.B(net4386),
.Y(net4395)
);

XOR2x2_ASAP7_75t_R c4359(
.A(net4291),
.B(net4210),
.Y(net4396)
);

CKINVDCx9p33_ASAP7_75t_R c4360(
.A(net4337),
.Y(net4397)
);

XOR2xp5_ASAP7_75t_R c4361(
.A(net2262),
.B(net9910),
.Y(net4398)
);

AND2x2_ASAP7_75t_R c4362(
.A(net693),
.B(net2537),
.Y(net4399)
);

AND2x4_ASAP7_75t_R c4363(
.A(net4101),
.B(net4399),
.Y(net4400)
);

HB1xp67_ASAP7_75t_R c4364(
.A(net4398),
.Y(net4401)
);

AND2x6_ASAP7_75t_R c4365(
.A(net4358),
.B(net4367),
.Y(net4402)
);

HB2xp67_ASAP7_75t_R c4366(
.A(net9941),
.Y(net4403)
);

HB3xp67_ASAP7_75t_R c4367(
.A(net10388),
.Y(net4404)
);

HB4xp67_ASAP7_75t_R c4368(
.A(net9898),
.Y(net4405)
);

INVx11_ASAP7_75t_R c4369(
.A(net9869),
.Y(net4406)
);

INVx13_ASAP7_75t_R c4370(
.A(net4400),
.Y(net4407)
);

INVx1_ASAP7_75t_R c4371(
.A(net4384),
.Y(net4408)
);

INVx2_ASAP7_75t_R c4372(
.A(net4081),
.Y(net4409)
);

HAxp5_ASAP7_75t_R c4373(
.A(net4391),
.B(net4364),
.CON(net4411),
.SN(net4410)
);

NAND2x1_ASAP7_75t_R c4374(
.A(net3373),
.B(net3477),
.Y(net4412)
);

INVx3_ASAP7_75t_R c4375(
.A(net9137),
.Y(net4413)
);

INVx4_ASAP7_75t_R c4376(
.A(net4397),
.Y(net4414)
);

AOI32xp33_ASAP7_75t_R c4377(
.A1(net4405),
.A2(net2584),
.A3(net4403),
.B1(net4353),
.B2(net4264),
.Y(net4415)
);

NAND2x1p5_ASAP7_75t_R c4378(
.A(net4371),
.B(net10228),
.Y(net4416)
);

MAJx3_ASAP7_75t_R c4379(
.A(net4372),
.B(net4404),
.C(net2463),
.Y(net4417)
);

NAND2x2_ASAP7_75t_R c4380(
.A(net4383),
.B(net4257),
.Y(net4418)
);

INVx5_ASAP7_75t_R c4381(
.A(net4412),
.Y(net4419)
);

OAI33xp33_ASAP7_75t_R c4382(
.A1(net4418),
.A2(net4110),
.A3(net4386),
.B1(net4294),
.B2(net4357),
.B3(net10228),
.Y(net4420)
);

NAND3x1_ASAP7_75t_R c4383(
.A(net4390),
.B(net4416),
.C(net4406),
.Y(net4421)
);

NAND3x2_ASAP7_75t_R c4384(
.B(net4382),
.C(net4405),
.A(net9805),
.Y(net4422)
);

INVx6_ASAP7_75t_R c4385(
.A(net10022),
.Y(net4423)
);

INVx8_ASAP7_75t_R c4386(
.A(net10133),
.Y(net4424)
);

NAND2xp33_ASAP7_75t_R c4387(
.A(net4382),
.B(net4409),
.Y(net4425)
);

INVxp33_ASAP7_75t_R c4388(
.A(net10172),
.Y(net4426)
);

NAND2xp5_ASAP7_75t_R c4389(
.A(net4414),
.B(net4425),
.Y(net4427)
);

NAND2xp67_ASAP7_75t_R c4390(
.A(net4367),
.B(net4409),
.Y(net4428)
);

NAND3xp33_ASAP7_75t_R c4391(
.A(net4411),
.B(net4352),
.C(net10153),
.Y(net4429)
);

NOR2x1_ASAP7_75t_R c4392(
.A(net4396),
.B(net10044),
.Y(net4430)
);

NOR3x1_ASAP7_75t_R c4393(
.A(net1250),
.B(net4391),
.C(net10044),
.Y(net4431)
);

NAND5xp2_ASAP7_75t_R c4394(
.A(net4370),
.B(net4095),
.C(net4335),
.D(net4373),
.E(net3432),
.Y(net4432)
);

NOR5xp2_ASAP7_75t_R c4395(
.A(net2537),
.B(net4407),
.C(net4431),
.D(net4294),
.E(net10169),
.Y(net4433)
);

AND4x2_ASAP7_75t_R c4396(
.A(net4423),
.B(net4427),
.C(net4363),
.D(net4431),
.Y(net4434)
);

NOR3x2_ASAP7_75t_R c4397(
.B(net4406),
.C(net4418),
.A(net4431),
.Y(net4435)
);

AO222x2_ASAP7_75t_R c4398(
.A1(net4424),
.A2(net4423),
.B1(net4432),
.B2(net4379),
.C1(net4386),
.C2(net4431),
.Y(net4436)
);

NOR3xp33_ASAP7_75t_R c4399(
.A(net3561),
.B(net4310),
.C(net3580),
.Y(net4437)
);

NOR2x1p5_ASAP7_75t_R c4400(
.A(net4110),
.B(net10244),
.Y(net4438)
);

SDFLx1_ASAP7_75t_R c4401(
.D(net2475),
.SE(net2668),
.SI(net9941),
.CLK(clk),
.QN(net4439)
);

INVxp67_ASAP7_75t_R c4402(
.A(net4202),
.Y(net4440)
);

NOR2x2_ASAP7_75t_R c4403(
.A(net2629),
.B(net2538),
.Y(out1)
);

NOR2xp33_ASAP7_75t_R c4404(
.A(net2538),
.B(net10198),
.Y(net4441)
);

BUFx10_ASAP7_75t_R c4405(
.A(net10155),
.Y(net4442)
);

NOR2xp67_ASAP7_75t_R c4406(
.A(net4441),
.B(net9683),
.Y(net4443)
);

OR2x2_ASAP7_75t_R c4407(
.A(net4355),
.B(net4409),
.Y(net4444)
);

OR2x4_ASAP7_75t_R c4408(
.A(net4438),
.B(net3442),
.Y(net4445)
);

BUFx12_ASAP7_75t_R c4409(
.A(net10429),
.Y(net4446)
);

BUFx12f_ASAP7_75t_R c4410(
.A(net1736),
.Y(net4447)
);

ICGx4DC_ASAP7_75t_R c4411(
.ENA(net3450),
.SE(net3580),
.CLK(clk),
.GCLK(net4448)
);

OR2x6_ASAP7_75t_R c4412(
.A(net4401),
.B(net1664),
.Y(net4449)
);

BUFx16f_ASAP7_75t_R c4413(
.A(net10117),
.Y(net4450)
);

XNOR2x1_ASAP7_75t_R c4414(
.B(net4417),
.A(net4310),
.Y(net4451)
);

XNOR2x2_ASAP7_75t_R c4415(
.A(net4450),
.B(net4446),
.Y(net4452)
);

XNOR2xp5_ASAP7_75t_R c4416(
.A(net3435),
.B(net4432),
.Y(net4453)
);

XOR2x1_ASAP7_75t_R c4417(
.A(net2668),
.B(net3360),
.Y(net4454)
);

XOR2x2_ASAP7_75t_R c4418(
.A(net667),
.B(net1664),
.Y(net4455)
);

OA21x2_ASAP7_75t_R c4419(
.A1(net3542),
.A2(net4435),
.B(net667),
.Y(net4456)
);

BUFx24_ASAP7_75t_R c4420(
.A(net10109),
.Y(net4457)
);

XOR2xp5_ASAP7_75t_R c4421(
.A(net4351),
.B(net667),
.Y(net4458)
);

OAI21x1_ASAP7_75t_R c4422(
.A1(net4451),
.A2(net4099),
.B(net10198),
.Y(net4459)
);

AND2x2_ASAP7_75t_R c4423(
.A(net3566),
.B(net790),
.Y(net4460)
);

AND2x4_ASAP7_75t_R c4424(
.A(net4409),
.B(net4454),
.Y(net4461)
);

OAI21xp33_ASAP7_75t_R c4425(
.A1(net660),
.A2(net4441),
.B(net4447),
.Y(net4462)
);

BUFx2_ASAP7_75t_R c4426(
.A(net10357),
.Y(net4463)
);

OAI21xp5_ASAP7_75t_R c4427(
.A1(net4158),
.A2(net1736),
.B(net4379),
.Y(net4464)
);

BUFx3_ASAP7_75t_R c4428(
.A(net1612),
.Y(net4465)
);

AND2x6_ASAP7_75t_R c4429(
.A(net2427),
.B(net4355),
.Y(net4466)
);

SDFLx2_ASAP7_75t_R c4430(
.D(net3591),
.SE(net750),
.SI(net1490),
.CLK(clk),
.QN(net4467)
);

HAxp5_ASAP7_75t_R c4431(
.A(net790),
.B(net4458),
.CON(net4469),
.SN(net4468)
);

NAND2x1_ASAP7_75t_R c4432(
.A(net3363),
.B(net4465),
.Y(net4470)
);

AO211x2_ASAP7_75t_R c4433(
.A1(net3552),
.A2(net2584),
.B(net4439),
.C(net10244),
.Y(net4471)
);

NAND2x1p5_ASAP7_75t_R c4434(
.A(net4454),
.B(net4462),
.Y(net4472)
);

NAND2x2_ASAP7_75t_R c4435(
.A(net775),
.B(net2661),
.Y(net4473)
);

NAND2xp33_ASAP7_75t_R c4436(
.A(net2337),
.B(net4446),
.Y(net4474)
);

BUFx4_ASAP7_75t_R c4437(
.A(net10428),
.Y(net4475)
);

NAND2xp5_ASAP7_75t_R c4438(
.A(net4455),
.B(net3578),
.Y(net4476)
);

BUFx4f_ASAP7_75t_R c4439(
.A(net10087),
.Y(net4477)
);

NAND2xp67_ASAP7_75t_R c4440(
.A(net4447),
.B(net3537),
.Y(net4478)
);

SDFLx3_ASAP7_75t_R c4441(
.D(net3585),
.SE(net4440),
.SI(net3557),
.CLK(clk),
.QN(net4479)
);

AO22x1_ASAP7_75t_R c4442(
.A1(net4457),
.A2(net2636),
.B1(net4440),
.B2(net4468),
.Y(net4480)
);

NOR2x1_ASAP7_75t_R c4443(
.A(net1709),
.B(net4210),
.Y(net4481)
);

NOR2x1p5_ASAP7_75t_R c4444(
.A(net4437),
.B(net4439),
.Y(net4482)
);

NOR2x2_ASAP7_75t_R c4445(
.A(net3360),
.B(net4478),
.Y(net4483)
);

NOR2xp33_ASAP7_75t_R c4446(
.A(net4449),
.B(net9647),
.Y(net4484)
);

OR3x1_ASAP7_75t_R c4447(
.A(net2380),
.B(net2538),
.C(net4479),
.Y(net4485)
);

NOR2xp67_ASAP7_75t_R c4448(
.A(net4463),
.B(net4483),
.Y(net4486)
);

OR2x2_ASAP7_75t_R c4449(
.A(net4463),
.B(net10169),
.Y(net4487)
);

OR3x2_ASAP7_75t_R c4450(
.A(net4482),
.B(net4476),
.C(net4425),
.Y(net4488)
);

OR2x4_ASAP7_75t_R c4451(
.A(net4459),
.B(net4481),
.Y(net4489)
);

OR3x4_ASAP7_75t_R c4452(
.A(net4486),
.B(net4487),
.C(net4446),
.Y(net4490)
);

BUFx5_ASAP7_75t_R c4453(
.A(net10364),
.Y(net4491)
);

SDFLx4_ASAP7_75t_R c4454(
.D(net4317),
.SE(net4490),
.SI(net3587),
.CLK(clk),
.QN(net4492)
);

AND3x1_ASAP7_75t_R c4455(
.A(net4443),
.B(net4492),
.C(net4447),
.Y(net4493)
);

OR2x6_ASAP7_75t_R c4456(
.A(net2605),
.B(net4492),
.Y(net4494)
);

AND3x2_ASAP7_75t_R c4457(
.A(net4471),
.B(net4417),
.C(net4479),
.Y(net4495)
);

DFFASRHQNx1_ASAP7_75t_R c4458(
.D(net4353),
.RESETN(net4487),
.SETN(net4448),
.CLK(clk),
.QN(net4496)
);

AND3x4_ASAP7_75t_R c4459(
.A(net4466),
.B(net4446),
.C(net4481),
.Y(net4497)
);

XNOR2x1_ASAP7_75t_R c4460(
.B(net4470),
.A(net4497),
.Y(net4498)
);

AO21x1_ASAP7_75t_R c4461(
.A1(net2569),
.A2(net4494),
.B(net4437),
.Y(net4499)
);

SDFHx1_ASAP7_75t_R c4462(
.D(net4490),
.SE(net1720),
.SI(net4496),
.CLK(clk),
.QN(net4500)
);

XNOR2x2_ASAP7_75t_R c4463(
.A(net4461),
.B(net4496),
.Y(net4501)
);

SDFHx2_ASAP7_75t_R c4464(
.D(net4476),
.SE(net4499),
.SI(net4501),
.CLK(clk),
.QN(net4502)
);

OA221x2_ASAP7_75t_R c4465(
.A1(net4460),
.A2(net4439),
.B1(net4502),
.B2(net3432),
.C(net4449),
.Y(net4503)
);

AO21x2_ASAP7_75t_R c4466(
.A1(net4474),
.A2(net4499),
.B(net4502),
.Y(net4504)
);

AOI21x1_ASAP7_75t_R c4467(
.A1(net4485),
.A2(net2601),
.B(net1664),
.Y(net4505)
);

AOI21xp33_ASAP7_75t_R c4468(
.A1(net4473),
.A2(net4500),
.B(net4495),
.Y(net4506)
);

AOI21xp5_ASAP7_75t_R c4469(
.A1(net4496),
.A2(net4500),
.B(net4503),
.Y(net4507)
);

XNOR2xp5_ASAP7_75t_R c4470(
.A(net4503),
.B(net4475),
.Y(net4508)
);

FAx1_ASAP7_75t_R c4471(
.A(net4508),
.B(net4507),
.CI(net3542),
.SN(net4509)
);

BUFx6f_ASAP7_75t_R c4472(
.A(net10155),
.Y(net4510)
);

MAJIxp5_ASAP7_75t_R c4473(
.A(net2636),
.B(net4444),
.C(net4487),
.Y(net4511)
);

MAJx2_ASAP7_75t_R c4474(
.A(net4506),
.B(net4449),
.C(net4463),
.Y(net4512)
);

XOR2x1_ASAP7_75t_R c4475(
.A(net4510),
.B(net4467),
.Y(net4513)
);

XOR2x2_ASAP7_75t_R c4476(
.A(net4210),
.B(net4491),
.Y(net4514)
);

MAJx3_ASAP7_75t_R c4477(
.A(net3560),
.B(net4501),
.C(net4483),
.Y(net4515)
);

AO22x2_ASAP7_75t_R c4478(
.A1(net4416),
.A2(net4500),
.B1(net4515),
.B2(net9916),
.Y(net4516)
);

NAND3x1_ASAP7_75t_R c4479(
.A(net4493),
.B(net9869),
.C(net10245),
.Y(net4517)
);

AO31x2_ASAP7_75t_R c4480(
.A1(net4514),
.A2(net4517),
.A3(net4515),
.B(net4432),
.Y(net4518)
);

AOI211x1_ASAP7_75t_R c4481(
.A1(net4512),
.A2(net4503),
.B(net4515),
.C(net9945),
.Y(net4519)
);

XOR2xp5_ASAP7_75t_R c4482(
.A(net3485),
.B(net2682),
.Y(net4520)
);

AND2x2_ASAP7_75t_R c4483(
.A(net3481),
.B(net784),
.Y(net4521)
);

AND2x4_ASAP7_75t_R c4484(
.A(net3512),
.B(net10230),
.Y(net4522)
);

AND2x6_ASAP7_75t_R c4485(
.A(net686),
.B(net1759),
.Y(net4523)
);

NAND3x2_ASAP7_75t_R c4486(
.B(net4394),
.C(net824),
.A(net10245),
.Y(net4524)
);

HAxp5_ASAP7_75t_R c4487(
.A(net2584),
.B(net3655),
.CON(net4526),
.SN(net4525)
);

NAND3xp33_ASAP7_75t_R c4488(
.A(net3617),
.B(net3655),
.C(net4495),
.Y(net4527)
);

NAND2x1_ASAP7_75t_R c4489(
.A(net4480),
.B(net2745),
.Y(net4528)
);

NOR3x1_ASAP7_75t_R c4490(
.A(net3632),
.B(net3617),
.C(net4357),
.Y(net4529)
);

SDFHx3_ASAP7_75t_R c4491(
.D(net2689),
.SE(net3660),
.SI(net3565),
.CLK(clk),
.QN(net4530)
);

NOR3x2_ASAP7_75t_R c4492(
.B(net3660),
.C(net2708),
.A(net10245),
.Y(net4531)
);

BUFx8_ASAP7_75t_R c4493(
.A(net10340),
.Y(net4532)
);

NOR3xp33_ASAP7_75t_R c4494(
.A(net3486),
.B(net2736),
.C(net3512),
.Y(net4533)
);

NAND2x1p5_ASAP7_75t_R c4495(
.A(net824),
.B(net3592),
.Y(net4534)
);

NAND2x2_ASAP7_75t_R c4496(
.A(net2714),
.B(net2735),
.Y(net4535)
);

NAND2xp33_ASAP7_75t_R c4497(
.A(net3609),
.B(net2714),
.Y(net4536)
);

OA21x2_ASAP7_75t_R c4498(
.A1(net4293),
.A2(net3633),
.B(net9794),
.Y(net4537)
);

OAI21x1_ASAP7_75t_R c4499(
.A1(net3646),
.A2(net838),
.B(net10231),
.Y(net4538)
);

OAI21xp33_ASAP7_75t_R c4500(
.A1(net3541),
.A2(net4534),
.B(net4480),
.Y(net4539)
);

NAND2xp5_ASAP7_75t_R c4501(
.A(net4472),
.B(net3628),
.Y(net4540)
);

NAND2xp67_ASAP7_75t_R c4502(
.A(net4357),
.B(net9962),
.Y(net4541)
);

CKINVDCx10_ASAP7_75t_R c4503(
.A(net10547),
.Y(net4542)
);

OAI21xp5_ASAP7_75t_R c4504(
.A1(net3611),
.A2(net3541),
.B(net3652),
.Y(net4543)
);

OR3x1_ASAP7_75t_R c4505(
.A(net2678),
.B(net3673),
.C(net3600),
.Y(net4544)
);

ICGx4_ASAP7_75t_R c4506(
.ENA(net4433),
.SE(net3565),
.CLK(clk),
.GCLK(net4545)
);

OR3x2_ASAP7_75t_R c4507(
.A(net2735),
.B(out1),
.C(net4166),
.Y(net4546)
);

AOI211xp5_ASAP7_75t_R c4508(
.A1(net4532),
.A2(net1720),
.B(net750),
.C(net10232),
.Y(net4547)
);

OR3x4_ASAP7_75t_R c4509(
.A(net750),
.B(net4530),
.C(net3600),
.Y(net4548)
);

SDFHx4_ASAP7_75t_R c4510(
.D(net3604),
.SE(net3603),
.SI(net4357),
.CLK(clk),
.QN(net4549)
);

AND3x1_ASAP7_75t_R c4511(
.A(net3656),
.B(net3640),
.C(net10234),
.Y(net4550)
);

NOR2x1_ASAP7_75t_R c4512(
.A(net876),
.B(net3650),
.Y(net4551)
);

SDFLx1_ASAP7_75t_R c4513(
.D(net2732),
.SE(net4522),
.SI(net2745),
.CLK(clk),
.QN(net4552)
);

AND3x2_ASAP7_75t_R c4514(
.A(net3592),
.B(net4534),
.C(net750),
.Y(net4553)
);

AOI22x1_ASAP7_75t_R c4515(
.A1(net4495),
.A2(net4536),
.B1(net3676),
.B2(net4552),
.Y(net4554)
);

AND3x4_ASAP7_75t_R c4516(
.A(net3663),
.B(net2707),
.C(net3512),
.Y(net4555)
);

NOR2x1p5_ASAP7_75t_R c4517(
.A(net3580),
.B(net4552),
.Y(net4556)
);

NOR2x2_ASAP7_75t_R c4518(
.A(net4544),
.B(net4521),
.Y(net4557)
);

NOR2xp33_ASAP7_75t_R c4519(
.A(net4548),
.B(net9836),
.Y(net4558)
);

AOI22xp33_ASAP7_75t_R c4520(
.A1(net4520),
.A2(net1823),
.B1(net4480),
.B2(net2747),
.Y(net4559)
);

AO21x1_ASAP7_75t_R c4521(
.A1(net1777),
.A2(net4558),
.B(net3656),
.Y(net4560)
);

OAI221xp5_ASAP7_75t_R c4522(
.A1(net3573),
.A2(net4495),
.B1(net4534),
.B2(net2617),
.C(net10246),
.Y(net4561)
);

AO21x2_ASAP7_75t_R c4523(
.A1(net2740),
.A2(net2590),
.B(net4548),
.Y(net4562)
);

AOI21x1_ASAP7_75t_R c4524(
.A1(net3484),
.A2(net2617),
.B(net9685),
.Y(net4563)
);

AOI21xp33_ASAP7_75t_R c4525(
.A1(net3640),
.A2(net3663),
.B(net2712),
.Y(net4564)
);

AOI21xp5_ASAP7_75t_R c4526(
.A1(net4548),
.A2(net4560),
.B(net3643),
.Y(net4565)
);

SDFLx2_ASAP7_75t_R c4527(
.D(net3666),
.SE(net4293),
.SI(net839),
.CLK(clk),
.QN(net4566)
);

NOR2xp67_ASAP7_75t_R c4528(
.A(net3646),
.B(net4552),
.Y(net4567)
);

CKINVDCx11_ASAP7_75t_R c4529(
.A(net10340),
.Y(net4568)
);

FAx1_ASAP7_75t_R c4530(
.A(net4527),
.B(net3619),
.CI(net4307),
.SN(net4569)
);

AO33x2_ASAP7_75t_R c4531(
.A1(net3603),
.A2(net3622),
.A3(net4552),
.B1(net3640),
.B2(net3604),
.B3(net3655),
.Y(net4570)
);

OR2x2_ASAP7_75t_R c4532(
.A(net4545),
.B(net1823),
.Y(net4571)
);

OR2x4_ASAP7_75t_R c4533(
.A(net1769),
.B(net2642),
.Y(net4572)
);

OR2x6_ASAP7_75t_R c4534(
.A(net9772),
.B(net10247),
.Y(net4573)
);

XNOR2x1_ASAP7_75t_R c4535(
.B(net3878),
.A(net4567),
.Y(net4574)
);

SDFLx3_ASAP7_75t_R c4536(
.D(net3480),
.SE(net4550),
.SI(net2691),
.CLK(clk),
.QN(net4575)
);

XNOR2x2_ASAP7_75t_R c4537(
.A(net3484),
.B(net4575),
.Y(net4576)
);

MAJIxp5_ASAP7_75t_R c4538(
.A(net3532),
.B(net686),
.C(net10234),
.Y(net4577)
);

MAJx2_ASAP7_75t_R c4539(
.A(net3633),
.B(net4529),
.C(net4573),
.Y(net4578)
);

MAJx3_ASAP7_75t_R c4540(
.A(net3599),
.B(net4573),
.C(net4540),
.Y(net4579)
);

NAND3x1_ASAP7_75t_R c4541(
.A(net4551),
.B(net4530),
.C(net10247),
.Y(net4580)
);

NAND3x2_ASAP7_75t_R c4542(
.B(net4552),
.C(net10232),
.A(net10246),
.Y(net4581)
);

AOI222xp33_ASAP7_75t_R c4543(
.A1(net2691),
.A2(net4469),
.B1(net4572),
.B2(net2689),
.C1(net4573),
.C2(net10246),
.Y(net4582)
);

SDFLx4_ASAP7_75t_R c4544(
.D(net4567),
.SE(net2747),
.SI(net4552),
.CLK(clk),
.QN(net4583)
);

NAND3xp33_ASAP7_75t_R c4545(
.A(net4541),
.B(net4577),
.C(net4545),
.Y(net4584)
);

NOR3x1_ASAP7_75t_R c4546(
.A(net4548),
.B(net9937),
.C(net10247),
.Y(net4585)
);

NOR3x2_ASAP7_75t_R c4547(
.B(net3629),
.C(net4542),
.A(net784),
.Y(net4586)
);

NOR3xp33_ASAP7_75t_R c4548(
.A(net4574),
.B(net4586),
.C(net10248),
.Y(net4587)
);

OA21x2_ASAP7_75t_R c4549(
.A1(net3239),
.A2(net4530),
.B(net803),
.Y(net4588)
);

OAI21x1_ASAP7_75t_R c4550(
.A1(net4524),
.A2(net4583),
.B(net9937),
.Y(net4589)
);

OAI21xp33_ASAP7_75t_R c4551(
.A1(net4528),
.A2(net4553),
.B(net4575),
.Y(net4590)
);

DFFASRHQNx1_ASAP7_75t_R c4552(
.D(net3636),
.RESETN(net3604),
.SETN(net3666),
.CLK(clk),
.QN(net4591)
);

SDFHx1_ASAP7_75t_R c4553(
.D(net1785),
.SE(net4575),
.SI(net4573),
.CLK(clk),
.QN(net4592)
);

SDFHx2_ASAP7_75t_R c4554(
.D(net4581),
.SE(net4589),
.SI(net9685),
.CLK(clk),
.QN(net4593)
);

SDFHx3_ASAP7_75t_R c4555(
.D(net2736),
.SE(net2747),
.SI(net3676),
.CLK(clk),
.QN(net4594)
);

OAI21xp5_ASAP7_75t_R c4556(
.A1(net4534),
.A2(net4568),
.B(net4566),
.Y(net4595)
);

OR3x1_ASAP7_75t_R c4557(
.A(net4562),
.B(net9754),
.C(net9962),
.Y(net4596)
);

AOI321xp33_ASAP7_75t_R c4558(
.A1(net1817),
.A2(net4592),
.A3(net4572),
.B1(net4573),
.B2(net3655),
.C(net3626),
.Y(net4597)
);

OR3x2_ASAP7_75t_R c4559(
.A(net784),
.B(net4567),
.C(net4594),
.Y(net4598)
);

SDFHx4_ASAP7_75t_R c4560(
.D(net4561),
.SE(net4596),
.SI(net4575),
.CLK(clk),
.QN(net4599)
);

OR3x4_ASAP7_75t_R c4561(
.A(net4599),
.B(net4587),
.C(net4594),
.Y(net4600)
);

AND3x1_ASAP7_75t_R c4562(
.A(net4547),
.B(net4592),
.C(net9892),
.Y(net4601)
);

AND3x2_ASAP7_75t_R c4563(
.A(net4601),
.B(net4599),
.C(net3618),
.Y(net4602)
);

AND3x4_ASAP7_75t_R c4564(
.A(net3565),
.B(net4600),
.C(net9815),
.Y(net4603)
);

CKINVDCx12_ASAP7_75t_R c4565(
.A(net3682),
.Y(net4604)
);

CKINVDCx14_ASAP7_75t_R c4566(
.A(net3751),
.Y(net4605)
);

CKINVDCx16_ASAP7_75t_R c4567(
.A(net3709),
.Y(net4606)
);

CKINVDCx20_ASAP7_75t_R c4568(
.A(net3702),
.Y(net4607)
);

XNOR2xp5_ASAP7_75t_R c4569(
.A(net1891),
.B(net3755),
.Y(net4608)
);

CKINVDCx5p33_ASAP7_75t_R c4570(
.A(net3700),
.Y(net4609)
);

CKINVDCx6p67_ASAP7_75t_R c4571(
.A(net975),
.Y(net4610)
);

CKINVDCx8_ASAP7_75t_R c4572(
.A(net1892),
.Y(net4611)
);

XOR2x1_ASAP7_75t_R c4573(
.A(net1827),
.B(in24),
.Y(net4612)
);

CKINVDCx9p33_ASAP7_75t_R c4574(
.A(net980),
.Y(net4613)
);

HB1xp67_ASAP7_75t_R c4575(
.A(net3716),
.Y(net4614)
);

HB2xp67_ASAP7_75t_R c4576(
.A(net3755),
.Y(net4615)
);

HB3xp67_ASAP7_75t_R c4577(
.A(net3746),
.Y(net4616)
);

HB4xp67_ASAP7_75t_R c4578(
.A(net1844),
.Y(net4617)
);

INVx11_ASAP7_75t_R c4579(
.A(in7),
.Y(net4618)
);

INVx13_ASAP7_75t_R c4580(
.A(net3699),
.Y(net4619)
);

INVx1_ASAP7_75t_R c4581(
.A(net4612),
.Y(net4620)
);

INVx2_ASAP7_75t_R c4582(
.A(net3726),
.Y(net4621)
);

XOR2x2_ASAP7_75t_R c4583(
.A(net3706),
.B(net3745),
.Y(net4622)
);

INVx3_ASAP7_75t_R c4584(
.A(net3733),
.Y(net4623)
);

INVx4_ASAP7_75t_R c4585(
.A(net1869),
.Y(net4624)
);

INVx5_ASAP7_75t_R c4586(
.A(net2810),
.Y(net4625)
);

INVx6_ASAP7_75t_R c4587(
.A(net3706),
.Y(net4626)
);

XOR2xp5_ASAP7_75t_R c4588(
.A(net4614),
.B(net4626),
.Y(net4627)
);

INVx8_ASAP7_75t_R c4589(
.A(net2792),
.Y(net4628)
);

INVxp33_ASAP7_75t_R c4590(
.A(net4622),
.Y(net4629)
);

INVxp67_ASAP7_75t_R c4591(
.A(net4620),
.Y(net4630)
);

AND2x2_ASAP7_75t_R c4592(
.A(in24),
.B(net3706),
.Y(net4631)
);

BUFx10_ASAP7_75t_R c4593(
.A(net4605),
.Y(net4632)
);

AND2x4_ASAP7_75t_R c4594(
.A(net4606),
.B(net4630),
.Y(net4633)
);

BUFx12_ASAP7_75t_R c4595(
.A(net3709),
.Y(net4634)
);

AND2x6_ASAP7_75t_R c4596(
.A(net4627),
.B(net2775),
.Y(net4635)
);

BUFx12f_ASAP7_75t_R c4597(
.A(net4632),
.Y(net4636)
);

HAxp5_ASAP7_75t_R c4598(
.A(net4629),
.B(net3760),
.CON(net4638),
.SN(net4637)
);

NAND2x1_ASAP7_75t_R c4599(
.A(net4623),
.B(net4628),
.Y(net4639)
);

AO21x1_ASAP7_75t_R c4600(
.A1(net4630),
.A2(net4631),
.B(net4628),
.Y(net4640)
);

BUFx16f_ASAP7_75t_R c4601(
.A(net9088),
.Y(net4641)
);

BUFx24_ASAP7_75t_R c4602(
.A(net3713),
.Y(net4642)
);

NAND2x1p5_ASAP7_75t_R c4603(
.A(net4621),
.B(net4633),
.Y(net4643)
);

NAND2x2_ASAP7_75t_R c4604(
.A(net4628),
.B(net4615),
.Y(net4644)
);

BUFx2_ASAP7_75t_R c4605(
.A(net4631),
.Y(net4645)
);

AO21x2_ASAP7_75t_R c4606(
.A1(net4617),
.A2(net4620),
.B(net4640),
.Y(net4646)
);

NAND2xp33_ASAP7_75t_R c4607(
.A(net2792),
.B(net4644),
.Y(net4647)
);

AOI21x1_ASAP7_75t_R c4608(
.A1(net4634),
.A2(net3725),
.B(net4611),
.Y(net4648)
);

AOI21xp33_ASAP7_75t_R c4609(
.A1(net4623),
.A2(net4626),
.B(net4634),
.Y(net4649)
);

NAND2xp5_ASAP7_75t_R c4610(
.A(net4640),
.B(net4612),
.Y(net4650)
);

BUFx3_ASAP7_75t_R c4611(
.A(net2823),
.Y(net4651)
);

ICGx5_ASAP7_75t_R c4612(
.ENA(net4637),
.SE(net4648),
.CLK(clk),
.GCLK(net4652)
);

BUFx4_ASAP7_75t_R c4613(
.A(net4636),
.Y(net4653)
);

NAND2xp67_ASAP7_75t_R c4614(
.A(net4643),
.B(net4636),
.Y(net4654)
);

NOR2x1_ASAP7_75t_R c4615(
.A(net4632),
.B(net4633),
.Y(net4655)
);

NOR2x1p5_ASAP7_75t_R c4616(
.A(net4648),
.B(net4606),
.Y(net4656)
);

NOR2x2_ASAP7_75t_R c4617(
.A(net4653),
.B(net4642),
.Y(net4657)
);

BUFx4f_ASAP7_75t_R c4618(
.A(net9088),
.Y(net4658)
);

NOR2xp33_ASAP7_75t_R c4619(
.A(net4605),
.B(net3755),
.Y(net4659)
);

NOR2xp67_ASAP7_75t_R c4620(
.A(net4659),
.B(net4645),
.Y(net4660)
);

OR2x2_ASAP7_75t_R c4621(
.A(net4607),
.B(net3751),
.Y(net4661)
);

OR2x4_ASAP7_75t_R c4622(
.A(net4649),
.B(net3751),
.Y(net4662)
);

OR2x6_ASAP7_75t_R c4623(
.A(net4640),
.B(net4662),
.Y(net4663)
);

XNOR2x1_ASAP7_75t_R c4624(
.B(net3725),
.A(net4663),
.Y(net4664)
);

XNOR2x2_ASAP7_75t_R c4625(
.A(net4622),
.B(net4625),
.Y(net4665)
);

AOI21xp5_ASAP7_75t_R c4626(
.A1(net4645),
.A2(net4608),
.B(net4623),
.Y(net4666)
);

FAx1_ASAP7_75t_R c4627(
.A(net4658),
.B(net3733),
.CI(net4666),
.SN(net4668),
.CON(net4667)
);

XNOR2xp5_ASAP7_75t_R c4628(
.A(net4664),
.B(net4665),
.Y(net4669)
);

XOR2x1_ASAP7_75t_R c4629(
.A(net3685),
.B(net4634),
.Y(net4670)
);

XOR2x2_ASAP7_75t_R c4630(
.A(net4661),
.B(net4662),
.Y(net4671)
);

MAJIxp5_ASAP7_75t_R c4631(
.A(net4614),
.B(net4656),
.C(net9727),
.Y(net4672)
);

ICGx5p33DC_ASAP7_75t_R c4632(
.ENA(net3726),
.SE(net4670),
.CLK(clk),
.GCLK(net4673)
);

AOI33xp33_ASAP7_75t_R c4633(
.A1(net4659),
.A2(net4626),
.A3(net4664),
.B1(net4673),
.B2(net4650),
.B3(net3701),
.Y(net4674)
);

AOI22xp5_ASAP7_75t_R c4634(
.A1(net4604),
.A2(net4641),
.B1(net4670),
.B2(net3747),
.Y(net4675)
);

MAJx2_ASAP7_75t_R c4635(
.A(net4673),
.B(net4647),
.C(net4628),
.Y(net4676)
);

MAJx3_ASAP7_75t_R c4636(
.A(net4662),
.B(net4672),
.C(net4639),
.Y(net4677)
);

XOR2xp5_ASAP7_75t_R c4637(
.A(net4641),
.B(net4671),
.Y(net4678)
);

AND2x2_ASAP7_75t_R c4638(
.A(net4673),
.B(net9727),
.Y(net4679)
);

AOI31xp33_ASAP7_75t_R c4639(
.A1(net4615),
.A2(net4653),
.A3(net4623),
.B(net3699),
.Y(net4680)
);

AND2x4_ASAP7_75t_R c4640(
.A(net4680),
.B(net3705),
.Y(net4681)
);

AOI31xp67_ASAP7_75t_R c4641(
.A1(net4670),
.A2(net4678),
.A3(net4643),
.B(net4681),
.Y(net4682)
);

OA222x2_ASAP7_75t_R c4642(
.A1(net4677),
.A2(net4663),
.B1(net4621),
.B2(net4656),
.C1(net3701),
.C2(net10250),
.Y(net4683)
);

AND2x6_ASAP7_75t_R c4643(
.A(net4666),
.B(net4662),
.Y(net4684)
);

HAxp5_ASAP7_75t_R c4644(
.A(net4672),
.B(net4671),
.CON(net4686),
.SN(net4685)
);

SDFLx1_ASAP7_75t_R c4645(
.D(net4680),
.SE(net4686),
.SI(net10251),
.CLK(clk),
.QN(net4687)
);

SDFLx2_ASAP7_75t_R c4646(
.D(net4686),
.SE(net10249),
.SI(net10251),
.CLK(clk),
.QN(net4688)
);

OAI311xp33_ASAP7_75t_R c4647(
.A1(net4684),
.A2(net4654),
.A3(net4685),
.B1(net4681),
.C1(net4613),
.Y(net4689)
);

NAND2x1_ASAP7_75t_R c4648(
.A(net3776),
.B(net2841),
.Y(net4690)
);

NAND3x1_ASAP7_75t_R c4649(
.A(net3809),
.B(net4646),
.C(net4633),
.Y(net4691)
);

BUFx5_ASAP7_75t_R c4650(
.A(net3812),
.Y(net4692)
);

NAND3x2_ASAP7_75t_R c4651(
.B(net1954),
.C(net2775),
.A(net3776),
.Y(net4693)
);

BUFx6f_ASAP7_75t_R c4652(
.A(net4633),
.Y(net4694)
);

NAND2x1p5_ASAP7_75t_R c4653(
.A(net3764),
.B(net3766),
.Y(net4695)
);

BUFx8_ASAP7_75t_R c4654(
.A(net3789),
.Y(net4696)
);

CKINVDCx10_ASAP7_75t_R c4655(
.A(net1989),
.Y(net4697)
);

CKINVDCx11_ASAP7_75t_R c4656(
.A(net10562),
.Y(net4698)
);

CKINVDCx12_ASAP7_75t_R c4657(
.A(net4697),
.Y(net4699)
);

CKINVDCx14_ASAP7_75t_R c4658(
.A(net4694),
.Y(net4700)
);

CKINVDCx16_ASAP7_75t_R c4659(
.A(net9176),
.Y(net4701)
);

NAND2x2_ASAP7_75t_R c4660(
.A(net4627),
.B(net3705),
.Y(net4702)
);

CKINVDCx20_ASAP7_75t_R c4661(
.A(net3680),
.Y(net4703)
);

NAND2xp33_ASAP7_75t_R c4662(
.A(net2885),
.B(net4646),
.Y(net4704)
);

CKINVDCx5p33_ASAP7_75t_R c4663(
.A(net9201),
.Y(net4705)
);

CKINVDCx6p67_ASAP7_75t_R c4664(
.A(net3792),
.Y(net4706)
);

CKINVDCx8_ASAP7_75t_R c4665(
.A(net4698),
.Y(net4707)
);

NAND2xp5_ASAP7_75t_R c4666(
.A(net2841),
.B(net2913),
.Y(net4708)
);

CKINVDCx9p33_ASAP7_75t_R c4667(
.A(net4699),
.Y(net4709)
);

ICGx6p67DC_ASAP7_75t_R c4668(
.ENA(net4638),
.SE(net4639),
.CLK(clk),
.GCLK(net4710)
);

HB1xp67_ASAP7_75t_R c4669(
.A(net9935),
.Y(net4711)
);

SDFLx3_ASAP7_75t_R c4670(
.D(net4693),
.SE(net4709),
.SI(net4706),
.CLK(clk),
.QN(net4712)
);

HB2xp67_ASAP7_75t_R c4671(
.A(net3810),
.Y(net4713)
);

HB3xp67_ASAP7_75t_R c4672(
.A(net4679),
.Y(net4714)
);

HB4xp67_ASAP7_75t_R c4673(
.A(net4702),
.Y(net4715)
);

NAND2xp67_ASAP7_75t_R c4674(
.A(net4647),
.B(net4663),
.Y(net4716)
);

SDFLx4_ASAP7_75t_R c4675(
.D(net4663),
.SE(net1974),
.SI(net4691),
.CLK(clk),
.QN(net4717)
);

INVx11_ASAP7_75t_R c4676(
.A(net2823),
.Y(net4718)
);

NOR2x1_ASAP7_75t_R c4677(
.A(net4713),
.B(net4711),
.Y(net4719)
);

NOR2x1p5_ASAP7_75t_R c4678(
.A(net4688),
.B(net4663),
.Y(net4720)
);

INVx13_ASAP7_75t_R c4679(
.A(net4703),
.Y(net4721)
);

NOR2x2_ASAP7_75t_R c4680(
.A(net2775),
.B(net3739),
.Y(net4722)
);

INVx1_ASAP7_75t_R c4681(
.A(net1844),
.Y(net4723)
);

NOR2xp33_ASAP7_75t_R c4682(
.A(net4687),
.B(net3782),
.Y(net4724)
);

NOR2xp67_ASAP7_75t_R c4683(
.A(net4712),
.B(net4710),
.Y(net4725)
);

OR2x2_ASAP7_75t_R c4684(
.A(net4725),
.B(net1988),
.Y(net4726)
);

INVx2_ASAP7_75t_R c4685(
.A(net4673),
.Y(net4727)
);

INVx3_ASAP7_75t_R c4686(
.A(net4721),
.Y(net4728)
);

INVx4_ASAP7_75t_R c4687(
.A(net4719),
.Y(net4729)
);

INVx5_ASAP7_75t_R c4688(
.A(net1961),
.Y(net4730)
);

OR2x4_ASAP7_75t_R c4689(
.A(net4707),
.B(net4726),
.Y(net4731)
);

ICGx8DC_ASAP7_75t_R c4690(
.ENA(net4704),
.SE(net4724),
.CLK(clk),
.GCLK(net4732)
);

OR2x6_ASAP7_75t_R c4691(
.A(net4731),
.B(net4613),
.Y(net4733)
);

XNOR2x1_ASAP7_75t_R c4692(
.B(net4690),
.A(net4733),
.Y(net4734)
);

INVx6_ASAP7_75t_R c4693(
.A(net10482),
.Y(net4735)
);

INVx8_ASAP7_75t_R c4694(
.A(net4626),
.Y(net4736)
);

NAND3xp33_ASAP7_75t_R c4695(
.A(net4726),
.B(net4706),
.C(net4712),
.Y(net4737)
);

DFFASRHQNx1_ASAP7_75t_R c4696(
.D(net4729),
.RESETN(net2877),
.SETN(net4715),
.CLK(clk),
.QN(net4738)
);

NOR3x1_ASAP7_75t_R c4697(
.A(net2913),
.B(net4671),
.C(net4724),
.Y(net4739)
);

INVxp33_ASAP7_75t_R c4698(
.A(net9176),
.Y(net4740)
);

XNOR2x2_ASAP7_75t_R c4699(
.A(net4628),
.B(net9870),
.Y(net4741)
);

ICGx1_ASAP7_75t_R c4700(
.ENA(net4730),
.SE(net4688),
.CLK(clk),
.GCLK(net4742)
);

INVxp67_ASAP7_75t_R c4701(
.A(net9684),
.Y(net4743)
);

XNOR2xp5_ASAP7_75t_R c4702(
.A(net4691),
.B(net4613),
.Y(net4744)
);

BUFx10_ASAP7_75t_R c4703(
.A(net10472),
.Y(net4745)
);

BUFx12_ASAP7_75t_R c4704(
.A(net4737),
.Y(net4746)
);

XOR2x1_ASAP7_75t_R c4705(
.A(net4733),
.B(net4734),
.Y(net4747)
);

NOR3x2_ASAP7_75t_R c4706(
.B(net4745),
.C(net4702),
.A(net4730),
.Y(net4748)
);

XOR2x2_ASAP7_75t_R c4707(
.A(net4727),
.B(net3739),
.Y(net4749)
);

XOR2xp5_ASAP7_75t_R c4708(
.A(net4712),
.B(net9807),
.Y(net4750)
);

BUFx12f_ASAP7_75t_R c4709(
.A(net4718),
.Y(net4751)
);

BUFx16f_ASAP7_75t_R c4710(
.A(net4751),
.Y(net4752)
);

AND2x2_ASAP7_75t_R c4711(
.A(net4613),
.B(net4741),
.Y(net4753)
);

NOR3xp33_ASAP7_75t_R c4712(
.A(net4750),
.B(net4742),
.C(net4711),
.Y(net4754)
);

BUFx24_ASAP7_75t_R c4713(
.A(net10406),
.Y(net4755)
);

AND2x4_ASAP7_75t_R c4714(
.A(net4723),
.B(net4714),
.Y(net4756)
);

AND2x6_ASAP7_75t_R c4715(
.A(net4753),
.B(net4733),
.Y(net4757)
);

BUFx2_ASAP7_75t_R c4716(
.A(net9935),
.Y(net4758)
);

HAxp5_ASAP7_75t_R c4717(
.A(net4741),
.B(net4645),
.CON(net4760),
.SN(net4759)
);

OA21x2_ASAP7_75t_R c4718(
.A1(net4755),
.A2(net3790),
.B(net9978),
.Y(net4761)
);

NAND2x1_ASAP7_75t_R c4719(
.A(net4760),
.B(net4752),
.Y(net4762)
);

NAND2x1p5_ASAP7_75t_R c4720(
.A(net4752),
.B(net4738),
.Y(net4763)
);

NAND2x2_ASAP7_75t_R c4721(
.A(net4756),
.B(net4713),
.Y(net4764)
);

NAND2xp33_ASAP7_75t_R c4722(
.A(net4709),
.B(net3813),
.Y(net4765)
);

OAI21x1_ASAP7_75t_R c4723(
.A1(net3682),
.A2(net4733),
.B(net4755),
.Y(net4766)
);

OA33x2_ASAP7_75t_R c4724(
.A1(net4725),
.A2(net4766),
.A3(net4697),
.B1(net4738),
.B2(net2877),
.B3(net4733),
.Y(net4767)
);

NAND2xp5_ASAP7_75t_R c4725(
.A(net4764),
.B(net4752),
.Y(net4768)
);

SDFHx1_ASAP7_75t_R c4726(
.D(net4757),
.SE(net4750),
.SI(net3699),
.CLK(clk),
.QN(net4769)
);

NAND2xp67_ASAP7_75t_R c4727(
.A(net4768),
.B(net4742),
.Y(net4770)
);

OAI21xp33_ASAP7_75t_R c4728(
.A1(net4765),
.A2(net4687),
.B(net9935),
.Y(net4771)
);

OAI222xp33_ASAP7_75t_R c4729(
.A1(net4765),
.A2(net4770),
.B1(net4738),
.B2(net3772),
.C1(net4707),
.C2(net9684),
.Y(net4772)
);

SDFHx2_ASAP7_75t_R c4730(
.D(net4639),
.SE(net4770),
.SI(net4768),
.CLK(clk),
.QN(net4773)
);

NOR2x1_ASAP7_75t_R c4731(
.A(net2991),
.B(net1861),
.Y(net4774)
);

NOR2x1p5_ASAP7_75t_R c4732(
.A(net2022),
.B(net4735),
.Y(net4775)
);

NOR2x2_ASAP7_75t_R c4733(
.A(net3926),
.B(net4775),
.Y(net4776)
);

NOR2xp33_ASAP7_75t_R c4734(
.A(net3705),
.B(net10190),
.Y(net4777)
);

NOR2xp67_ASAP7_75t_R c4735(
.A(net4695),
.B(net3804),
.Y(net4778)
);

BUFx3_ASAP7_75t_R c4736(
.A(net1957),
.Y(net4779)
);

BUFx4_ASAP7_75t_R c4737(
.A(net2779),
.Y(net4780)
);

BUFx4f_ASAP7_75t_R c4738(
.A(net4611),
.Y(net4781)
);

BUFx5_ASAP7_75t_R c4739(
.A(net3821),
.Y(net4782)
);

BUFx6f_ASAP7_75t_R c4740(
.A(net10567),
.Y(net4783)
);

BUFx8_ASAP7_75t_R c4741(
.A(net2934),
.Y(net4784)
);

OR2x2_ASAP7_75t_R c4742(
.A(net4777),
.B(net4706),
.Y(net4785)
);

CKINVDCx10_ASAP7_75t_R c4743(
.A(net4775),
.Y(net4786)
);

OR2x4_ASAP7_75t_R c4744(
.A(net4781),
.B(net4717),
.Y(net4787)
);

OR2x6_ASAP7_75t_R c4745(
.A(net3790),
.B(net10113),
.Y(net4788)
);

XNOR2x1_ASAP7_75t_R c4746(
.B(net4779),
.A(net2022),
.Y(net4789)
);

CKINVDCx11_ASAP7_75t_R c4747(
.A(net10387),
.Y(net4790)
);

CKINVDCx12_ASAP7_75t_R c4748(
.A(net3901),
.Y(net4791)
);

CKINVDCx14_ASAP7_75t_R c4749(
.A(net4787),
.Y(net4792)
);

CKINVDCx16_ASAP7_75t_R c4750(
.A(net9827),
.Y(net4793)
);

XNOR2x2_ASAP7_75t_R c4751(
.A(net2052),
.B(net3854),
.Y(net4794)
);

CKINVDCx20_ASAP7_75t_R c4752(
.A(net3776),
.Y(net4795)
);

CKINVDCx5p33_ASAP7_75t_R c4753(
.A(net4794),
.Y(net4796)
);

OAI21xp5_ASAP7_75t_R c4754(
.A1(net4608),
.A2(net4795),
.B(net3813),
.Y(net4797)
);

XNOR2xp5_ASAP7_75t_R c4755(
.A(net4785),
.B(net4795),
.Y(net4798)
);

CKINVDCx6p67_ASAP7_75t_R c4756(
.A(net9169),
.Y(net4799)
);

CKINVDCx8_ASAP7_75t_R c4757(
.A(net4776),
.Y(net4800)
);

CKINVDCx9p33_ASAP7_75t_R c4758(
.A(net9966),
.Y(net4801)
);

HB1xp67_ASAP7_75t_R c4759(
.A(net4796),
.Y(net4802)
);

XOR2x1_ASAP7_75t_R c4760(
.A(net3873),
.B(net4795),
.Y(net4803)
);

HB2xp67_ASAP7_75t_R c4761(
.A(net4776),
.Y(net4804)
);

XOR2x2_ASAP7_75t_R c4762(
.A(net4646),
.B(net4802),
.Y(net4805)
);

HB3xp67_ASAP7_75t_R c4763(
.A(net2810),
.Y(net4806)
);

HB4xp67_ASAP7_75t_R c4764(
.A(net9169),
.Y(net4807)
);

INVx11_ASAP7_75t_R c4765(
.A(net10438),
.Y(net4808)
);

OR3x1_ASAP7_75t_R c4766(
.A(net4786),
.B(net4746),
.C(net4806),
.Y(net4809)
);

INVx13_ASAP7_75t_R c4767(
.A(net4806),
.Y(net4810)
);

XOR2xp5_ASAP7_75t_R c4768(
.A(net4810),
.B(net4802),
.Y(net4811)
);

OR3x2_ASAP7_75t_R c4769(
.A(net4795),
.B(net4794),
.C(net4650),
.Y(net4812)
);

SDFHx3_ASAP7_75t_R c4770(
.D(net3790),
.SE(net4797),
.SI(net3903),
.CLK(clk),
.QN(net4813)
);

AND2x2_ASAP7_75t_R c4771(
.A(net3911),
.B(net10016),
.Y(net4814)
);

OAI32xp33_ASAP7_75t_R c4772(
.A1(net4717),
.A2(net4794),
.A3(net3760),
.B1(net4770),
.B2(net4796),
.Y(net4815)
);

AND2x4_ASAP7_75t_R c4773(
.A(net4808),
.B(net4712),
.Y(net4816)
);

AND2x6_ASAP7_75t_R c4774(
.A(net4799),
.B(net4773),
.Y(net4817)
);

INVx1_ASAP7_75t_R c4775(
.A(net10564),
.Y(net4818)
);

HAxp5_ASAP7_75t_R c4776(
.A(net4803),
.B(net4806),
.CON(net4819)
);

OR3x4_ASAP7_75t_R c4777(
.A(net4679),
.B(net3892),
.C(net4793),
.Y(net4820)
);

INVx2_ASAP7_75t_R c4778(
.A(net3927),
.Y(net4821)
);

NAND2x1_ASAP7_75t_R c4779(
.A(net4804),
.B(net4796),
.Y(net4822)
);

AND3x1_ASAP7_75t_R c4780(
.A(net4811),
.B(net3906),
.C(net4702),
.Y(net4823)
);

NAND2x1p5_ASAP7_75t_R c4781(
.A(net3903),
.B(net4714),
.Y(net4824)
);

NAND2x2_ASAP7_75t_R c4782(
.A(net4801),
.B(net3906),
.Y(net4825)
);

INVx3_ASAP7_75t_R c4783(
.A(net9242),
.Y(net4826)
);

SDFHx4_ASAP7_75t_R c4784(
.D(net4811),
.SE(net2954),
.SI(net9663),
.CLK(clk),
.QN(net4827)
);

INVx4_ASAP7_75t_R c4785(
.A(net4825),
.Y(net4828)
);

INVx5_ASAP7_75t_R c4786(
.A(net4819),
.Y(net4829)
);

OR5x1_ASAP7_75t_R c4787(
.A(net4829),
.B(net4796),
.C(net4811),
.D(net4806),
.E(net3922),
.Y(net4830)
);

INVx6_ASAP7_75t_R c4788(
.A(net9242),
.Y(net4831)
);

AND3x2_ASAP7_75t_R c4789(
.A(net4820),
.B(net4695),
.C(net4813),
.Y(net4832)
);

OR5x2_ASAP7_75t_R c4790(
.A(net4796),
.B(net2999),
.C(net4789),
.D(net2934),
.E(net4793),
.Y(net4833)
);

INVx8_ASAP7_75t_R c4791(
.A(net2954),
.Y(net4834)
);

SDFLx1_ASAP7_75t_R c4792(
.D(net4701),
.SE(net4827),
.SI(net4828),
.CLK(clk),
.QN(net4835)
);

INVxp33_ASAP7_75t_R c4793(
.A(net4790),
.Y(net4836)
);

INVxp67_ASAP7_75t_R c4794(
.A(net4831),
.Y(net4837)
);

BUFx10_ASAP7_75t_R c4795(
.A(net4779),
.Y(net4838)
);

BUFx12_ASAP7_75t_R c4796(
.A(net10418),
.Y(net4839)
);

BUFx12f_ASAP7_75t_R c4797(
.A(net4839),
.Y(net4840)
);

AND3x4_ASAP7_75t_R c4798(
.A(net3766),
.B(net4776),
.C(net4816),
.Y(net4841)
);

NAND2xp33_ASAP7_75t_R c4799(
.A(net4837),
.B(net4793),
.Y(net4842)
);

BUFx16f_ASAP7_75t_R c4800(
.A(net9201),
.Y(net4843)
);

BUFx24_ASAP7_75t_R c4801(
.A(net10039),
.Y(net4844)
);

SDFLx2_ASAP7_75t_R c4802(
.D(net4842),
.SE(net4828),
.SI(net4843),
.CLK(clk),
.QN(net4845)
);

NAND2xp5_ASAP7_75t_R c4803(
.A(net4838),
.B(net4843),
.Y(net4846)
);

NAND2xp67_ASAP7_75t_R c4804(
.A(net4841),
.B(net4788),
.Y(net4847)
);

AO21x1_ASAP7_75t_R c4805(
.A1(net4782),
.A2(net3908),
.B(net4840),
.Y(net4848)
);

BUFx2_ASAP7_75t_R c4806(
.A(net10560),
.Y(net4849)
);

AO21x2_ASAP7_75t_R c4807(
.A1(net4791),
.A2(net4837),
.B(net9845),
.Y(net4850)
);

AOI21x1_ASAP7_75t_R c4808(
.A1(net4850),
.A2(net4806),
.B(net4611),
.Y(net4851)
);

NOR2x1_ASAP7_75t_R c4809(
.A(net3927),
.B(net10013),
.Y(net4852)
);

BUFx3_ASAP7_75t_R c4810(
.A(net10387),
.Y(net4853)
);

AOI21xp33_ASAP7_75t_R c4811(
.A1(net4608),
.A2(net4852),
.B(net9909),
.Y(net4854)
);

BUFx4_ASAP7_75t_R c4812(
.A(net10039),
.Y(net4855)
);

AOI21xp5_ASAP7_75t_R c4813(
.A1(net4855),
.A2(net4827),
.B(net4842),
.Y(net4856)
);

BUFx4f_ASAP7_75t_R c4814(
.A(net10079),
.Y(net4857)
);

NOR2x1p5_ASAP7_75t_R c4815(
.A(net3976),
.B(net4818),
.Y(net4858)
);

NOR2x2_ASAP7_75t_R c4816(
.A(net3881),
.B(net3034),
.Y(net4859)
);

BUFx5_ASAP7_75t_R c4817(
.A(net3892),
.Y(net4860)
);

NOR2xp33_ASAP7_75t_R c4818(
.A(net4742),
.B(net1229),
.Y(net4861)
);

NOR2xp67_ASAP7_75t_R c4819(
.A(net4799),
.B(net4857),
.Y(net4862)
);

OR2x2_ASAP7_75t_R c4820(
.A(net3990),
.B(net3941),
.Y(net4863)
);

OR2x4_ASAP7_75t_R c4821(
.A(net3782),
.B(net2984),
.Y(net4864)
);

BUFx6f_ASAP7_75t_R c4822(
.A(net3974),
.Y(net4865)
);

OR2x6_ASAP7_75t_R c4823(
.A(net4702),
.B(net4738),
.Y(net4866)
);

SDFLx3_ASAP7_75t_R c4824(
.D(net4774),
.SE(net3087),
.SI(net3015),
.CLK(clk),
.QN(net4867)
);

BUFx8_ASAP7_75t_R c4825(
.A(net3906),
.Y(net4868)
);

CKINVDCx10_ASAP7_75t_R c4826(
.A(net10019),
.Y(net4869)
);

XNOR2x1_ASAP7_75t_R c4827(
.B(net4865),
.A(net10019),
.Y(net4870)
);

XNOR2x2_ASAP7_75t_R c4828(
.A(net3848),
.B(net4722),
.Y(net4871)
);

CKINVDCx11_ASAP7_75t_R c4829(
.A(net3902),
.Y(net4872)
);

XNOR2xp5_ASAP7_75t_R c4830(
.A(net3930),
.B(net3708),
.Y(net4873)
);

XOR2x1_ASAP7_75t_R c4831(
.A(net4865),
.B(net2983),
.Y(net4874)
);

XOR2x2_ASAP7_75t_R c4832(
.A(net2962),
.B(net4743),
.Y(net4875)
);

CKINVDCx12_ASAP7_75t_R c4833(
.A(net4712),
.Y(net4876)
);

XOR2xp5_ASAP7_75t_R c4834(
.A(net245),
.B(net4826),
.Y(net4877)
);

AND2x2_ASAP7_75t_R c4835(
.A(net3983),
.B(net2942),
.Y(net4878)
);

AND2x4_ASAP7_75t_R c4836(
.A(net4857),
.B(net4742),
.Y(net4879)
);

AND2x6_ASAP7_75t_R c4837(
.A(net4878),
.B(net4802),
.Y(net4880)
);

HAxp5_ASAP7_75t_R c4838(
.A(net4826),
.B(net2842),
.CON(net4881)
);

FAx1_ASAP7_75t_R c4839(
.A(net4864),
.B(net3922),
.CI(net4875),
.SN(net4882)
);

CKINVDCx14_ASAP7_75t_R c4840(
.A(net4844),
.Y(net4883)
);

NAND2x1_ASAP7_75t_R c4841(
.A(net4879),
.B(net4875),
.Y(net4884)
);

NAND2x1p5_ASAP7_75t_R c4842(
.A(net4866),
.B(net3772),
.Y(net4885)
);

NAND2x2_ASAP7_75t_R c4843(
.A(net4884),
.B(net3878),
.Y(net4886)
);

NAND2xp33_ASAP7_75t_R c4844(
.A(net2983),
.B(net3782),
.Y(net4887)
);

NAND2xp5_ASAP7_75t_R c4845(
.A(net3760),
.B(net4789),
.Y(net4888)
);

NAND2xp67_ASAP7_75t_R c4846(
.A(net4880),
.B(net2034),
.Y(net4889)
);

MAJIxp5_ASAP7_75t_R c4847(
.A(net4859),
.B(net3977),
.C(net4875),
.Y(net4890)
);

CKINVDCx16_ASAP7_75t_R c4848(
.A(net10569),
.Y(net4891)
);

MAJx2_ASAP7_75t_R c4849(
.A(net3087),
.B(net4880),
.C(net3079),
.Y(net4892)
);

MAJx3_ASAP7_75t_R c4850(
.A(net4813),
.B(net3995),
.C(net4875),
.Y(net4893)
);

NOR2x1_ASAP7_75t_R c4851(
.A(net4869),
.B(net4843),
.Y(net4894)
);

NAND3x1_ASAP7_75t_R c4852(
.A(net4881),
.B(net4644),
.C(net4858),
.Y(net4895)
);

CKINVDCx20_ASAP7_75t_R c4853(
.A(net10066),
.Y(net4896)
);

NOR2x1p5_ASAP7_75t_R c4854(
.A(net4859),
.B(net10036),
.Y(net4897)
);

CKINVDCx5p33_ASAP7_75t_R c4855(
.A(net10024),
.Y(net4898)
);

NAND3x2_ASAP7_75t_R c4856(
.B(net4894),
.C(net4891),
.A(net3952),
.Y(net4899)
);

NAND3xp33_ASAP7_75t_R c4857(
.A(net4003),
.B(net4895),
.C(net4799),
.Y(net4900)
);

NOR2x2_ASAP7_75t_R c4858(
.A(net3995),
.B(net4874),
.Y(net4901)
);

NOR2xp33_ASAP7_75t_R c4859(
.A(net4891),
.B(net9977),
.Y(net4902)
);

NOR2xp67_ASAP7_75t_R c4860(
.A(net4901),
.B(net4887),
.Y(net4903)
);

OR2x2_ASAP7_75t_R c4861(
.A(net3895),
.B(net4840),
.Y(net4904)
);

OR2x4_ASAP7_75t_R c4862(
.A(net3710),
.B(net4894),
.Y(net4905)
);

OR2x6_ASAP7_75t_R c4863(
.A(net4826),
.B(net10190),
.Y(net4906)
);

CKINVDCx6p67_ASAP7_75t_R c4864(
.A(net10085),
.Y(net4907)
);

CKINVDCx8_ASAP7_75t_R c4865(
.A(net10345),
.Y(net4908)
);

NOR3x1_ASAP7_75t_R c4866(
.A(net4861),
.B(net4897),
.C(net4893),
.Y(net4909)
);

A2O1A1O1Ixp25_ASAP7_75t_R c4867(
.A1(net4888),
.A2(net4813),
.B(net3989),
.C(net4875),
.D(net4858),
.Y(net4910)
);

CKINVDCx9p33_ASAP7_75t_R c4868(
.A(net10383),
.Y(net4911)
);

XNOR2x1_ASAP7_75t_R c4869(
.B(net3864),
.A(net2045),
.Y(net4912)
);

NOR3x2_ASAP7_75t_R c4870(
.B(net4907),
.C(net4895),
.A(net4844),
.Y(net4913)
);

XNOR2x2_ASAP7_75t_R c4871(
.A(net4769),
.B(net4906),
.Y(net4914)
);

XNOR2xp5_ASAP7_75t_R c4872(
.A(net4876),
.B(net4866),
.Y(net4915)
);

XOR2x1_ASAP7_75t_R c4873(
.A(net4743),
.B(net4857),
.Y(net4916)
);

NAND4xp25_ASAP7_75t_R c4874(
.A(net4873),
.B(net4906),
.C(net4904),
.D(net4905),
.Y(net4917)
);

XOR2x2_ASAP7_75t_R c4875(
.A(net4894),
.B(net4896),
.Y(net4918)
);

NOR3xp33_ASAP7_75t_R c4876(
.A(net4916),
.B(net4893),
.C(net3990),
.Y(net4919)
);

HB1xp67_ASAP7_75t_R c4877(
.A(net10561),
.Y(net4920)
);

XOR2xp5_ASAP7_75t_R c4878(
.A(net4902),
.B(net4874),
.Y(net4921)
);

AND2x2_ASAP7_75t_R c4879(
.A(net4828),
.B(net4887),
.Y(net4922)
);

AND2x4_ASAP7_75t_R c4880(
.A(net4866),
.B(net10048),
.Y(net4923)
);

HB2xp67_ASAP7_75t_R c4881(
.A(net10399),
.Y(net4924)
);

OA21x2_ASAP7_75t_R c4882(
.A1(net4896),
.A2(net4769),
.B(net4923),
.Y(net4925)
);

OAI21x1_ASAP7_75t_R c4883(
.A1(net4883),
.A2(net4887),
.B(net4915),
.Y(net4926)
);

NAND4xp75_ASAP7_75t_R c4884(
.A(net4921),
.B(net3938),
.C(net4875),
.D(net10223),
.Y(net4927)
);

AND2x6_ASAP7_75t_R c4885(
.A(net4904),
.B(net4914),
.Y(net4928)
);

OAI21xp33_ASAP7_75t_R c4886(
.A1(net4871),
.A2(net4901),
.B(net4868),
.Y(net4929)
);

HAxp5_ASAP7_75t_R c4887(
.A(net4923),
.B(net9876),
.CON(net4931),
.SN(net4930)
);

NAND2x1_ASAP7_75t_R c4888(
.A(net4791),
.B(net4894),
.Y(net4932)
);

HB3xp67_ASAP7_75t_R c4889(
.A(net10345),
.Y(net4933)
);

OAI21xp5_ASAP7_75t_R c4890(
.A1(net4898),
.A2(net4933),
.B(net4925),
.Y(net4934)
);

NOR4xp25_ASAP7_75t_R c4891(
.A(net3970),
.B(net4933),
.C(net3977),
.D(net10091),
.Y(net4935)
);

NOR4xp75_ASAP7_75t_R c4892(
.A(net4932),
.B(net4887),
.C(net4865),
.D(net4789),
.Y(net4936)
);

O2A1O1Ixp33_ASAP7_75t_R c4893(
.A1(net4913),
.A2(net4868),
.B(net4001),
.C(net4826),
.Y(net4937)
);

OR3x1_ASAP7_75t_R c4894(
.A(net4915),
.B(net4920),
.C(net10085),
.Y(net4938)
);

OR3x2_ASAP7_75t_R c4895(
.A(net4789),
.B(net4609),
.C(net4925),
.Y(net4939)
);

OR3x4_ASAP7_75t_R c4896(
.A(net4928),
.B(net4932),
.C(net4923),
.Y(net4940)
);

HB4xp67_ASAP7_75t_R c4897(
.A(net9777),
.Y(net4941)
);

NAND2x1p5_ASAP7_75t_R c4898(
.A(net4802),
.B(net3150),
.Y(net4942)
);

INVx11_ASAP7_75t_R c4899(
.A(net9219),
.Y(net4943)
);

INVx13_ASAP7_75t_R c4900(
.A(net10253),
.Y(net4944)
);

INVx1_ASAP7_75t_R c4901(
.A(net9102),
.Y(net4945)
);

NAND2x2_ASAP7_75t_R c4902(
.A(net3169),
.B(net4785),
.Y(net4946)
);

INVx2_ASAP7_75t_R c4903(
.A(net4014),
.Y(net4947)
);

ICGx2_ASAP7_75t_R c4904(
.ENA(net4062),
.SE(net4891),
.CLK(clk),
.GCLK(net4948)
);

ICGx2p67DC_ASAP7_75t_R c4905(
.ENA(net4926),
.SE(net3872),
.CLK(clk),
.GCLK(net4949)
);

INVx3_ASAP7_75t_R c4906(
.A(net10363),
.Y(net4950)
);

NAND2xp33_ASAP7_75t_R c4907(
.A(net3708),
.B(net10253),
.Y(net4951)
);

INVx4_ASAP7_75t_R c4908(
.A(net10019),
.Y(net4952)
);

INVx5_ASAP7_75t_R c4909(
.A(net4763),
.Y(net4953)
);

NAND2xp5_ASAP7_75t_R c4910(
.A(net4912),
.B(net10223),
.Y(net4954)
);

NAND2xp67_ASAP7_75t_R c4911(
.A(net1256),
.B(net4763),
.Y(net4955)
);

INVx6_ASAP7_75t_R c4912(
.A(net4785),
.Y(net4956)
);

NOR2x1_ASAP7_75t_R c4913(
.A(net4900),
.B(net4895),
.Y(net4957)
);

NOR2x1p5_ASAP7_75t_R c4914(
.A(net4956),
.B(net2779),
.Y(net4958)
);

NOR2x2_ASAP7_75t_R c4915(
.A(net4918),
.B(net4033),
.Y(net4959)
);

SDFLx4_ASAP7_75t_R c4916(
.D(net4952),
.SE(net4062),
.SI(net4059),
.CLK(clk),
.QN(net4960)
);

NOR2xp33_ASAP7_75t_R c4917(
.A(net3938),
.B(net4944),
.Y(net4961)
);

NOR2xp67_ASAP7_75t_R c4918(
.A(net4706),
.B(net3104),
.Y(net4962)
);

OR2x2_ASAP7_75t_R c4919(
.A(net3104),
.B(net4962),
.Y(net4963)
);

OR2x4_ASAP7_75t_R c4920(
.A(net4033),
.B(net4952),
.Y(net4964)
);

OR2x6_ASAP7_75t_R c4921(
.A(net3150),
.B(net245),
.Y(net4965)
);

INVx8_ASAP7_75t_R c4922(
.A(net10530),
.Y(net4966)
);

XNOR2x1_ASAP7_75t_R c4923(
.B(net4059),
.A(net4957),
.Y(net4967)
);

XNOR2x2_ASAP7_75t_R c4924(
.A(net4885),
.B(net4963),
.Y(net4968)
);

XNOR2xp5_ASAP7_75t_R c4925(
.A(net4949),
.B(net4948),
.Y(net4969)
);

INVxp33_ASAP7_75t_R c4926(
.A(net4969),
.Y(net4970)
);

XOR2x1_ASAP7_75t_R c4927(
.A(net4915),
.B(net4952),
.Y(net4971)
);

XOR2x2_ASAP7_75t_R c4928(
.A(net3142),
.B(net1861),
.Y(net4972)
);

INVxp67_ASAP7_75t_R c4929(
.A(net3067),
.Y(net4973)
);

XOR2xp5_ASAP7_75t_R c4930(
.A(net4644),
.B(net4863),
.Y(net4974)
);

AND3x1_ASAP7_75t_R c4931(
.A(net4780),
.B(net4950),
.C(net4948),
.Y(net4975)
);

BUFx10_ASAP7_75t_R c4932(
.A(net2942),
.Y(net4976)
);

BUFx12_ASAP7_75t_R c4933(
.A(net10573),
.Y(net4977)
);

BUFx12f_ASAP7_75t_R c4934(
.A(net10409),
.Y(net4978)
);

AND3x2_ASAP7_75t_R c4935(
.A(net4912),
.B(net2180),
.C(net4926),
.Y(net4979)
);

AND2x2_ASAP7_75t_R c4936(
.A(net2164),
.B(net4949),
.Y(net4980)
);

AND2x4_ASAP7_75t_R c4937(
.A(net4948),
.B(net4954),
.Y(net4981)
);

BUFx16f_ASAP7_75t_R c4938(
.A(net9102),
.Y(net4982)
);

BUFx24_ASAP7_75t_R c4939(
.A(net10520),
.Y(net4983)
);

DFFASRHQNx1_ASAP7_75t_R c4940(
.D(net4961),
.RESETN(net4982),
.SETN(net4936),
.CLK(clk),
.QN(net4984)
);

AND3x4_ASAP7_75t_R c4941(
.A(net4874),
.B(net4964),
.C(net4950),
.Y(net4985)
);

BUFx2_ASAP7_75t_R c4942(
.A(net4017),
.Y(net4986)
);

AND2x6_ASAP7_75t_R c4943(
.A(net4895),
.B(net4970),
.Y(net4987)
);

HAxp5_ASAP7_75t_R c4944(
.A(net4945),
.B(net4971),
.CON(net4988)
);

NAND2x1_ASAP7_75t_R c4945(
.A(net4982),
.B(net4944),
.Y(net4989)
);

NAND2x1p5_ASAP7_75t_R c4946(
.A(net4051),
.B(net4959),
.Y(net4990)
);

BUFx3_ASAP7_75t_R c4947(
.A(net10067),
.Y(net4991)
);

NAND2x2_ASAP7_75t_R c4948(
.A(net4988),
.B(net1190),
.Y(net4992)
);

NAND2xp33_ASAP7_75t_R c4949(
.A(net4984),
.B(net4963),
.Y(net4993)
);

BUFx4_ASAP7_75t_R c4950(
.A(net10475),
.Y(net4994)
);

AND5x1_ASAP7_75t_R c4951(
.A(net4976),
.B(net4994),
.C(net4983),
.D(net4961),
.E(net3086),
.Y(net4995)
);

AO21x1_ASAP7_75t_R c4952(
.A1(net4966),
.A2(net4897),
.B(net4978),
.Y(net4996)
);

OAI321xp33_ASAP7_75t_R c4953(
.A1(net4038),
.A2(net3142),
.A3(net3977),
.B1(net4027),
.B2(net4957),
.C(net4962),
.Y(net4997)
);

AO21x2_ASAP7_75t_R c4954(
.A1(net4958),
.A2(net4964),
.B(net2180),
.Y(net4998)
);

NAND2xp5_ASAP7_75t_R c4955(
.A(net1190),
.B(net4993),
.Y(net4999)
);

NAND2xp67_ASAP7_75t_R c4956(
.A(net4990),
.B(net4982),
.Y(net5000)
);

NOR2x1_ASAP7_75t_R c4957(
.A(net4993),
.B(net9946),
.Y(net5001)
);

NOR2x1p5_ASAP7_75t_R c4958(
.A(net4980),
.B(net4959),
.Y(net5002)
);

AOI21x1_ASAP7_75t_R c4959(
.A1(net4983),
.A2(net4049),
.B(net4994),
.Y(net5003)
);

AOI21xp33_ASAP7_75t_R c4960(
.A1(net4987),
.A2(net3067),
.B(net10255),
.Y(net5004)
);

BUFx4f_ASAP7_75t_R c4961(
.A(net10532),
.Y(net5005)
);

NOR2x2_ASAP7_75t_R c4962(
.A(net4961),
.B(net9670),
.Y(net5006)
);

O2A1O1Ixp5_ASAP7_75t_R c4963(
.A1(net4995),
.A2(net3142),
.B(net5005),
.C(net4027),
.Y(net5007)
);

AOI21xp5_ASAP7_75t_R c4964(
.A1(net4999),
.A2(net4961),
.B(net10168),
.Y(net5008)
);

FAx1_ASAP7_75t_R c4965(
.A(net4860),
.B(net4984),
.CI(net10255),
.SN(net5010),
.CON(net5009)
);

MAJIxp5_ASAP7_75t_R c4966(
.A(net5009),
.B(net2180),
.C(net9788),
.Y(net5011)
);

NOR2xp33_ASAP7_75t_R c4967(
.A(net4991),
.B(net5005),
.Y(net5012)
);

MAJx2_ASAP7_75t_R c4968(
.A(net4986),
.B(net4984),
.C(net4961),
.Y(net5013)
);

NOR2xp67_ASAP7_75t_R c4969(
.A(net4950),
.B(net10120),
.Y(net5014)
);

BUFx5_ASAP7_75t_R c4970(
.A(net10543),
.Y(net5015)
);

OR2x2_ASAP7_75t_R c4971(
.A(net4993),
.B(net5015),
.Y(net5016)
);

SDFHx1_ASAP7_75t_R c4972(
.D(net4936),
.SE(net4995),
.SI(net10224),
.CLK(clk),
.QN(net5017)
);

MAJx3_ASAP7_75t_R c4973(
.A(net4047),
.B(net5017),
.C(net9670),
.Y(net5018)
);

OAI33xp33_ASAP7_75t_R c4974(
.A1(net4994),
.A2(net2164),
.A3(net5017),
.B1(net4962),
.B2(net3772),
.B3(net10120),
.Y(net5019)
);

NAND3x1_ASAP7_75t_R c4975(
.A(net5017),
.B(net5019),
.C(net5016),
.Y(net5020)
);

OR2x4_ASAP7_75t_R c4976(
.A(net4965),
.B(net3132),
.Y(net5021)
);

NAND3x2_ASAP7_75t_R c4977(
.B(net5014),
.C(net5017),
.A(net10168),
.Y(net5022)
);

AO222x2_ASAP7_75t_R c4978(
.A1(net3132),
.A2(net5012),
.B1(net5017),
.B2(net4827),
.C1(net4059),
.C2(net10255),
.Y(net5023)
);

NAND3xp33_ASAP7_75t_R c4979(
.A(net5019),
.B(net5018),
.C(net3877),
.Y(net5024)
);

BUFx6f_ASAP7_75t_R c4980(
.A(net5021),
.Y(net5025)
);

OR2x6_ASAP7_75t_R c4981(
.A(net4989),
.B(net4992),
.Y(net5026)
);

BUFx8_ASAP7_75t_R c4982(
.A(net2214),
.Y(net5027)
);

XNOR2x1_ASAP7_75t_R c4983(
.B(net4977),
.A(net3246),
.Y(net5028)
);

XNOR2x2_ASAP7_75t_R c4984(
.A(net4045),
.B(net4166),
.Y(net5029)
);

SDFHx2_ASAP7_75t_R c4985(
.D(net4137),
.SE(net5028),
.SI(net5002),
.CLK(clk),
.QN(net5030)
);

XNOR2xp5_ASAP7_75t_R c4986(
.A(net5018),
.B(net4116),
.Y(net5031)
);

CKINVDCx10_ASAP7_75t_R c4987(
.A(net4992),
.Y(net5032)
);

CKINVDCx11_ASAP7_75t_R c4988(
.A(net9151),
.Y(net5033)
);

XOR2x1_ASAP7_75t_R c4989(
.A(net4040),
.B(net4109),
.Y(net5034)
);

CKINVDCx12_ASAP7_75t_R c4990(
.A(net9151),
.Y(net5035)
);

NOR3x1_ASAP7_75t_R c4991(
.A(net5027),
.B(net4049),
.C(net4027),
.Y(net5036)
);

NOR3x2_ASAP7_75t_R c4992(
.B(net5031),
.C(net5012),
.A(net4148),
.Y(net5037)
);

CKINVDCx14_ASAP7_75t_R c4993(
.A(net10110),
.Y(net5038)
);

CKINVDCx16_ASAP7_75t_R c4994(
.A(net9208),
.Y(net5039)
);

XOR2x2_ASAP7_75t_R c4995(
.A(net5037),
.B(net4925),
.Y(net5040)
);

CKINVDCx20_ASAP7_75t_R c4996(
.A(net1238),
.Y(net5041)
);

NOR3xp33_ASAP7_75t_R c4997(
.A(net3246),
.B(net5025),
.C(net5023),
.Y(net5042)
);

XOR2xp5_ASAP7_75t_R c4998(
.A(net4056),
.B(net1348),
.Y(net5043)
);

AND2x2_ASAP7_75t_R c4999(
.A(net5029),
.B(net4173),
.Y(net5044)
);

AND2x4_ASAP7_75t_R c5000(
.A(net4943),
.B(net5033),
.Y(net5045)
);

CKINVDCx5p33_ASAP7_75t_R c5001(
.A(net5041),
.Y(net5046)
);

AND2x6_ASAP7_75t_R c5002(
.A(net4154),
.B(net4116),
.Y(net5047)
);

CKINVDCx6p67_ASAP7_75t_R c5003(
.A(net9219),
.Y(net5048)
);

CKINVDCx8_ASAP7_75t_R c5004(
.A(net5046),
.Y(net5049)
);

HAxp5_ASAP7_75t_R c5005(
.A(net4080),
.B(net5016),
.CON(net5050)
);

CKINVDCx9p33_ASAP7_75t_R c5006(
.A(net10489),
.Y(net5051)
);

HB1xp67_ASAP7_75t_R c5007(
.A(net5048),
.Y(net5052)
);

OA21x2_ASAP7_75t_R c5008(
.A1(net4128),
.A2(net5046),
.B(net10138),
.Y(net5053)
);

NAND2x1_ASAP7_75t_R c5009(
.A(net4992),
.B(net10138),
.Y(net5054)
);

OAI21x1_ASAP7_75t_R c5010(
.A1(net5025),
.A2(net5035),
.B(net3246),
.Y(net5055)
);

OAI21xp33_ASAP7_75t_R c5011(
.A1(net5040),
.A2(net5039),
.B(net4148),
.Y(net5056)
);

NAND2x1p5_ASAP7_75t_R c5012(
.A(net4818),
.B(net4019),
.Y(net5057)
);

SDFHx3_ASAP7_75t_R c5013(
.D(net4019),
.SE(net5018),
.SI(net5056),
.CLK(clk),
.QN(net5058)
);

HB2xp67_ASAP7_75t_R c5014(
.A(net4891),
.Y(net5059)
);

HB3xp67_ASAP7_75t_R c5015(
.A(net4155),
.Y(net5060)
);

NAND2x2_ASAP7_75t_R c5016(
.A(net4890),
.B(net5057),
.Y(net5061)
);

NAND2xp33_ASAP7_75t_R c5017(
.A(net3232),
.B(net4978),
.Y(net5062)
);

HB4xp67_ASAP7_75t_R c5018(
.A(net9227),
.Y(net5063)
);

NAND2xp5_ASAP7_75t_R c5019(
.A(net5052),
.B(net4045),
.Y(net5064)
);

NAND2xp67_ASAP7_75t_R c5020(
.A(net5049),
.B(net5059),
.Y(net5065)
);

INVx11_ASAP7_75t_R c5021(
.A(net10517),
.Y(net5066)
);

NOR2x1_ASAP7_75t_R c5022(
.A(net5054),
.B(net10124),
.Y(net5067)
);

INVx13_ASAP7_75t_R c5023(
.A(net10544),
.Y(net5068)
);

OAI21xp5_ASAP7_75t_R c5024(
.A1(net5060),
.A2(net5057),
.B(net5065),
.Y(net5069)
);

OR3x1_ASAP7_75t_R c5025(
.A(net5051),
.B(net4116),
.C(net4047),
.Y(net5070)
);

INVx1_ASAP7_75t_R c5026(
.A(net10465),
.Y(net5071)
);

INVx2_ASAP7_75t_R c5027(
.A(net10529),
.Y(net5072)
);

OR3x2_ASAP7_75t_R c5028(
.A(net5065),
.B(net5054),
.C(net5018),
.Y(net5073)
);

AND5x2_ASAP7_75t_R c5029(
.A(net5056),
.B(net4121),
.C(net5001),
.D(net5035),
.E(net5033),
.Y(net5074)
);

OR3x4_ASAP7_75t_R c5030(
.A(net5053),
.B(net5057),
.C(net4121),
.Y(net5075)
);

NOR2x1p5_ASAP7_75t_R c5031(
.A(net3227),
.B(net4148),
.Y(net5076)
);

ICGx3_ASAP7_75t_R c5032(
.ENA(net2292),
.SE(net3049),
.CLK(clk),
.GCLK(net5077)
);

INVx3_ASAP7_75t_R c5033(
.A(net10110),
.Y(net5078)
);

NOR2x2_ASAP7_75t_R c5034(
.A(net5078),
.B(net4931),
.Y(net5079)
);

AND3x1_ASAP7_75t_R c5035(
.A(net4117),
.B(net5079),
.C(net4891),
.Y(net5080)
);

NOR2xp33_ASAP7_75t_R c5036(
.A(net5063),
.B(net3227),
.Y(net5081)
);

NOR2xp67_ASAP7_75t_R c5037(
.A(net4176),
.B(net5065),
.Y(net5082)
);

OR2x2_ASAP7_75t_R c5038(
.A(net5042),
.B(net4981),
.Y(net5083)
);

ICGx4DC_ASAP7_75t_R c5039(
.ENA(net5028),
.SE(net5037),
.CLK(clk),
.GCLK(net5084)
);

AND3x2_ASAP7_75t_R c5040(
.A(net4047),
.B(net4173),
.C(net10084),
.Y(net5085)
);

OR2x4_ASAP7_75t_R c5041(
.A(net4147),
.B(net5015),
.Y(net5086)
);

AND3x4_ASAP7_75t_R c5042(
.A(net5084),
.B(net5036),
.C(net9910),
.Y(net5087)
);

OR2x6_ASAP7_75t_R c5043(
.A(net5084),
.B(net4749),
.Y(net5088)
);

XNOR2x1_ASAP7_75t_R c5044(
.B(net5079),
.A(net452),
.Y(net5089)
);

AO21x1_ASAP7_75t_R c5045(
.A1(net5086),
.A2(net5085),
.B(net4818),
.Y(net5090)
);

XNOR2x2_ASAP7_75t_R c5046(
.A(net5088),
.B(net5077),
.Y(net5091)
);

XNOR2xp5_ASAP7_75t_R c5047(
.A(net4180),
.B(net5077),
.Y(net5092)
);

XOR2x1_ASAP7_75t_R c5048(
.A(net5045),
.B(net5088),
.Y(net5093)
);

INVx4_ASAP7_75t_R c5049(
.A(net10489),
.Y(net5094)
);

INVx5_ASAP7_75t_R c5050(
.A(net10166),
.Y(net5095)
);

SDFHx4_ASAP7_75t_R c5051(
.D(net5089),
.SE(net5088),
.SI(net5062),
.CLK(clk),
.QN(net5096)
);

AO221x1_ASAP7_75t_R c5052(
.A1(net4934),
.A2(net5096),
.B1(net2292),
.B2(net5072),
.C(net5047),
.Y(net5097)
);

AO221x2_ASAP7_75t_R c5053(
.A1(net4026),
.A2(net4897),
.B1(net4139),
.B2(net5072),
.C(net3086),
.Y(net5098)
);

AO21x2_ASAP7_75t_R c5054(
.A1(net5034),
.A2(net5065),
.B(net5088),
.Y(net5099)
);

XOR2x2_ASAP7_75t_R c5055(
.A(net5068),
.B(net5093),
.Y(net5100)
);

AO32x1_ASAP7_75t_R c5056(
.A1(net5090),
.A2(net5100),
.A3(net5097),
.B1(net5059),
.B2(net5072),
.Y(net5101)
);

XOR2xp5_ASAP7_75t_R c5057(
.A(net5038),
.B(net9775),
.Y(net5102)
);

AOI21x1_ASAP7_75t_R c5058(
.A1(net5102),
.A2(net5100),
.B(net5072),
.Y(net5103)
);

AOI21xp33_ASAP7_75t_R c5059(
.A1(net5066),
.A2(net5103),
.B(net5078),
.Y(net5104)
);

AO33x2_ASAP7_75t_R c5060(
.A1(net5071),
.A2(net5104),
.A3(net5064),
.B1(net5084),
.B2(net5058),
.B3(net5077),
.Y(net5105)
);

AND2x2_ASAP7_75t_R c5061(
.A(net5103),
.B(net5104),
.Y(net5106)
);

AOI222xp33_ASAP7_75t_R c5062(
.A1(net5106),
.A2(net5103),
.B1(net5104),
.B2(net4110),
.C1(net5077),
.C2(net9859),
.Y(net5107)
);

AND2x4_ASAP7_75t_R c5063(
.A(net4109),
.B(net4198),
.Y(net5108)
);

AND2x6_ASAP7_75t_R c5064(
.A(net5058),
.B(net10101),
.Y(net5109)
);

INVx6_ASAP7_75t_R c5065(
.A(net907),
.Y(net5110)
);

INVx8_ASAP7_75t_R c5066(
.A(net4652),
.Y(net5111)
);

INVxp33_ASAP7_75t_R c5067(
.A(net2364),
.Y(net5112)
);

HAxp5_ASAP7_75t_R c5068(
.A(net4251),
.B(net5091),
.CON(net5113)
);

INVxp67_ASAP7_75t_R c5069(
.A(net4862),
.Y(net5114)
);

NAND2x1_ASAP7_75t_R c5070(
.A(net4027),
.B(net4247),
.Y(net5115)
);

BUFx10_ASAP7_75t_R c5071(
.A(net4049),
.Y(net5116)
);

BUFx12_ASAP7_75t_R c5072(
.A(net4722),
.Y(net5117)
);

BUFx12f_ASAP7_75t_R c5073(
.A(net9191),
.Y(net5118)
);

NAND2x1p5_ASAP7_75t_R c5074(
.A(net5057),
.B(net4247),
.Y(net5119)
);

NAND2x2_ASAP7_75t_R c5075(
.A(net4217),
.B(net4049),
.Y(net5120)
);

BUFx16f_ASAP7_75t_R c5076(
.A(net9191),
.Y(net5121)
);

BUFx24_ASAP7_75t_R c5077(
.A(net4247),
.Y(net5122)
);

BUFx2_ASAP7_75t_R c5078(
.A(net4944),
.Y(net5123)
);

BUFx3_ASAP7_75t_R c5079(
.A(net10157),
.Y(net5124)
);

BUFx4_ASAP7_75t_R c5080(
.A(net4182),
.Y(net5125)
);

BUFx4f_ASAP7_75t_R c5081(
.A(net5064),
.Y(net5126)
);

BUFx5_ASAP7_75t_R c5082(
.A(net5096),
.Y(net5127)
);

BUFx6f_ASAP7_75t_R c5083(
.A(net3257),
.Y(net5128)
);

AOI21xp5_ASAP7_75t_R c5084(
.A1(net5122),
.A2(net531),
.B(net5128),
.Y(net5129)
);

BUFx8_ASAP7_75t_R c5085(
.A(net5108),
.Y(net5130)
);

NAND2xp33_ASAP7_75t_R c5086(
.A(net5091),
.B(net4243),
.Y(net5131)
);

CKINVDCx10_ASAP7_75t_R c5087(
.A(net9204),
.Y(net5132)
);

CKINVDCx11_ASAP7_75t_R c5088(
.A(net4198),
.Y(net5133)
);

CKINVDCx12_ASAP7_75t_R c5089(
.A(net4974),
.Y(net5134)
);

SDFLx1_ASAP7_75t_R c5090(
.D(net5117),
.SE(net5070),
.SI(net5002),
.CLK(clk),
.QN(net5135)
);

CKINVDCx14_ASAP7_75t_R c5091(
.A(net9955),
.Y(net5136)
);

CKINVDCx16_ASAP7_75t_R c5092(
.A(net5119),
.Y(net5137)
);

CKINVDCx20_ASAP7_75t_R c5093(
.A(net10456),
.Y(net5138)
);

AO32x2_ASAP7_75t_R c5094(
.A1(net4925),
.A2(net3267),
.A3(net5135),
.B1(net4897),
.B2(net5111),
.Y(net5139)
);

CKINVDCx5p33_ASAP7_75t_R c5095(
.A(net4219),
.Y(net5140)
);

NAND2xp5_ASAP7_75t_R c5096(
.A(net4179),
.B(net5138),
.Y(net5141)
);

OA211x2_ASAP7_75t_R c5097(
.A1(net5137),
.A2(net5128),
.B(net5057),
.C(net2400),
.Y(net5142)
);

NAND2xp67_ASAP7_75t_R c5098(
.A(net4113),
.B(net4217),
.Y(net5143)
);

OA22x2_ASAP7_75t_R c5099(
.A1(net3298),
.A2(net5096),
.B1(net4246),
.B2(net5111),
.Y(net5144)
);

NOR2x1_ASAP7_75t_R c5100(
.A(net5136),
.B(net4219),
.Y(net5145)
);

NOR2x1p5_ASAP7_75t_R c5101(
.A(net5070),
.B(net4195),
.Y(net5146)
);

CKINVDCx6p67_ASAP7_75t_R c5102(
.A(net9229),
.Y(net5147)
);

FAx1_ASAP7_75t_R c5103(
.A(net5132),
.B(net4113),
.CI(net4049),
.SN(net5149),
.CON(net5148)
);

NOR2x2_ASAP7_75t_R c5104(
.A(net1424),
.B(net5124),
.Y(net5150)
);

CKINVDCx8_ASAP7_75t_R c5105(
.A(net5095),
.Y(net5151)
);

ICGx4_ASAP7_75t_R c5106(
.ENA(net5151),
.SE(net2381),
.CLK(clk),
.GCLK(net5152)
);

NOR2xp33_ASAP7_75t_R c5107(
.A(net5131),
.B(net5148),
.Y(net5153)
);

NOR2xp67_ASAP7_75t_R c5108(
.A(net5120),
.B(net4264),
.Y(net5154)
);

OR2x2_ASAP7_75t_R c5109(
.A(net4218),
.B(net5154),
.Y(net5155)
);

CKINVDCx9p33_ASAP7_75t_R c5110(
.A(net10484),
.Y(net5156)
);

OR2x4_ASAP7_75t_R c5111(
.A(net5109),
.B(net5072),
.Y(net5157)
);

MAJIxp5_ASAP7_75t_R c5112(
.A(net5139),
.B(net5156),
.C(net5058),
.Y(net5158)
);

OR2x6_ASAP7_75t_R c5113(
.A(net5092),
.B(net4219),
.Y(net5159)
);

HB1xp67_ASAP7_75t_R c5114(
.A(net10548),
.Y(net5160)
);

OA31x2_ASAP7_75t_R c5115(
.A1(net5149),
.A2(net5058),
.A3(net5154),
.B1(net5111),
.Y(net5161)
);

XNOR2x1_ASAP7_75t_R c5116(
.B(net5158),
.A(net5030),
.Y(net5162)
);

XNOR2x2_ASAP7_75t_R c5117(
.A(net5133),
.B(net5143),
.Y(net5163)
);

XNOR2xp5_ASAP7_75t_R c5118(
.A(net5126),
.B(net4134),
.Y(net5164)
);

HB2xp67_ASAP7_75t_R c5119(
.A(net10445),
.Y(net5165)
);

XOR2x1_ASAP7_75t_R c5120(
.A(net5160),
.B(net5164),
.Y(net5166)
);

HB3xp67_ASAP7_75t_R c5121(
.A(net9672),
.Y(net5167)
);

MAJx2_ASAP7_75t_R c5122(
.A(net3218),
.B(net5156),
.C(net10257),
.Y(net5168)
);

ICGx5_ASAP7_75t_R c5123(
.ENA(net5166),
.SE(net5154),
.CLK(clk),
.GCLK(net5169)
);

HB4xp67_ASAP7_75t_R c5124(
.A(net5169),
.Y(net5170)
);

INVx11_ASAP7_75t_R c5125(
.A(net10257),
.Y(net5171)
);

XOR2x2_ASAP7_75t_R c5126(
.A(net5156),
.B(net4027),
.Y(net5172)
);

XOR2xp5_ASAP7_75t_R c5127(
.A(net5114),
.B(net5030),
.Y(net5173)
);

OAI211xp5_ASAP7_75t_R c5128(
.A1(net5016),
.A2(net4113),
.B(net5156),
.C(net5096),
.Y(net5174)
);

MAJx3_ASAP7_75t_R c5129(
.A(net5146),
.B(net4045),
.C(net5169),
.Y(net5175)
);

AND2x2_ASAP7_75t_R c5130(
.A(net5175),
.B(net5167),
.Y(net5176)
);

OAI22x1_ASAP7_75t_R c5131(
.A1(net4906),
.A2(net2390),
.B1(net5165),
.B2(net4962),
.Y(net5177)
);

AND2x4_ASAP7_75t_R c5132(
.A(net5116),
.B(net5172),
.Y(net5178)
);

INVx13_ASAP7_75t_R c5133(
.A(net10536),
.Y(net5179)
);

NAND3x1_ASAP7_75t_R c5134(
.A(net4134),
.B(net5175),
.C(net5172),
.Y(net5180)
);

AND2x6_ASAP7_75t_R c5135(
.A(net5179),
.B(net5170),
.Y(net5181)
);

SDFLx2_ASAP7_75t_R c5136(
.D(net5178),
.SE(net5035),
.SI(net9672),
.CLK(clk),
.QN(net5182)
);

HAxp5_ASAP7_75t_R c5137(
.A(net5169),
.B(net9917),
.CON(net5183)
);

ICGx5p33DC_ASAP7_75t_R c5138(
.ENA(net5180),
.SE(net10256),
.CLK(clk),
.GCLK(net5184)
);

ICGx6p67DC_ASAP7_75t_R c5139(
.ENA(net5142),
.SE(net4262),
.CLK(clk),
.GCLK(net5185)
);

NAND3x2_ASAP7_75t_R c5140(
.B(net5177),
.C(net5184),
.A(net4251),
.Y(net5186)
);

INVx1_ASAP7_75t_R c5141(
.A(net10547),
.Y(net5187)
);

NAND3xp33_ASAP7_75t_R c5142(
.A(net5186),
.B(net5182),
.C(net4179),
.Y(net5188)
);

NAND2x1_ASAP7_75t_R c5143(
.A(net5183),
.B(net5182),
.Y(net5189)
);

INVx2_ASAP7_75t_R c5144(
.A(net10042),
.Y(net5190)
);

NAND2x1p5_ASAP7_75t_R c5145(
.A(net5189),
.B(net5190),
.Y(net5191)
);

INVx3_ASAP7_75t_R c5146(
.A(net5170),
.Y(net5192)
);

INVx4_ASAP7_75t_R c5147(
.A(net9145),
.Y(net5193)
);

INVx5_ASAP7_75t_R c5148(
.A(net5159),
.Y(net5194)
);

INVx6_ASAP7_75t_R c5149(
.A(net5128),
.Y(net5195)
);

INVx8_ASAP7_75t_R c5150(
.A(net10516),
.Y(net5196)
);

NAND2x2_ASAP7_75t_R c5151(
.A(net5157),
.B(net5168),
.Y(net5197)
);

NAND2xp33_ASAP7_75t_R c5152(
.A(net4344),
.B(net5129),
.Y(net5198)
);

NOR3x1_ASAP7_75t_R c5153(
.A(net2499),
.B(net4252),
.C(net10242),
.Y(net5199)
);

INVxp33_ASAP7_75t_R c5154(
.A(net9145),
.Y(net5200)
);

INVxp67_ASAP7_75t_R c5155(
.A(net4288),
.Y(net5201)
);

NAND2xp5_ASAP7_75t_R c5156(
.A(net4170),
.B(net5123),
.Y(net5202)
);

NOR3x2_ASAP7_75t_R c5157(
.B(net5196),
.C(net5035),
.A(net5187),
.Y(net5203)
);

BUFx10_ASAP7_75t_R c5158(
.A(net10061),
.Y(net5204)
);

NAND2xp67_ASAP7_75t_R c5159(
.A(net5201),
.B(net5072),
.Y(net5205)
);

BUFx12_ASAP7_75t_R c5160(
.A(net5002),
.Y(net5206)
);

BUFx12f_ASAP7_75t_R c5161(
.A(net9229),
.Y(net5207)
);

NOR2x1_ASAP7_75t_R c5162(
.A(net4347),
.B(net5077),
.Y(net5208)
);

BUFx16f_ASAP7_75t_R c5163(
.A(net5202),
.Y(net5209)
);

NOR2x1p5_ASAP7_75t_R c5164(
.A(net5150),
.B(net4308),
.Y(net5210)
);

BUFx24_ASAP7_75t_R c5165(
.A(net10502),
.Y(net5211)
);

BUFx2_ASAP7_75t_R c5166(
.A(net4243),
.Y(net5212)
);

BUFx3_ASAP7_75t_R c5167(
.A(net5208),
.Y(net5213)
);

BUFx4_ASAP7_75t_R c5168(
.A(net5204),
.Y(net5214)
);

BUFx4f_ASAP7_75t_R c5169(
.A(net3406),
.Y(net5215)
);

BUFx5_ASAP7_75t_R c5170(
.A(net10084),
.Y(net5216)
);

NOR2x2_ASAP7_75t_R c5171(
.A(net5195),
.B(net4206),
.Y(net5217)
);

NOR2xp33_ASAP7_75t_R c5172(
.A(net5216),
.B(net9735),
.Y(net5218)
);

BUFx6f_ASAP7_75t_R c5173(
.A(net10443),
.Y(net5219)
);

NOR3xp33_ASAP7_75t_R c5174(
.A(net5141),
.B(net5047),
.C(net5217),
.Y(net5220)
);

NOR2xp67_ASAP7_75t_R c5175(
.A(net5212),
.B(net3412),
.Y(net5221)
);

OR2x2_ASAP7_75t_R c5176(
.A(net5216),
.B(net5035),
.Y(net5222)
);

BUFx8_ASAP7_75t_R c5177(
.A(net3389),
.Y(net5223)
);

OR2x4_ASAP7_75t_R c5178(
.A(net5207),
.B(net4229),
.Y(net5224)
);

SDFLx3_ASAP7_75t_R c5179(
.D(net5194),
.SE(net4302),
.SI(net5200),
.CLK(clk),
.QN(net5225)
);

OR2x6_ASAP7_75t_R c5180(
.A(net5209),
.B(net5224),
.Y(net5226)
);

XNOR2x1_ASAP7_75t_R c5181(
.B(net5210),
.A(net5047),
.Y(net5227)
);

XNOR2x2_ASAP7_75t_R c5182(
.A(net5226),
.B(net5208),
.Y(net5228)
);

XNOR2xp5_ASAP7_75t_R c5183(
.A(net4206),
.B(net5208),
.Y(net5229)
);

XOR2x1_ASAP7_75t_R c5184(
.A(net2497),
.B(net5217),
.Y(net5230)
);

XOR2x2_ASAP7_75t_R c5185(
.A(net4002),
.B(net5210),
.Y(net5231)
);

XOR2xp5_ASAP7_75t_R c5186(
.A(net5214),
.B(net2452),
.Y(net5232)
);

AND2x2_ASAP7_75t_R c5187(
.A(net5203),
.B(net5167),
.Y(net5233)
);

AND2x4_ASAP7_75t_R c5188(
.A(net5231),
.B(net5225),
.Y(net5234)
);

AND2x6_ASAP7_75t_R c5189(
.A(net5205),
.B(net4272),
.Y(net5235)
);

HAxp5_ASAP7_75t_R c5190(
.A(net5199),
.B(net5072),
.CON(net5237),
.SN(net5236)
);

CKINVDCx10_ASAP7_75t_R c5191(
.A(net10361),
.Y(net5238)
);

CKINVDCx11_ASAP7_75t_R c5192(
.A(net5072),
.Y(net5239)
);

NAND2x1_ASAP7_75t_R c5193(
.A(net5190),
.B(net5224),
.Y(net5240)
);

OA21x2_ASAP7_75t_R c5194(
.A1(net5215),
.A2(net3416),
.B(net3412),
.Y(net5241)
);

CKINVDCx12_ASAP7_75t_R c5195(
.A(net10538),
.Y(net5242)
);

CKINVDCx14_ASAP7_75t_R c5196(
.A(net10137),
.Y(net5243)
);

CKINVDCx16_ASAP7_75t_R c5197(
.A(net10148),
.Y(net5244)
);

NAND2x1p5_ASAP7_75t_R c5198(
.A(net5129),
.B(net5229),
.Y(net5245)
);

CKINVDCx20_ASAP7_75t_R c5199(
.A(net4272),
.Y(net5246)
);

NAND2x2_ASAP7_75t_R c5200(
.A(net5235),
.B(net9656),
.Y(net5247)
);

NAND2xp33_ASAP7_75t_R c5201(
.A(net5244),
.B(net5192),
.Y(net5248)
);

NAND2xp5_ASAP7_75t_R c5202(
.A(net5248),
.B(net2498),
.Y(net5249)
);

OAI21x1_ASAP7_75t_R c5203(
.A1(net5233),
.A2(net5168),
.B(net5147),
.Y(net5250)
);

NAND2xp67_ASAP7_75t_R c5204(
.A(net1348),
.B(net5244),
.Y(net5251)
);

CKINVDCx5p33_ASAP7_75t_R c5205(
.A(net5035),
.Y(net5252)
);

NOR2x1_ASAP7_75t_R c5206(
.A(net4321),
.B(net1490),
.Y(net5253)
);

NOR2x1p5_ASAP7_75t_R c5207(
.A(net5206),
.B(net5216),
.Y(net5254)
);

OAI22xp33_ASAP7_75t_R c5208(
.A1(net4994),
.A2(net5238),
.B1(net5077),
.B2(net10254),
.Y(net5255)
);

NOR2x2_ASAP7_75t_R c5209(
.A(net5235),
.B(net5254),
.Y(net5256)
);

CKINVDCx6p67_ASAP7_75t_R c5210(
.A(net10135),
.Y(net5257)
);

OAI21xp33_ASAP7_75t_R c5211(
.A1(net5254),
.A2(net4257),
.B(net4229),
.Y(net5258)
);

OAI21xp5_ASAP7_75t_R c5212(
.A1(net5256),
.A2(net5242),
.B(net5257),
.Y(net5259)
);

NOR2xp33_ASAP7_75t_R c5213(
.A(net5258),
.B(net5246),
.Y(net5260)
);

NOR2xp67_ASAP7_75t_R c5214(
.A(net5243),
.B(net5260),
.Y(net5261)
);

OR2x2_ASAP7_75t_R c5215(
.A(net5123),
.B(net5254),
.Y(net5262)
);

OR3x1_ASAP7_75t_R c5216(
.A(net4305),
.B(net5223),
.C(net3406),
.Y(net5263)
);

OR2x4_ASAP7_75t_R c5217(
.A(net5224),
.B(net5201),
.Y(net5264)
);

OR3x2_ASAP7_75t_R c5218(
.A(net5218),
.B(net5210),
.C(net9835),
.Y(net5265)
);

SDFLx4_ASAP7_75t_R c5219(
.D(net5265),
.SE(net5263),
.SI(net5262),
.CLK(clk),
.QN(net5266)
);

OR2x6_ASAP7_75t_R c5220(
.A(net3941),
.B(net5231),
.Y(net5267)
);

AOI321xp33_ASAP7_75t_R c5221(
.A1(net5264),
.A2(net5242),
.A3(net5255),
.B1(net5224),
.B2(net5257),
.C(net10242),
.Y(net5268)
);

XNOR2x1_ASAP7_75t_R c5222(
.B(net5219),
.A(net5257),
.Y(net5269)
);

AOI221x1_ASAP7_75t_R c5223(
.A1(net5200),
.A2(net5221),
.B1(net5263),
.B2(net5260),
.C(net5203),
.Y(net5270)
);

XNOR2x2_ASAP7_75t_R c5224(
.A(net4252),
.B(net5265),
.Y(net5271)
);

AOI221xp5_ASAP7_75t_R c5225(
.A1(net5238),
.A2(net5167),
.B1(net5265),
.B2(net5225),
.C(net5260),
.Y(net5272)
);

AOI311xp33_ASAP7_75t_R c5226(
.A1(net5259),
.A2(net4272),
.A3(net5225),
.B(net5257),
.C(net5077),
.Y(net5273)
);

DFFASRHQNx1_ASAP7_75t_R c5227(
.D(net5271),
.RESETN(net5262),
.SETN(net10258),
.CLK(clk),
.QN(net5274)
);

SDFHx1_ASAP7_75t_R c5228(
.D(net5273),
.SE(net5240),
.SI(net4960),
.CLK(clk),
.QN(net5275)
);

XNOR2xp5_ASAP7_75t_R c5229(
.A(net4427),
.B(net5221),
.Y(net5276)
);

XOR2x1_ASAP7_75t_R c5230(
.A(net4399),
.B(net1078),
.Y(net5277)
);

CKINVDCx8_ASAP7_75t_R c5231(
.A(net9467),
.Y(out25)
);

XOR2x2_ASAP7_75t_R c5232(
.A(net5220),
.B(net2399),
.Y(net5278)
);

CKINVDCx9p33_ASAP7_75t_R c5233(
.A(net10129),
.Y(net5279)
);

OR3x4_ASAP7_75t_R c5234(
.A(net3424),
.B(net5227),
.C(net5276),
.Y(net5280)
);

HB1xp67_ASAP7_75t_R c5235(
.A(net10015),
.Y(net5281)
);

XOR2xp5_ASAP7_75t_R c5236(
.A(net5269),
.B(net5262),
.Y(net5282)
);

AND2x2_ASAP7_75t_R c5237(
.A(net5279),
.B(net4373),
.Y(net5283)
);

AND2x4_ASAP7_75t_R c5238(
.A(net3460),
.B(net10147),
.Y(net5284)
);

AND2x6_ASAP7_75t_R c5239(
.A(net2400),
.B(net5275),
.Y(net5285)
);

HAxp5_ASAP7_75t_R c5240(
.A(net5281),
.B(net5077),
.CON(net5286)
);

NAND2x1_ASAP7_75t_R c5241(
.A(net4429),
.B(net5284),
.Y(net5287)
);

HB2xp67_ASAP7_75t_R c5242(
.A(net5230),
.Y(net5288)
);

NAND2x1p5_ASAP7_75t_R c5243(
.A(net4426),
.B(net4399),
.Y(net5289)
);

NAND2x2_ASAP7_75t_R c5244(
.A(net4356),
.B(net4380),
.Y(net5290)
);

NAND2xp33_ASAP7_75t_R c5245(
.A(net9710),
.B(net10242),
.Y(net5291)
);

NAND2xp5_ASAP7_75t_R c5246(
.A(net4236),
.B(net2400),
.Y(net5292)
);

HB3xp67_ASAP7_75t_R c5247(
.A(net4403),
.Y(net5293)
);

NAND2xp67_ASAP7_75t_R c5248(
.A(net5187),
.B(net5293),
.Y(net5294)
);

NOR2x1_ASAP7_75t_R c5249(
.A(net4362),
.B(net4329),
.Y(net5295)
);

NOR2x1p5_ASAP7_75t_R c5250(
.A(net686),
.B(net9911),
.Y(net5296)
);

NOR2x2_ASAP7_75t_R c5251(
.A(net5278),
.B(net5257),
.Y(net5297)
);

HB4xp67_ASAP7_75t_R c5252(
.A(net5287),
.Y(net5298)
);

NOR2xp33_ASAP7_75t_R c5253(
.A(net5221),
.B(net3491),
.Y(net5299)
);

NOR2xp67_ASAP7_75t_R c5254(
.A(net5298),
.B(net4329),
.Y(net5300)
);

OR2x2_ASAP7_75t_R c5255(
.A(net4407),
.B(net3438),
.Y(net5301)
);

INVx11_ASAP7_75t_R c5256(
.A(net4047),
.Y(net5302)
);

OR2x4_ASAP7_75t_R c5257(
.A(net4380),
.B(net9696),
.Y(net5303)
);

OR2x6_ASAP7_75t_R c5258(
.A(net5222),
.B(net3483),
.Y(net5304)
);

INVx13_ASAP7_75t_R c5259(
.A(net4298),
.Y(net5305)
);

XNOR2x1_ASAP7_75t_R c5260(
.B(net4434),
.A(net4957),
.Y(net5306)
);

INVx1_ASAP7_75t_R c5261(
.A(net10386),
.Y(net5307)
);

INVx2_ASAP7_75t_R c5262(
.A(net10122),
.Y(net5308)
);

XNOR2x2_ASAP7_75t_R c5263(
.A(net5253),
.B(net3443),
.Y(net5309)
);

INVx3_ASAP7_75t_R c5264(
.A(net10169),
.Y(net5310)
);

XNOR2xp5_ASAP7_75t_R c5265(
.A(net5282),
.B(net4110),
.Y(net5311)
);

XOR2x1_ASAP7_75t_R c5266(
.A(net4368),
.B(net9710),
.Y(net5312)
);

XOR2x2_ASAP7_75t_R c5267(
.A(net5239),
.B(net4407),
.Y(net5313)
);

XOR2xp5_ASAP7_75t_R c5268(
.A(net5302),
.B(net4166),
.Y(net5314)
);

AND2x2_ASAP7_75t_R c5269(
.A(net5295),
.B(net5312),
.Y(net5315)
);

INVx4_ASAP7_75t_R c5270(
.A(net10133),
.Y(net5316)
);

AND2x4_ASAP7_75t_R c5271(
.A(net5283),
.B(net5277),
.Y(net5317)
);

INVx5_ASAP7_75t_R c5272(
.A(net9467),
.Y(net5318)
);

INVx6_ASAP7_75t_R c5273(
.A(net10533),
.Y(net5319)
);

AND2x6_ASAP7_75t_R c5274(
.A(net4389),
.B(net4310),
.Y(net5320)
);

HAxp5_ASAP7_75t_R c5275(
.A(net5304),
.B(net5293),
.CON(net5321)
);

INVx8_ASAP7_75t_R c5276(
.A(net10419),
.Y(net5322)
);

AND3x1_ASAP7_75t_R c5277(
.A(net4336),
.B(net677),
.C(net4425),
.Y(net5323)
);

NAND2x1_ASAP7_75t_R c5278(
.A(net5321),
.B(net4827),
.Y(net5324)
);

ICGx8DC_ASAP7_75t_R c5279(
.ENA(net4428),
.SE(net5306),
.CLK(clk),
.GCLK(net5325)
);

INVxp33_ASAP7_75t_R c5280(
.A(net5310),
.Y(net5326)
);

INVxp67_ASAP7_75t_R c5281(
.A(net5317),
.Y(net5327)
);

NAND2x1p5_ASAP7_75t_R c5282(
.A(net5323),
.B(net5325),
.Y(net5328)
);

NAND2x2_ASAP7_75t_R c5283(
.A(net5303),
.B(net4380),
.Y(net5329)
);

NAND2xp33_ASAP7_75t_R c5284(
.A(net5329),
.B(net5274),
.Y(net5330)
);

NAND2xp5_ASAP7_75t_R c5285(
.A(net5292),
.B(net5328),
.Y(net5331)
);

NAND2xp67_ASAP7_75t_R c5286(
.A(net4368),
.B(net5319),
.Y(net5332)
);

NOR2x1_ASAP7_75t_R c5287(
.A(net2399),
.B(net5140),
.Y(net5333)
);

NOR2x1p5_ASAP7_75t_R c5288(
.A(net4413),
.B(net5325),
.Y(net5334)
);

NOR2x2_ASAP7_75t_R c5289(
.A(net5327),
.B(net5274),
.Y(net5335)
);

AND3x2_ASAP7_75t_R c5290(
.A(net5313),
.B(net5330),
.C(net5325),
.Y(net5336)
);

NOR2xp33_ASAP7_75t_R c5291(
.A(net5328),
.B(net5336),
.Y(net5337)
);

NOR2xp67_ASAP7_75t_R c5292(
.A(net4264),
.B(net5221),
.Y(net5338)
);

BUFx10_ASAP7_75t_R c5293(
.A(net10118),
.Y(net5339)
);

OR2x2_ASAP7_75t_R c5294(
.A(net5326),
.B(net5173),
.Y(net5340)
);

AOI33xp33_ASAP7_75t_R c5295(
.A1(net5277),
.A2(net5340),
.A3(net4379),
.B1(net5290),
.B2(net10044),
.B3(net10259),
.Y(net5341)
);

OR2x4_ASAP7_75t_R c5296(
.A(net5333),
.B(net5332),
.Y(net5342)
);

BUFx12_ASAP7_75t_R c5297(
.A(net10451),
.Y(net5343)
);

AND3x4_ASAP7_75t_R c5298(
.A(net5341),
.B(net5305),
.C(net3878),
.Y(net5344)
);

OA222x2_ASAP7_75t_R c5299(
.A1(net3428),
.A2(net5340),
.B1(net5341),
.B2(out25),
.C1(net5325),
.C2(net4373),
.Y(net5345)
);

AO21x1_ASAP7_75t_R c5300(
.A1(net5339),
.A2(net4968),
.B(net5334),
.Y(net5346)
);

BUFx12f_ASAP7_75t_R c5301(
.A(net10129),
.Y(net5347)
);

AO21x2_ASAP7_75t_R c5302(
.A1(net5289),
.A2(net5344),
.B(net5347),
.Y(net5348)
);

SDFHx2_ASAP7_75t_R c5303(
.D(net5331),
.SE(net5328),
.SI(net5347),
.CLK(clk),
.QN(net5349)
);

AOI32xp33_ASAP7_75t_R c5304(
.A1(net4827),
.A2(net5340),
.A3(net5343),
.B1(net5325),
.B2(out25),
.Y(net5350)
);

OA33x2_ASAP7_75t_R c5305(
.A1(net5307),
.A2(net5346),
.A3(net5347),
.B1(net4264),
.B2(net5135),
.B3(net10044),
.Y(net5351)
);

OR2x6_ASAP7_75t_R c5306(
.A(net5308),
.B(net5347),
.Y(net5352)
);

OAI222xp33_ASAP7_75t_R c5307(
.A1(net5352),
.A2(net4302),
.B1(net5290),
.B2(net5325),
.C1(net9790),
.C2(net10242),
.Y(net5353)
);

AOI21x1_ASAP7_75t_R c5308(
.A1(net5147),
.A2(net5348),
.B(net10100),
.Y(net5354)
);

NAND5xp2_ASAP7_75t_R c5309(
.A(net5350),
.B(net5341),
.C(net4399),
.D(net5347),
.E(net4357),
.Y(net5355)
);

AOI21xp33_ASAP7_75t_R c5310(
.A1(net5353),
.A2(net5354),
.B(net5322),
.Y(net5356)
);

SDFHx3_ASAP7_75t_R c5311(
.D(net5356),
.SE(net5347),
.SI(net5230),
.CLK(clk),
.QN(net5357)
);

XNOR2x1_ASAP7_75t_R c5312(
.B(net4379),
.A(net3537),
.Y(net5358)
);

NOR5xp2_ASAP7_75t_R c5313(
.A(net4445),
.B(net4379),
.C(net4446),
.D(net5182),
.E(net3557),
.Y(net5359)
);

BUFx16f_ASAP7_75t_R c5314(
.A(net10571),
.Y(net5360)
);

XNOR2x2_ASAP7_75t_R c5315(
.A(net4500),
.B(net3556),
.Y(net5361)
);

BUFx24_ASAP7_75t_R c5316(
.A(net10109),
.Y(net5362)
);

AOI21xp5_ASAP7_75t_R c5317(
.A1(net5362),
.A2(net4431),
.B(net5058),
.Y(net5363)
);

XNOR2xp5_ASAP7_75t_R c5318(
.A(net5285),
.B(net3564),
.Y(net5364)
);

XOR2x1_ASAP7_75t_R c5319(
.A(net4329),
.B(net5361),
.Y(net5365)
);

BUFx2_ASAP7_75t_R c5320(
.A(net10403),
.Y(net5366)
);

BUFx3_ASAP7_75t_R c5321(
.A(net10042),
.Y(net5367)
);

XOR2x2_ASAP7_75t_R c5322(
.A(net3578),
.B(net10229),
.Y(net5368)
);

XOR2xp5_ASAP7_75t_R c5323(
.A(net4464),
.B(net5293),
.Y(net5369)
);

BUFx4_ASAP7_75t_R c5324(
.A(net10078),
.Y(net5370)
);

AND2x2_ASAP7_75t_R c5325(
.A(net5153),
.B(net5361),
.Y(net5371)
);

AND2x4_ASAP7_75t_R c5326(
.A(net3578),
.B(net5314),
.Y(net5372)
);

AND2x6_ASAP7_75t_R c5327(
.A(net5316),
.B(net5334),
.Y(net5373)
);

HAxp5_ASAP7_75t_R c5328(
.A(net3315),
.B(net5348),
.CON(net5375),
.SN(net5374)
);

NAND2x1_ASAP7_75t_R c5329(
.A(net3543),
.B(net803),
.Y(net5376)
);

NAND2x1p5_ASAP7_75t_R c5330(
.A(net5227),
.B(net5373),
.Y(net5377)
);

NAND2x2_ASAP7_75t_R c5331(
.A(net5257),
.B(net5367),
.Y(net5378)
);

NAND2xp33_ASAP7_75t_R c5332(
.A(net5348),
.B(net4431),
.Y(net5379)
);

NAND2xp5_ASAP7_75t_R c5333(
.A(net5378),
.B(net5362),
.Y(net5380)
);

NAND2xp67_ASAP7_75t_R c5334(
.A(net5277),
.B(net5348),
.Y(net5381)
);

BUFx4f_ASAP7_75t_R c5335(
.A(net10054),
.Y(net5382)
);

BUFx5_ASAP7_75t_R c5336(
.A(net10352),
.Y(net5383)
);

FAx1_ASAP7_75t_R c5337(
.A(net5140),
.B(net2390),
.CI(net10259),
.SN(net5385),
.CON(net5384)
);

NOR2x1_ASAP7_75t_R c5338(
.A(net452),
.B(net5374),
.Y(net5386)
);

MAJIxp5_ASAP7_75t_R c5339(
.A(net3556),
.B(net5357),
.C(net4479),
.Y(net5387)
);

NOR2x1p5_ASAP7_75t_R c5340(
.A(net3562),
.B(net2990),
.Y(net5388)
);

NOR2x2_ASAP7_75t_R c5341(
.A(net4442),
.B(net5318),
.Y(net5389)
);

BUFx6f_ASAP7_75t_R c5342(
.A(net10159),
.Y(net5390)
);

NOR2xp33_ASAP7_75t_R c5343(
.A(net3571),
.B(net4110),
.Y(net5391)
);

NOR2xp67_ASAP7_75t_R c5344(
.A(net5335),
.B(net4501),
.Y(net5392)
);

MAJx2_ASAP7_75t_R c5345(
.A(net3582),
.B(net3315),
.C(net9641),
.Y(net5393)
);

OR2x2_ASAP7_75t_R c5346(
.A(net4505),
.B(net4479),
.Y(net5394)
);

OR2x4_ASAP7_75t_R c5347(
.A(net5375),
.B(net5394),
.Y(net5395)
);

MAJx3_ASAP7_75t_R c5348(
.A(net4380),
.B(net5290),
.C(net5314),
.Y(net5396)
);

OR2x6_ASAP7_75t_R c5349(
.A(net4425),
.B(net5369),
.Y(net5397)
);

XNOR2x1_ASAP7_75t_R c5350(
.B(net5389),
.A(net4442),
.Y(net5398)
);

NAND3x1_ASAP7_75t_R c5351(
.A(net5361),
.B(net5390),
.C(net4968),
.Y(net5399)
);

SDFHx4_ASAP7_75t_R c5352(
.D(net1664),
.SE(net5377),
.SI(net10228),
.CLK(clk),
.QN(net5400)
);

XNOR2x2_ASAP7_75t_R c5353(
.A(net4452),
.B(net5300),
.Y(net5401)
);

XNOR2xp5_ASAP7_75t_R c5354(
.A(net5360),
.B(net5375),
.Y(net5402)
);

XOR2x1_ASAP7_75t_R c5355(
.A(net5383),
.B(net5400),
.Y(net5403)
);

BUFx8_ASAP7_75t_R c5356(
.A(net10349),
.Y(net5404)
);

XOR2x2_ASAP7_75t_R c5357(
.A(net5381),
.B(net5390),
.Y(net5405)
);

XOR2xp5_ASAP7_75t_R c5358(
.A(net5398),
.B(net9697),
.Y(net5406)
);

AND2x2_ASAP7_75t_R c5359(
.A(net5366),
.B(net9754),
.Y(net5407)
);

AND2x4_ASAP7_75t_R c5360(
.A(net5391),
.B(net5376),
.Y(net5408)
);

SDFLx1_ASAP7_75t_R c5361(
.D(net5135),
.SE(net5400),
.SI(net3562),
.CLK(clk),
.QN(net5409)
);

AND2x6_ASAP7_75t_R c5362(
.A(net5380),
.B(net5408),
.Y(net5410)
);

NAND3x2_ASAP7_75t_R c5363(
.B(net748),
.C(net5376),
.A(net5257),
.Y(net5411)
);

HAxp5_ASAP7_75t_R c5364(
.A(net4110),
.B(net5409),
.CON(net5413),
.SN(net5412)
);

ICGx1_ASAP7_75t_R c5365(
.ENA(net5276),
.SE(net5406),
.CLK(clk),
.GCLK(net5414)
);

CKINVDCx10_ASAP7_75t_R c5366(
.A(net10456),
.Y(net5415)
);

NAND2x1_ASAP7_75t_R c5367(
.A(net5364),
.B(net5362),
.Y(net5416)
);

NAND2x1p5_ASAP7_75t_R c5368(
.A(net5405),
.B(net5416),
.Y(net5417)
);

NAND2x2_ASAP7_75t_R c5369(
.A(net5416),
.B(net10259),
.Y(net5418)
);

NAND3xp33_ASAP7_75t_R c5370(
.A(net4435),
.B(net5416),
.C(net5414),
.Y(net5419)
);

NAND2xp33_ASAP7_75t_R c5371(
.A(net3316),
.B(net5362),
.Y(net5420)
);

ICGx2_ASAP7_75t_R c5372(
.ENA(net2390),
.SE(net5392),
.CLK(clk),
.GCLK(net5421)
);

CKINVDCx11_ASAP7_75t_R c5373(
.A(net10484),
.Y(net5422)
);

NOR3x1_ASAP7_75t_R c5374(
.A(net4416),
.B(net5395),
.C(net5361),
.Y(net5423)
);

SDFLx2_ASAP7_75t_R c5375(
.D(net5382),
.SE(net5422),
.SI(net5417),
.CLK(clk),
.QN(net5424)
);

CKINVDCx12_ASAP7_75t_R c5376(
.A(net10500),
.Y(net5425)
);

NAND2xp5_ASAP7_75t_R c5377(
.A(net5358),
.B(net5368),
.Y(net5426)
);

NAND2xp67_ASAP7_75t_R c5378(
.A(net5192),
.B(net5418),
.Y(net5427)
);

NOR2x1_ASAP7_75t_R c5379(
.A(net5418),
.B(net5408),
.Y(net5428)
);

NOR3x2_ASAP7_75t_R c5380(
.B(net5318),
.C(net5404),
.A(net5427),
.Y(net5429)
);

NOR2x1p5_ASAP7_75t_R c5381(
.A(net5429),
.B(net5198),
.Y(net5430)
);

NOR2x2_ASAP7_75t_R c5382(
.A(net5173),
.B(net5410),
.Y(net5431)
);

NOR2xp33_ASAP7_75t_R c5383(
.A(net5424),
.B(net9641),
.Y(net5432)
);

OA221x2_ASAP7_75t_R c5384(
.A1(net5395),
.A2(net5432),
.B1(net4445),
.B2(net5361),
.C(net5419),
.Y(net5433)
);

OAI221xp5_ASAP7_75t_R c5385(
.A1(net5419),
.A2(net5370),
.B1(net5432),
.B2(net5418),
.C(net5411),
.Y(net5434)
);

NOR2xp67_ASAP7_75t_R c5386(
.A(net5372),
.B(net5379),
.Y(net5435)
);

OR2x2_ASAP7_75t_R c5387(
.A(net5425),
.B(net9779),
.Y(net5436)
);

OR2x4_ASAP7_75t_R c5388(
.A(net5420),
.B(net5396),
.Y(net5437)
);

OR2x6_ASAP7_75t_R c5389(
.A(net2601),
.B(net5427),
.Y(net5438)
);

NOR3xp33_ASAP7_75t_R c5390(
.A(net5390),
.B(net5417),
.C(net10260),
.Y(net5439)
);

OA21x2_ASAP7_75t_R c5391(
.A1(net5435),
.A2(net5374),
.B(net9949),
.Y(net5440)
);

OAI311xp33_ASAP7_75t_R c5392(
.A1(net4511),
.A2(net5428),
.A3(net4468),
.B1(net5414),
.C1(net10260),
.Y(net5441)
);

XNOR2x1_ASAP7_75t_R c5393(
.B(net5334),
.A(net5436),
.Y(net5442)
);

CKINVDCx14_ASAP7_75t_R c5394(
.A(net10109),
.Y(net5443)
);

OAI21x1_ASAP7_75t_R c5395(
.A1(net1798),
.A2(net3628),
.B(net5421),
.Y(net5444)
);

XNOR2x2_ASAP7_75t_R c5396(
.A(net3517),
.B(net5182),
.Y(net5445)
);

XNOR2xp5_ASAP7_75t_R c5397(
.A(net4307),
.B(net10218),
.Y(net5446)
);

XOR2x1_ASAP7_75t_R c5398(
.A(net5441),
.B(net3600),
.Y(net5447)
);

XOR2x2_ASAP7_75t_R c5399(
.A(net5421),
.B(net4432),
.Y(net5448)
);

CKINVDCx16_ASAP7_75t_R c5400(
.A(net10344),
.Y(net5449)
);

OAI22xp5_ASAP7_75t_R c5401(
.A1(net4571),
.A2(net4538),
.B1(net2707),
.B2(net4523),
.Y(net5450)
);

OAI321xp33_ASAP7_75t_R c5402(
.A1(net3626),
.A2(net4507),
.A3(net5357),
.B1(net4573),
.B2(net10245),
.C(net10247),
.Y(net5451)
);

ICGx2p67DC_ASAP7_75t_R c5403(
.ENA(net5288),
.SE(net4526),
.CLK(clk),
.GCLK(net5452)
);

OAI21xp33_ASAP7_75t_R c5404(
.A1(net5182),
.A2(net4598),
.B(net4589),
.Y(net5453)
);

OAI21xp5_ASAP7_75t_R c5405(
.A1(net1759),
.A2(net3673),
.B(net3537),
.Y(net5454)
);

OR3x1_ASAP7_75t_R c5406(
.A(net4546),
.B(net4598),
.C(net10248),
.Y(net5455)
);

SDFLx3_ASAP7_75t_R c5407(
.D(net4585),
.SE(net4535),
.SI(net5438),
.CLK(clk),
.QN(net5456)
);

CKINVDCx20_ASAP7_75t_R c5408(
.A(net10494),
.Y(net5457)
);

XOR2xp5_ASAP7_75t_R c5409(
.A(net4522),
.B(net3674),
.Y(net5458)
);

AND2x2_ASAP7_75t_R c5410(
.A(net4598),
.B(net4546),
.Y(net5459)
);

AND2x4_ASAP7_75t_R c5411(
.A(net2590),
.B(net4357),
.Y(net5460)
);

AND2x6_ASAP7_75t_R c5412(
.A(net4432),
.B(net9772),
.Y(net5461)
);

HAxp5_ASAP7_75t_R c5413(
.A(net5458),
.B(net5288),
.CON(out16),
.SN(net5462)
);

OR3x2_ASAP7_75t_R c5414(
.A(net5438),
.B(net3667),
.C(net9858),
.Y(net5463)
);

OR3x4_ASAP7_75t_R c5415(
.A(net2682),
.B(net5438),
.C(net5456),
.Y(net5464)
);

AND3x1_ASAP7_75t_R c5416(
.A(net4507),
.B(net5455),
.C(net2578),
.Y(net5465)
);

NAND2x1_ASAP7_75t_R c5417(
.A(net5445),
.B(net2712),
.Y(net5466)
);

NAND2x1p5_ASAP7_75t_R c5418(
.A(net4591),
.B(net5424),
.Y(net5467)
);

NAND2x2_ASAP7_75t_R c5419(
.A(net4556),
.B(net4566),
.Y(net5468)
);

NAND2xp33_ASAP7_75t_R c5420(
.A(net3644),
.B(net10248),
.Y(net5469)
);

AND3x2_ASAP7_75t_R c5421(
.A(net3667),
.B(net3626),
.C(net4572),
.Y(net5470)
);

SDFLx4_ASAP7_75t_R c5422(
.D(net3650),
.SE(net5441),
.SI(net3676),
.CLK(clk),
.QN(net5471)
);

NAND2xp5_ASAP7_75t_R c5423(
.A(net4446),
.B(net677),
.Y(net5472)
);

NAND2xp67_ASAP7_75t_R c5424(
.A(net5459),
.B(net5454),
.Y(net5473)
);

NOR2x1_ASAP7_75t_R c5425(
.A(net5455),
.B(net5290),
.Y(net5474)
);

AND3x4_ASAP7_75t_R c5426(
.A(net5376),
.B(net4478),
.C(net10245),
.Y(net5475)
);

AO21x1_ASAP7_75t_R c5427(
.A1(net3643),
.A2(net5456),
.B(net9836),
.Y(net5476)
);

AO21x2_ASAP7_75t_R c5428(
.A1(net5403),
.A2(net2617),
.B(net4099),
.Y(net5477)
);

NOR2x1p5_ASAP7_75t_R c5429(
.A(net5454),
.B(net10248),
.Y(net5478)
);

NOR2x2_ASAP7_75t_R c5430(
.A(net5475),
.B(net3652),
.Y(net5479)
);

AOI21x1_ASAP7_75t_R c5431(
.A1(net5468),
.A2(net2682),
.B(net3639),
.Y(net5480)
);

ICGx3_ASAP7_75t_R c5432(
.ENA(net3608),
.SE(net5376),
.CLK(clk),
.GCLK(net5481)
);

AOI21xp33_ASAP7_75t_R c5433(
.A1(net4579),
.A2(net2708),
.B(net3639),
.Y(net5482)
);

CKINVDCx5p33_ASAP7_75t_R c5434(
.A(net10428),
.Y(net5483)
);

NOR2xp33_ASAP7_75t_R c5435(
.A(net3673),
.B(net10203),
.Y(net5484)
);

AOI21xp5_ASAP7_75t_R c5436(
.A1(net1720),
.A2(net5478),
.B(net9707),
.Y(net5485)
);

DFFASRHQNx1_ASAP7_75t_R c5437(
.D(net4572),
.RESETN(net5475),
.SETN(net3655),
.CLK(clk),
.QN(net5486)
);

FAx1_ASAP7_75t_R c5438(
.A(net4478),
.B(net2578),
.CI(net4432),
.SN(net5488),
.CON(net5487)
);

NOR2xp67_ASAP7_75t_R c5439(
.A(net2463),
.B(net5485),
.Y(net5489)
);

MAJIxp5_ASAP7_75t_R c5440(
.A(net5457),
.B(net4540),
.C(net10247),
.Y(net5490)
);

MAJx2_ASAP7_75t_R c5441(
.A(net4539),
.B(net4572),
.C(net4535),
.Y(net5491)
);

SDFHx1_ASAP7_75t_R c5442(
.D(net5399),
.SE(net5481),
.SI(net5475),
.CLK(clk),
.QN(net5492)
);

OR2x2_ASAP7_75t_R c5443(
.A(net5480),
.B(net5481),
.Y(net5493)
);

MAJx3_ASAP7_75t_R c5444(
.A(net5471),
.B(net4522),
.C(net5475),
.Y(net5494)
);

OR2x4_ASAP7_75t_R c5445(
.A(net5489),
.B(net5421),
.Y(net5495)
);

SDFHx2_ASAP7_75t_R c5446(
.D(net5450),
.SE(net5487),
.SI(net3650),
.CLK(clk),
.QN(net5496)
);

CKINVDCx6p67_ASAP7_75t_R c5447(
.A(net10344),
.Y(net5497)
);

NAND3x1_ASAP7_75t_R c5448(
.A(net5497),
.B(net2682),
.C(net9895),
.Y(net5498)
);

OR2x6_ASAP7_75t_R c5449(
.A(net3600),
.B(net4540),
.Y(net5499)
);

XNOR2x1_ASAP7_75t_R c5450(
.B(net5476),
.A(net2712),
.Y(net5500)
);

NAND3x2_ASAP7_75t_R c5451(
.B(net5474),
.C(net5475),
.A(net5471),
.Y(net5501)
);

CKINVDCx8_ASAP7_75t_R c5452(
.A(net10468),
.Y(net5502)
);

XNOR2x2_ASAP7_75t_R c5453(
.A(net5498),
.B(net5474),
.Y(net5503)
);

SDFHx3_ASAP7_75t_R c5454(
.D(net5469),
.SE(net5503),
.SI(net4591),
.CLK(clk),
.QN(net5504)
);

NAND3xp33_ASAP7_75t_R c5455(
.A(net5500),
.B(net5467),
.C(net10218),
.Y(net5505)
);

SDFHx4_ASAP7_75t_R c5456(
.D(net5477),
.SE(net5488),
.SI(net5495),
.CLK(clk),
.QN(net5506)
);

SDFLx1_ASAP7_75t_R c5457(
.D(net5488),
.SE(net3618),
.SI(net5403),
.CLK(clk),
.QN(net5507)
);

NOR3x1_ASAP7_75t_R c5458(
.A(net5504),
.B(net5486),
.C(net5467),
.Y(net5508)
);

NOR3x2_ASAP7_75t_R c5459(
.B(net3537),
.C(net4573),
.A(net5504),
.Y(net5509)
);

NOR3xp33_ASAP7_75t_R c5460(
.A(net4526),
.B(net5473),
.C(net5454),
.Y(net5510)
);

XNOR2xp5_ASAP7_75t_R c5461(
.A(net5506),
.B(net5504),
.Y(net5511)
);

OA21x2_ASAP7_75t_R c5462(
.A1(net5509),
.A2(net5424),
.B(net5495),
.Y(net5512)
);

SDFLx2_ASAP7_75t_R c5463(
.D(net4562),
.SE(net5505),
.SI(net5485),
.CLK(clk),
.QN(net5513)
);

CKINVDCx9p33_ASAP7_75t_R c5464(
.A(net10419),
.Y(net5514)
);

XOR2x1_ASAP7_75t_R c5465(
.A(net4563),
.B(net5501),
.Y(net5515)
);

SDFLx3_ASAP7_75t_R c5466(
.D(net5499),
.SE(net5506),
.SI(net5489),
.CLK(clk),
.QN(net5516)
);

OAI21x1_ASAP7_75t_R c5467(
.A1(net4595),
.A2(net5422),
.B(net5512),
.Y(net5517)
);

OAI21xp33_ASAP7_75t_R c5468(
.A1(net5493),
.A2(net5509),
.B(net5495),
.Y(net5518)
);

OAI21xp5_ASAP7_75t_R c5469(
.A1(net5454),
.A2(net5504),
.B(net5459),
.Y(net5519)
);

SDFLx4_ASAP7_75t_R c5470(
.D(net5508),
.SE(net4525),
.SI(net9871),
.CLK(clk),
.QN(net5520)
);

OAI31xp33_ASAP7_75t_R c5471(
.A1(net5484),
.A2(net5486),
.A3(net5520),
.B(net10218),
.Y(net5521)
);

XOR2x2_ASAP7_75t_R c5472(
.A(net4565),
.B(net5498),
.Y(net5522)
);

OR3x1_ASAP7_75t_R c5473(
.A(net5466),
.B(net5492),
.C(net9943),
.Y(net5523)
);

OAI33xp33_ASAP7_75t_R c5474(
.A1(net5441),
.A2(net5492),
.A3(out25),
.B1(net5456),
.B2(net9911),
.B3(net10203),
.Y(net5524)
);

AO222x2_ASAP7_75t_R c5475(
.A1(net5522),
.A2(net5523),
.B1(net5520),
.B2(net5376),
.C1(out25),
.C2(net10228),
.Y(net5525)
);

OR3x2_ASAP7_75t_R c5476(
.A(net5519),
.B(net5521),
.C(net10262),
.Y(net5526)
);

OR3x4_ASAP7_75t_R c5477(
.A(net5497),
.B(net5526),
.C(net10262),
.Y(net5527)
);

XOR2xp5_ASAP7_75t_R c5478(
.A(net4665),
.B(net2795),
.Y(net5528)
);

HB1xp67_ASAP7_75t_R c5479(
.A(net4635),
.Y(net5529)
);

HB2xp67_ASAP7_75t_R c5480(
.A(net4657),
.Y(net5530)
);

HB3xp67_ASAP7_75t_R c5481(
.A(net4635),
.Y(net5531)
);

HB4xp67_ASAP7_75t_R c5482(
.A(net4651),
.Y(net5532)
);

INVx11_ASAP7_75t_R c5483(
.A(net2795),
.Y(net5533)
);

INVx13_ASAP7_75t_R c5484(
.A(net4619),
.Y(net5534)
);

INVx1_ASAP7_75t_R c5485(
.A(net5530),
.Y(net5535)
);

INVx2_ASAP7_75t_R c5486(
.A(net3694),
.Y(net5536)
);

ICGx4DC_ASAP7_75t_R c5487(
.ENA(net4624),
.SE(net4681),
.CLK(clk),
.GCLK(net5537)
);

INVx3_ASAP7_75t_R c5488(
.A(net4668),
.Y(net5538)
);

INVx4_ASAP7_75t_R c5489(
.A(net5535),
.Y(net5539)
);

INVx5_ASAP7_75t_R c5490(
.A(net4684),
.Y(net5540)
);

INVx6_ASAP7_75t_R c5491(
.A(net3722),
.Y(net5541)
);

AND2x2_ASAP7_75t_R c5492(
.A(net4618),
.B(net5541),
.Y(net5542)
);

AND2x4_ASAP7_75t_R c5493(
.A(net4617),
.B(net5541),
.Y(net5543)
);

INVx8_ASAP7_75t_R c5494(
.A(net4676),
.Y(net5544)
);

AND2x6_ASAP7_75t_R c5495(
.A(net4656),
.B(net2754),
.Y(net5545)
);

INVxp33_ASAP7_75t_R c5496(
.A(net3760),
.Y(net5546)
);

INVxp67_ASAP7_75t_R c5497(
.A(net947),
.Y(net5547)
);

BUFx10_ASAP7_75t_R c5498(
.A(net9184),
.Y(net5548)
);

BUFx12_ASAP7_75t_R c5499(
.A(net4676),
.Y(net5549)
);

BUFx12f_ASAP7_75t_R c5500(
.A(net9184),
.Y(net5550)
);

BUFx16f_ASAP7_75t_R c5501(
.A(net5538),
.Y(net5551)
);

BUFx24_ASAP7_75t_R c5502(
.A(net9203),
.Y(net5552)
);

HAxp5_ASAP7_75t_R c5503(
.A(net975),
.B(net4619),
.CON(net5554),
.SN(net5553)
);

ICGx4_ASAP7_75t_R c5504(
.ENA(net5531),
.SE(net10249),
.CLK(clk),
.GCLK(net5555)
);

BUFx2_ASAP7_75t_R c5505(
.A(net5544),
.Y(net5556)
);

BUFx3_ASAP7_75t_R c5506(
.A(net4660),
.Y(net5557)
);

ICGx5_ASAP7_75t_R c5507(
.ENA(net5535),
.SE(net3701),
.CLK(clk),
.GCLK(net5558)
);

AND3x1_ASAP7_75t_R c5508(
.A(net5538),
.B(net4667),
.C(net4616),
.Y(net5559)
);

NAND2x1_ASAP7_75t_R c5509(
.A(net5550),
.B(net5535),
.Y(net5560)
);

BUFx4_ASAP7_75t_R c5510(
.A(net10252),
.Y(net5561)
);

NAND2x1p5_ASAP7_75t_R c5511(
.A(net5557),
.B(net10249),
.Y(net5562)
);

BUFx4f_ASAP7_75t_R c5512(
.A(net9660),
.Y(net5563)
);

BUFx5_ASAP7_75t_R c5513(
.A(net3746),
.Y(net5564)
);

BUFx6f_ASAP7_75t_R c5514(
.A(net5558),
.Y(net5565)
);

AND3x2_ASAP7_75t_R c5515(
.A(net5564),
.B(net5535),
.C(net5551),
.Y(net5566)
);

NAND2x2_ASAP7_75t_R c5516(
.A(net3694),
.B(net4656),
.Y(net5567)
);

BUFx8_ASAP7_75t_R c5517(
.A(net5562),
.Y(net5568)
);

CKINVDCx10_ASAP7_75t_R c5518(
.A(net5537),
.Y(net5569)
);

CKINVDCx11_ASAP7_75t_R c5519(
.A(net9310),
.Y(net5570)
);

CKINVDCx12_ASAP7_75t_R c5520(
.A(net5564),
.Y(net5571)
);

CKINVDCx14_ASAP7_75t_R c5521(
.A(net5542),
.Y(net5572)
);

NAND2xp33_ASAP7_75t_R c5522(
.A(net5568),
.B(net5549),
.Y(net5573)
);

CKINVDCx16_ASAP7_75t_R c5523(
.A(net4629),
.Y(net5574)
);

CKINVDCx20_ASAP7_75t_R c5524(
.A(net5570),
.Y(net5575)
);

CKINVDCx5p33_ASAP7_75t_R c5525(
.A(net9233),
.Y(net5576)
);

NAND2xp5_ASAP7_75t_R c5526(
.A(net5550),
.B(net5551),
.Y(net5577)
);

NAND2xp67_ASAP7_75t_R c5527(
.A(net1904),
.B(net5559),
.Y(net5578)
);

AND3x4_ASAP7_75t_R c5528(
.A(net5565),
.B(net5575),
.C(net4609),
.Y(net5579)
);

ICGx5p33DC_ASAP7_75t_R c5529(
.ENA(net4624),
.SE(net5529),
.CLK(clk),
.GCLK(net5580)
);

CKINVDCx6p67_ASAP7_75t_R c5530(
.A(net9247),
.Y(net5581)
);

CKINVDCx8_ASAP7_75t_R c5531(
.A(net5559),
.Y(net5582)
);

CKINVDCx9p33_ASAP7_75t_R c5532(
.A(net4651),
.Y(net5583)
);

HB1xp67_ASAP7_75t_R c5533(
.A(net5555),
.Y(net5584)
);

HB2xp67_ASAP7_75t_R c5534(
.A(net5552),
.Y(net5585)
);

HB3xp67_ASAP7_75t_R c5535(
.A(net5580),
.Y(net5586)
);

NOR2x1_ASAP7_75t_R c5536(
.A(net5577),
.B(net5586),
.Y(net5587)
);

ICGx6p67DC_ASAP7_75t_R c5537(
.ENA(net5582),
.SE(net2795),
.CLK(clk),
.GCLK(net5588)
);

HB4xp67_ASAP7_75t_R c5538(
.A(net5547),
.Y(net5589)
);

INVx11_ASAP7_75t_R c5539(
.A(net5579),
.Y(net5590)
);

INVx13_ASAP7_75t_R c5540(
.A(net9282),
.Y(net5591)
);

DFFASRHQNx1_ASAP7_75t_R c5541(
.D(net5578),
.RESETN(net5591),
.SETN(net5561),
.CLK(clk),
.QN(net5592)
);

AO21x1_ASAP7_75t_R c5542(
.A1(net5575),
.A2(net5564),
.B(net5591),
.Y(net5593)
);

AO21x2_ASAP7_75t_R c5543(
.A1(net5566),
.A2(net5558),
.B(net5565),
.Y(net5594)
);

AOI21x1_ASAP7_75t_R c5544(
.A1(net5583),
.A2(net5593),
.B(net5584),
.Y(net5595)
);

SDFHx1_ASAP7_75t_R c5545(
.D(net5591),
.SE(net5555),
.SI(net5536),
.CLK(clk),
.QN(net5596)
);

ICGx8DC_ASAP7_75t_R c5546(
.ENA(net5533),
.SE(net5595),
.CLK(clk),
.GCLK(net5597)
);

NOR2x1p5_ASAP7_75t_R c5547(
.A(net5592),
.B(net5597),
.Y(net5598)
);

AOI21xp33_ASAP7_75t_R c5548(
.A1(net5555),
.A2(net5584),
.B(net5591),
.Y(net5599)
);

AOI21xp5_ASAP7_75t_R c5549(
.A1(net5593),
.A2(net5563),
.B(net9665),
.Y(net5600)
);

OAI31xp67_ASAP7_75t_R c5550(
.A1(net5595),
.A2(net5580),
.A3(net5528),
.B(net5584),
.Y(net5601)
);

FAx1_ASAP7_75t_R c5551(
.A(net4625),
.B(net5597),
.CI(net10252),
.SN(net5603),
.CON(net5602)
);

NOR2x2_ASAP7_75t_R c5552(
.A(net5583),
.B(net9665),
.Y(net5604)
);

MAJIxp5_ASAP7_75t_R c5553(
.A(net5585),
.B(net5602),
.C(net3759),
.Y(net5605)
);

AO33x2_ASAP7_75t_R c5554(
.A1(net5569),
.A2(net5596),
.A3(net5580),
.B1(net5551),
.B2(net5574),
.B3(net4681),
.Y(net5606)
);

MAJx2_ASAP7_75t_R c5555(
.A(net5576),
.B(net5599),
.C(net10263),
.Y(net5607)
);

SDFHx2_ASAP7_75t_R c5556(
.D(net5603),
.SE(net3722),
.SI(net5574),
.CLK(clk),
.QN(net5608)
);

NOR2xp33_ASAP7_75t_R c5557(
.A(net5607),
.B(net5562),
.Y(net5609)
);

MAJx3_ASAP7_75t_R c5558(
.A(net5590),
.B(net5609),
.C(net975),
.Y(net5610)
);

OR4x1_ASAP7_75t_R c5559(
.A(net5608),
.B(net5604),
.C(net5607),
.D(net5610),
.Y(net5611)
);

OR4x2_ASAP7_75t_R c5560(
.A(net5586),
.B(net5608),
.C(net5542),
.D(net5609),
.Y(net5612)
);

INVx1_ASAP7_75t_R c5561(
.A(net4705),
.Y(net5613)
);

INVx2_ASAP7_75t_R c5562(
.A(net9951),
.Y(net5614)
);

NOR2xp67_ASAP7_75t_R c5563(
.A(net5543),
.B(net4697),
.Y(net5615)
);

OR2x2_ASAP7_75t_R c5564(
.A(net1974),
.B(net4762),
.Y(net5616)
);

INVx3_ASAP7_75t_R c5565(
.A(net4671),
.Y(net5617)
);

ICGx1_ASAP7_75t_R c5566(
.ENA(net4752),
.SE(net5529),
.CLK(clk),
.GCLK(net5618)
);

OR2x4_ASAP7_75t_R c5567(
.A(net5529),
.B(net9978),
.Y(net5619)
);

NAND3x1_ASAP7_75t_R c5568(
.A(net4755),
.B(net5553),
.C(net4711),
.Y(net5620)
);

OR2x6_ASAP7_75t_R c5569(
.A(net5545),
.B(net4715),
.Y(net5621)
);

XNOR2x1_ASAP7_75t_R c5570(
.B(net4645),
.A(net5618),
.Y(net5622)
);

XNOR2x2_ASAP7_75t_R c5571(
.A(net3772),
.B(net4650),
.Y(net5623)
);

XNOR2xp5_ASAP7_75t_R c5572(
.A(net1974),
.B(net10265),
.Y(net5624)
);

INVx4_ASAP7_75t_R c5573(
.A(net9113),
.Y(net5625)
);

XOR2x1_ASAP7_75t_R c5574(
.A(net4734),
.B(net5563),
.Y(net5626)
);

XOR2x2_ASAP7_75t_R c5575(
.A(net3747),
.B(net10250),
.Y(net5627)
);

INVx5_ASAP7_75t_R c5576(
.A(net4759),
.Y(net5628)
);

XOR2xp5_ASAP7_75t_R c5577(
.A(net3780),
.B(net4755),
.Y(net5629)
);

AND2x2_ASAP7_75t_R c5578(
.A(net4655),
.B(net5592),
.Y(net5630)
);

INVx6_ASAP7_75t_R c5579(
.A(net9930),
.Y(net5631)
);

INVx8_ASAP7_75t_R c5580(
.A(net9113),
.Y(net5632)
);

AND2x4_ASAP7_75t_R c5581(
.A(net4655),
.B(net9677),
.Y(net5633)
);

AND2x6_ASAP7_75t_R c5582(
.A(net5604),
.B(net5543),
.Y(net5634)
);

INVxp33_ASAP7_75t_R c5583(
.A(net5572),
.Y(net5635)
);

NAND3x2_ASAP7_75t_R c5584(
.B(net5634),
.C(net3780),
.A(net4692),
.Y(net5636)
);

INVxp67_ASAP7_75t_R c5585(
.A(net10527),
.Y(net5637)
);

BUFx10_ASAP7_75t_R c5586(
.A(net4711),
.Y(net5638)
);

BUFx12_ASAP7_75t_R c5587(
.A(net10575),
.Y(net5639)
);

NAND3xp33_ASAP7_75t_R c5588(
.A(net5534),
.B(net5529),
.C(net1833),
.Y(net5640)
);

BUFx12f_ASAP7_75t_R c5589(
.A(net5596),
.Y(net5641)
);

BUFx16f_ASAP7_75t_R c5590(
.A(net900),
.Y(net5642)
);

BUFx24_ASAP7_75t_R c5591(
.A(net9247),
.Y(net5643)
);

BUFx2_ASAP7_75t_R c5592(
.A(net2891),
.Y(net5644)
);

BUFx3_ASAP7_75t_R c5593(
.A(net10446),
.Y(net5645)
);

ICGx2_ASAP7_75t_R c5594(
.ENA(net5637),
.SE(net2877),
.CLK(clk),
.GCLK(net5646)
);

HAxp5_ASAP7_75t_R c5595(
.A(net4655),
.B(net2754),
.CON(net5647)
);

NAND2x1_ASAP7_75t_R c5596(
.A(net4723),
.B(net4705),
.Y(net5648)
);

NAND2x1p5_ASAP7_75t_R c5597(
.A(net5622),
.B(net5645),
.Y(net5649)
);

NAND2x2_ASAP7_75t_R c5598(
.A(net5646),
.B(net5622),
.Y(net5650)
);

BUFx4_ASAP7_75t_R c5599(
.A(net5614),
.Y(net5651)
);

BUFx4f_ASAP7_75t_R c5600(
.A(net9233),
.Y(net5652)
);

BUFx5_ASAP7_75t_R c5601(
.A(net10576),
.Y(net5653)
);

NAND2xp33_ASAP7_75t_R c5602(
.A(net5642),
.B(net9862),
.Y(net5654)
);

NAND2xp5_ASAP7_75t_R c5603(
.A(net5643),
.B(net4735),
.Y(net5655)
);

NAND2xp67_ASAP7_75t_R c5604(
.A(net5642),
.B(net5628),
.Y(net5656)
);

NOR2x1_ASAP7_75t_R c5605(
.A(net5644),
.B(net2891),
.Y(net5657)
);

BUFx6f_ASAP7_75t_R c5606(
.A(net5641),
.Y(net5658)
);

BUFx8_ASAP7_75t_R c5607(
.A(net10406),
.Y(net5659)
);

NOR2x1p5_ASAP7_75t_R c5608(
.A(net5638),
.B(net10250),
.Y(net5660)
);

SDFHx3_ASAP7_75t_R c5609(
.D(net5646),
.SE(net5657),
.SI(net4740),
.CLK(clk),
.QN(net5661)
);

NOR2x2_ASAP7_75t_R c5610(
.A(net5563),
.B(net4758),
.Y(net5662)
);

CKINVDCx10_ASAP7_75t_R c5611(
.A(net5571),
.Y(net5663)
);

CKINVDCx11_ASAP7_75t_R c5612(
.A(net5650),
.Y(net5664)
);

NOR3x1_ASAP7_75t_R c5613(
.A(net5635),
.B(net5649),
.C(net5623),
.Y(net5665)
);

ICGx2p67DC_ASAP7_75t_R c5614(
.ENA(net5627),
.SE(net5663),
.CLK(clk),
.GCLK(net5666)
);

NOR2xp33_ASAP7_75t_R c5615(
.A(net5662),
.B(net4773),
.Y(net5667)
);

CKINVDCx12_ASAP7_75t_R c5616(
.A(net9951),
.Y(net5668)
);

NOR2xp67_ASAP7_75t_R c5617(
.A(net5667),
.B(net5615),
.Y(net5669)
);

NOR3x2_ASAP7_75t_R c5618(
.B(net3827),
.C(net5662),
.A(net5661),
.Y(net5670)
);

OR2x2_ASAP7_75t_R c5619(
.A(net5669),
.B(net5667),
.Y(net5671)
);

A2O1A1Ixp33_ASAP7_75t_R c5620(
.A1(net4715),
.A2(net5635),
.B(net142),
.C(net10265),
.Y(net5672)
);

NOR3xp33_ASAP7_75t_R c5621(
.A(net5651),
.B(net5656),
.C(net4696),
.Y(net5673)
);

CKINVDCx14_ASAP7_75t_R c5622(
.A(net10412),
.Y(net5674)
);

OR2x4_ASAP7_75t_R c5623(
.A(net5653),
.B(net5645),
.Y(net5675)
);

OR2x6_ASAP7_75t_R c5624(
.A(net5652),
.B(net5635),
.Y(net5676)
);

OA21x2_ASAP7_75t_R c5625(
.A1(net5615),
.A2(net5656),
.B(net9766),
.Y(net5677)
);

XNOR2x1_ASAP7_75t_R c5626(
.B(net5654),
.A(net5656),
.Y(net5678)
);

AND4x1_ASAP7_75t_R c5627(
.A(net5671),
.B(net5629),
.C(net5661),
.D(net5610),
.Y(net5679)
);

XNOR2x2_ASAP7_75t_R c5628(
.A(net5673),
.B(net4732),
.Y(net5680)
);

CKINVDCx16_ASAP7_75t_R c5629(
.A(net9930),
.Y(net5681)
);

OAI21x1_ASAP7_75t_R c5630(
.A1(net5612),
.A2(net5667),
.B(net9929),
.Y(net5682)
);

XNOR2xp5_ASAP7_75t_R c5631(
.A(net5658),
.B(net3813),
.Y(net5683)
);

XOR2x1_ASAP7_75t_R c5632(
.A(net5663),
.B(net4681),
.Y(net5684)
);

AND4x2_ASAP7_75t_R c5633(
.A(net5677),
.B(net5643),
.C(net2891),
.D(net5657),
.Y(net5685)
);

OAI21xp33_ASAP7_75t_R c5634(
.A1(net5681),
.A2(net9884),
.B(net10266),
.Y(net5686)
);

SDFHx4_ASAP7_75t_R c5635(
.D(net5529),
.SE(net5641),
.SI(net9862),
.CLK(clk),
.QN(net5687)
);

CKINVDCx20_ASAP7_75t_R c5636(
.A(net10530),
.Y(net5688)
);

SDFLx1_ASAP7_75t_R c5637(
.D(net5687),
.SE(net5621),
.SI(net9930),
.CLK(clk),
.QN(net5689)
);

OAI21xp5_ASAP7_75t_R c5638(
.A1(net5683),
.A2(net5664),
.B(net4716),
.Y(net5690)
);

OR3x1_ASAP7_75t_R c5639(
.A(net5687),
.B(net5572),
.C(net10250),
.Y(net5691)
);

XOR2x2_ASAP7_75t_R c5640(
.A(net5691),
.B(net5681),
.Y(net5692)
);

OR3x2_ASAP7_75t_R c5641(
.A(net5675),
.B(net5691),
.C(net10266),
.Y(net5693)
);

AO211x2_ASAP7_75t_R c5642(
.A1(net5686),
.A2(net5677),
.B(net3701),
.C(net5691),
.Y(net5694)
);

AOI222xp33_ASAP7_75t_R c5643(
.A1(net5693),
.A2(net2877),
.B1(net5621),
.B2(net5657),
.C1(net5691),
.C2(net5548),
.Y(net5695)
);

CKINVDCx5p33_ASAP7_75t_R c5644(
.A(net4735),
.Y(net5696)
);

CKINVDCx6p67_ASAP7_75t_R c5645(
.A(net3836),
.Y(net5697)
);

XOR2xp5_ASAP7_75t_R c5646(
.A(net3699),
.B(net2891),
.Y(net5698)
);

AND2x2_ASAP7_75t_R c5647(
.A(net4736),
.B(net5624),
.Y(net5699)
);

CKINVDCx8_ASAP7_75t_R c5648(
.A(net9235),
.Y(net5700)
);

CKINVDCx9p33_ASAP7_75t_R c5649(
.A(net9162),
.Y(net5701)
);

HB1xp67_ASAP7_75t_R c5650(
.A(net10268),
.Y(net5702)
);

HB2xp67_ASAP7_75t_R c5651(
.A(net4628),
.Y(net5703)
);

HB3xp67_ASAP7_75t_R c5652(
.A(net3813),
.Y(net5704)
);

OR3x4_ASAP7_75t_R c5653(
.A(net4758),
.B(net5702),
.C(net4851),
.Y(net5705)
);

AO22x1_ASAP7_75t_R c5654(
.A1(net4851),
.A2(net4735),
.B1(net5699),
.B2(net3922),
.Y(net5706)
);

AND2x4_ASAP7_75t_R c5655(
.A(net5659),
.B(net5705),
.Y(net5707)
);

AND2x6_ASAP7_75t_R c5656(
.A(net5666),
.B(net4681),
.Y(net5708)
);

HB4xp67_ASAP7_75t_R c5657(
.A(net9162),
.Y(net5709)
);

INVx11_ASAP7_75t_R c5658(
.A(net5699),
.Y(net5710)
);

HAxp5_ASAP7_75t_R c5659(
.A(net3925),
.B(net10268),
.CON(net5711)
);

INVx13_ASAP7_75t_R c5660(
.A(net9216),
.Y(net5712)
);

INVx1_ASAP7_75t_R c5661(
.A(net4761),
.Y(net5713)
);

NAND2x1_ASAP7_75t_R c5662(
.A(net5705),
.B(net5709),
.Y(net5714)
);

NAND2x1p5_ASAP7_75t_R c5663(
.A(net5655),
.B(net5592),
.Y(net5715)
);

INVx2_ASAP7_75t_R c5664(
.A(net5709),
.Y(net5716)
);

INVx3_ASAP7_75t_R c5665(
.A(net5624),
.Y(net5717)
);

INVx4_ASAP7_75t_R c5666(
.A(net10400),
.Y(net5718)
);

NAND2x2_ASAP7_75t_R c5667(
.A(net2996),
.B(net4840),
.Y(net5719)
);

AO22x2_ASAP7_75t_R c5668(
.A1(net5717),
.A2(net5699),
.B1(net5705),
.B2(net5702),
.Y(net5720)
);

AO31x2_ASAP7_75t_R c5669(
.A1(net5699),
.A2(net5666),
.A3(net5625),
.B(net5709),
.Y(net5721)
);

NAND2xp33_ASAP7_75t_R c5670(
.A(net5710),
.B(net4728),
.Y(net5722)
);

INVx5_ASAP7_75t_R c5671(
.A(net10438),
.Y(net5723)
);

NAND2xp5_ASAP7_75t_R c5672(
.A(net5713),
.B(net5702),
.Y(net5724)
);

NAND2xp67_ASAP7_75t_R c5673(
.A(net4681),
.B(net2891),
.Y(net5725)
);

INVx6_ASAP7_75t_R c5674(
.A(net4699),
.Y(net5726)
);

INVx8_ASAP7_75t_R c5675(
.A(net9926),
.Y(net5727)
);

NOR2x1_ASAP7_75t_R c5676(
.A(net5707),
.B(net5698),
.Y(net5728)
);

NOR2x1p5_ASAP7_75t_R c5677(
.A(net5724),
.B(net2891),
.Y(net5729)
);

AND3x1_ASAP7_75t_R c5678(
.A(net4807),
.B(net3872),
.C(net5645),
.Y(net5730)
);

INVxp33_ASAP7_75t_R c5679(
.A(net5719),
.Y(net5731)
);

INVxp67_ASAP7_75t_R c5680(
.A(net9870),
.Y(net5732)
);

BUFx10_ASAP7_75t_R c5681(
.A(net10016),
.Y(net5733)
);

BUFx12_ASAP7_75t_R c5682(
.A(net10402),
.Y(net5734)
);

BUFx12f_ASAP7_75t_R c5683(
.A(net5722),
.Y(net5735)
);

NOR2x2_ASAP7_75t_R c5684(
.A(net5698),
.B(net5713),
.Y(net5736)
);

BUFx16f_ASAP7_75t_R c5685(
.A(net5537),
.Y(net5737)
);

AND3x2_ASAP7_75t_R c5686(
.A(net4851),
.B(net4840),
.C(net9776),
.Y(net5738)
);

BUFx24_ASAP7_75t_R c5687(
.A(net9275),
.Y(net5739)
);

BUFx2_ASAP7_75t_R c5688(
.A(net10463),
.Y(net5740)
);

AND3x4_ASAP7_75t_R c5689(
.A(net5700),
.B(net5739),
.C(net4738),
.Y(net5741)
);

BUFx3_ASAP7_75t_R c5690(
.A(net5648),
.Y(net5742)
);

NOR2xp33_ASAP7_75t_R c5691(
.A(net5714),
.B(net5629),
.Y(net5743)
);

BUFx4_ASAP7_75t_R c5692(
.A(net9677),
.Y(net5744)
);

NOR2xp67_ASAP7_75t_R c5693(
.A(net5731),
.B(net5702),
.Y(net5745)
);

BUFx4f_ASAP7_75t_R c5694(
.A(net5737),
.Y(net5746)
);

OR2x2_ASAP7_75t_R c5695(
.A(net5664),
.B(net5709),
.Y(net5747)
);

AO21x1_ASAP7_75t_R c5696(
.A1(net5733),
.A2(net4793),
.B(net10268),
.Y(net5748)
);

AO21x2_ASAP7_75t_R c5697(
.A1(net5739),
.A2(net5746),
.B(net4788),
.Y(net5749)
);

OR2x4_ASAP7_75t_R c5698(
.A(net5727),
.B(net4788),
.Y(net5750)
);

OR2x6_ASAP7_75t_R c5699(
.A(net5715),
.B(net5696),
.Y(net5751)
);

BUFx5_ASAP7_75t_R c5700(
.A(net5732),
.Y(net5752)
);

XNOR2x1_ASAP7_75t_R c5701(
.B(net5740),
.A(net5692),
.Y(net5753)
);

BUFx6f_ASAP7_75t_R c5702(
.A(net4853),
.Y(net5754)
);

XNOR2x2_ASAP7_75t_R c5703(
.A(net5720),
.B(net5753),
.Y(net5755)
);

XNOR2xp5_ASAP7_75t_R c5704(
.A(net5750),
.B(net5698),
.Y(net5756)
);

XOR2x1_ASAP7_75t_R c5705(
.A(net4728),
.B(net5753),
.Y(net5757)
);

AOI21x1_ASAP7_75t_R c5706(
.A1(net5746),
.A2(net3922),
.B(net5753),
.Y(net5758)
);

BUFx8_ASAP7_75t_R c5707(
.A(net9993),
.Y(net5759)
);

AOI211x1_ASAP7_75t_R c5708(
.A1(net4824),
.A2(net5567),
.B(net5624),
.C(net4851),
.Y(net5760)
);

XOR2x2_ASAP7_75t_R c5709(
.A(net5749),
.B(net4714),
.Y(net5761)
);

CKINVDCx10_ASAP7_75t_R c5710(
.A(net10418),
.Y(net5762)
);

CKINVDCx11_ASAP7_75t_R c5711(
.A(net5762),
.Y(net5763)
);

CKINVDCx12_ASAP7_75t_R c5712(
.A(net10404),
.Y(net5764)
);

XOR2xp5_ASAP7_75t_R c5713(
.A(net5758),
.B(net4834),
.Y(net5765)
);

AND2x2_ASAP7_75t_R c5714(
.A(net5639),
.B(net5707),
.Y(net5766)
);

CKINVDCx14_ASAP7_75t_R c5715(
.A(net10116),
.Y(net5767)
);

AOI21xp33_ASAP7_75t_R c5716(
.A1(net4817),
.A2(net5766),
.B(net5758),
.Y(net5768)
);

AND2x4_ASAP7_75t_R c5717(
.A(net5764),
.B(net5766),
.Y(net5769)
);

SDFLx2_ASAP7_75t_R c5718(
.D(net5755),
.SE(net5736),
.SI(net5767),
.CLK(clk),
.QN(net5770)
);

AOI21xp5_ASAP7_75t_R c5719(
.A1(net5716),
.A2(net5718),
.B(net5705),
.Y(net5771)
);

SDFLx3_ASAP7_75t_R c5720(
.D(net5761),
.SE(net5736),
.SI(net5697),
.CLK(clk),
.QN(net5772)
);

FAx1_ASAP7_75t_R c5721(
.A(net5759),
.B(net5705),
.CI(net4851),
.SN(net5774),
.CON(net5773)
);

AND2x6_ASAP7_75t_R c5722(
.A(net5767),
.B(net10171),
.Y(net5775)
);

HAxp5_ASAP7_75t_R c5723(
.A(net5773),
.B(net9693),
.CON(net5776)
);

NAND2x1_ASAP7_75t_R c5724(
.A(net5739),
.B(net9909),
.Y(net5777)
);

MAJIxp5_ASAP7_75t_R c5725(
.A(net5754),
.B(net5755),
.C(net5777),
.Y(net5778)
);

SDFLx4_ASAP7_75t_R c5726(
.D(net5777),
.SE(net5778),
.SI(net5769),
.CLK(clk),
.QN(net5779)
);

MAJx2_ASAP7_75t_R c5727(
.A(net5585),
.B(net4736),
.C(net5748),
.Y(net5780)
);

AOI211xp5_ASAP7_75t_R c5728(
.A1(net4859),
.A2(net5599),
.B(net3989),
.C(net2891),
.Y(net5781)
);

CKINVDCx16_ASAP7_75t_R c5729(
.A(net5723),
.Y(net5782)
);

CKINVDCx20_ASAP7_75t_R c5730(
.A(net10070),
.Y(net5783)
);

CKINVDCx5p33_ASAP7_75t_R c5731(
.A(net5753),
.Y(net5784)
);

NAND2x1p5_ASAP7_75t_R c5732(
.A(net5692),
.B(net4908),
.Y(net5785)
);

CKINVDCx6p67_ASAP7_75t_R c5733(
.A(net5632),
.Y(net5786)
);

CKINVDCx8_ASAP7_75t_R c5734(
.A(net3086),
.Y(net5787)
);

NAND2x2_ASAP7_75t_R c5735(
.A(net1196),
.B(net4905),
.Y(net5788)
);

CKINVDCx9p33_ASAP7_75t_R c5736(
.A(net2095),
.Y(net5789)
);

HB1xp67_ASAP7_75t_R c5737(
.A(net9160),
.Y(net5790)
);

HB2xp67_ASAP7_75t_R c5738(
.A(net9160),
.Y(net5791)
);

NAND2xp33_ASAP7_75t_R c5739(
.A(net4879),
.B(net5775),
.Y(net5792)
);

ICGx3_ASAP7_75t_R c5740(
.ENA(net2149),
.SE(net272),
.CLK(clk),
.GCLK(net5793)
);

HB3xp67_ASAP7_75t_R c5741(
.A(net9275),
.Y(net5794)
);

HB4xp67_ASAP7_75t_R c5742(
.A(net4914),
.Y(net5795)
);

NAND2xp5_ASAP7_75t_R c5743(
.A(net5592),
.B(net5748),
.Y(net5796)
);

INVx11_ASAP7_75t_R c5744(
.A(net5782),
.Y(net5797)
);

NAND2xp67_ASAP7_75t_R c5745(
.A(net5789),
.B(net4843),
.Y(net5798)
);

NOR2x1_ASAP7_75t_R c5746(
.A(net4938),
.B(net3079),
.Y(net5799)
);

INVx13_ASAP7_75t_R c5747(
.A(net4923),
.Y(net5800)
);

OAI32xp33_ASAP7_75t_R c5748(
.A1(net5799),
.A2(net4920),
.A3(net2034),
.B1(net3942),
.B2(net5797),
.Y(net5801)
);

INVx1_ASAP7_75t_R c5749(
.A(net4843),
.Y(net5802)
);

INVx2_ASAP7_75t_R c5750(
.A(net10460),
.Y(net5803)
);

NOR2x1p5_ASAP7_75t_R c5751(
.A(net3952),
.B(net10269),
.Y(net5804)
);

INVx3_ASAP7_75t_R c5752(
.A(net5803),
.Y(net5805)
);

INVx4_ASAP7_75t_R c5753(
.A(net5785),
.Y(net5806)
);

INVx5_ASAP7_75t_R c5754(
.A(net2117),
.Y(net5807)
);

NOR2x2_ASAP7_75t_R c5755(
.A(net5744),
.B(net3054),
.Y(net5808)
);

NOR2xp33_ASAP7_75t_R c5756(
.A(net5783),
.B(net4773),
.Y(net5809)
);

NOR2xp67_ASAP7_75t_R c5757(
.A(net5798),
.B(net4859),
.Y(net5810)
);

OR2x2_ASAP7_75t_R c5758(
.A(net4714),
.B(net5798),
.Y(net5811)
);

OR2x4_ASAP7_75t_R c5759(
.A(net5794),
.B(net4933),
.Y(net5812)
);

OR2x6_ASAP7_75t_R c5760(
.A(net5797),
.B(net4879),
.Y(net5813)
);

INVx6_ASAP7_75t_R c5761(
.A(net10556),
.Y(net5814)
);

XNOR2x1_ASAP7_75t_R c5762(
.B(net1163),
.A(net5814),
.Y(net5815)
);

INVx8_ASAP7_75t_R c5763(
.A(net4773),
.Y(net5816)
);

INVxp33_ASAP7_75t_R c5764(
.A(net9218),
.Y(net5817)
);

ICGx4DC_ASAP7_75t_R c5765(
.ENA(net4893),
.SE(net3942),
.CLK(clk),
.GCLK(net5818)
);

XNOR2x2_ASAP7_75t_R c5766(
.A(net5805),
.B(net5798),
.Y(net5819)
);

INVxp67_ASAP7_75t_R c5767(
.A(net5817),
.Y(net5820)
);

XNOR2xp5_ASAP7_75t_R c5768(
.A(net5792),
.B(net5819),
.Y(net5821)
);

BUFx10_ASAP7_75t_R c5769(
.A(net5812),
.Y(net5822)
);

BUFx12_ASAP7_75t_R c5770(
.A(net4875),
.Y(net5823)
);

XOR2x1_ASAP7_75t_R c5771(
.A(net5787),
.B(net5818),
.Y(net5824)
);

MAJx3_ASAP7_75t_R c5772(
.A(net5782),
.B(net5745),
.C(net5802),
.Y(net5825)
);

AOI22x1_ASAP7_75t_R c5773(
.A1(net4935),
.A2(net5628),
.B1(net5802),
.B2(net10266),
.Y(net5826)
);

XOR2x2_ASAP7_75t_R c5774(
.A(net5678),
.B(net5747),
.Y(net5827)
);

XOR2xp5_ASAP7_75t_R c5775(
.A(net5554),
.B(net5763),
.Y(net5828)
);

BUFx12f_ASAP7_75t_R c5776(
.A(net5828),
.Y(net5829)
);

AND2x2_ASAP7_75t_R c5777(
.A(net4010),
.B(net4870),
.Y(net5830)
);

BUFx16f_ASAP7_75t_R c5778(
.A(net4858),
.Y(net5831)
);

BUFx24_ASAP7_75t_R c5779(
.A(net5814),
.Y(net5832)
);

AND2x4_ASAP7_75t_R c5780(
.A(net3963),
.B(net5795),
.Y(net5833)
);

BUFx2_ASAP7_75t_R c5781(
.A(net5811),
.Y(net5834)
);

AND2x6_ASAP7_75t_R c5782(
.A(net5795),
.B(net5797),
.Y(net5835)
);

BUFx3_ASAP7_75t_R c5783(
.A(net4917),
.Y(net5836)
);

HAxp5_ASAP7_75t_R c5784(
.A(net5789),
.B(net4920),
.CON(net5837)
);

NAND2x1_ASAP7_75t_R c5785(
.A(net5825),
.B(net3772),
.Y(net5838)
);

BUFx4_ASAP7_75t_R c5786(
.A(net10128),
.Y(net5839)
);

AOI22xp33_ASAP7_75t_R c5787(
.A1(net5832),
.A2(net5810),
.B1(net5824),
.B2(net10269),
.Y(net5840)
);

NAND2x1p5_ASAP7_75t_R c5788(
.A(net5816),
.B(net3015),
.Y(net5841)
);

BUFx4f_ASAP7_75t_R c5789(
.A(net5822),
.Y(net5842)
);

NAND3x1_ASAP7_75t_R c5790(
.A(net5806),
.B(net5837),
.C(net5819),
.Y(net5843)
);

NAND2x2_ASAP7_75t_R c5791(
.A(net5800),
.B(net5810),
.Y(net5844)
);

NAND2xp33_ASAP7_75t_R c5792(
.A(net2090),
.B(net5844),
.Y(net5845)
);

NAND2xp5_ASAP7_75t_R c5793(
.A(net5833),
.B(net10164),
.Y(net5846)
);

NAND2xp67_ASAP7_75t_R c5794(
.A(net5838),
.B(net5835),
.Y(net5847)
);

BUFx5_ASAP7_75t_R c5795(
.A(net10487),
.Y(net5848)
);

NAND3x2_ASAP7_75t_R c5796(
.B(net5743),
.C(net5818),
.A(net5835),
.Y(net5849)
);

NAND3xp33_ASAP7_75t_R c5797(
.A(net5844),
.B(net5849),
.C(net4938),
.Y(net5850)
);

NOR3x1_ASAP7_75t_R c5798(
.A(net3859),
.B(net5834),
.C(net5848),
.Y(net5851)
);

NOR2x1_ASAP7_75t_R c5799(
.A(net5840),
.B(net5838),
.Y(net5852)
);

NOR2x1p5_ASAP7_75t_R c5800(
.A(net5784),
.B(net5703),
.Y(net5853)
);

AOI22xp5_ASAP7_75t_R c5801(
.A1(net5808),
.A2(net5843),
.B1(net5853),
.B2(net5846),
.Y(net5854)
);

OR5x1_ASAP7_75t_R c5802(
.A(net5734),
.B(net3015),
.C(net4911),
.D(net5779),
.E(net5853),
.Y(net5855)
);

NOR3x2_ASAP7_75t_R c5803(
.B(net5809),
.C(net5797),
.A(net10020),
.Y(net5856)
);

BUFx6f_ASAP7_75t_R c5804(
.A(net10557),
.Y(net5857)
);

NOR3xp33_ASAP7_75t_R c5805(
.A(net5745),
.B(net5857),
.C(net10145),
.Y(net5858)
);

NOR2x2_ASAP7_75t_R c5806(
.A(net5856),
.B(net5846),
.Y(net5859)
);

NOR2xp33_ASAP7_75t_R c5807(
.A(net4835),
.B(net10145),
.Y(net5860)
);

OR5x2_ASAP7_75t_R c5808(
.A(net5830),
.B(net5804),
.C(net5853),
.D(net3079),
.E(net3015),
.Y(net5861)
);

A2O1A1O1Ixp25_ASAP7_75t_R c5809(
.A1(net5842),
.A2(net4843),
.B(net5853),
.C(net3977),
.D(net9826),
.Y(net5862)
);

NOR2xp67_ASAP7_75t_R c5810(
.A(net4058),
.B(net4867),
.Y(net5863)
);

OR2x2_ASAP7_75t_R c5811(
.A(net5697),
.B(net10161),
.Y(net5864)
);

BUFx8_ASAP7_75t_R c5812(
.A(net4732),
.Y(net5865)
);

OA21x2_ASAP7_75t_R c5813(
.A1(net4920),
.A2(net5006),
.B(net5846),
.Y(net5866)
);

OR2x4_ASAP7_75t_R c5814(
.A(net5609),
.B(net5000),
.Y(net5867)
);

OR2x6_ASAP7_75t_R c5815(
.A(net5613),
.B(net4954),
.Y(net5868)
);

CKINVDCx10_ASAP7_75t_R c5816(
.A(net5721),
.Y(net5869)
);

OAI21x1_ASAP7_75t_R c5817(
.A1(net4746),
.A2(net5831),
.B(net5747),
.Y(net5870)
);

XNOR2x1_ASAP7_75t_R c5818(
.B(net5865),
.A(net4971),
.Y(net5871)
);

CKINVDCx11_ASAP7_75t_R c5819(
.A(net10120),
.Y(net5872)
);

CKINVDCx12_ASAP7_75t_R c5820(
.A(net10329),
.Y(net5873)
);

OAI21xp33_ASAP7_75t_R c5821(
.A1(net4867),
.A2(net4870),
.B(net4963),
.Y(net5874)
);

CKINVDCx14_ASAP7_75t_R c5822(
.A(net10329),
.Y(net5875)
);

CKINVDCx16_ASAP7_75t_R c5823(
.A(net10168),
.Y(net5876)
);

XNOR2x2_ASAP7_75t_R c5824(
.A(net3079),
.B(net5645),
.Y(net5877)
);

CKINVDCx20_ASAP7_75t_R c5825(
.A(net5000),
.Y(net5878)
);

CKINVDCx5p33_ASAP7_75t_R c5826(
.A(net5813),
.Y(net5879)
);

XNOR2xp5_ASAP7_75t_R c5827(
.A(net5873),
.B(net4957),
.Y(net5880)
);

CKINVDCx6p67_ASAP7_75t_R c5828(
.A(net5863),
.Y(net5881)
);

CKINVDCx8_ASAP7_75t_R c5829(
.A(net10471),
.Y(net5882)
);

XOR2x1_ASAP7_75t_R c5830(
.A(net4954),
.B(net5721),
.Y(net5883)
);

ICGx4_ASAP7_75t_R c5831(
.ENA(net5815),
.SE(net5004),
.CLK(clk),
.GCLK(net5884)
);

CKINVDCx9p33_ASAP7_75t_R c5832(
.A(net5790),
.Y(net5885)
);

HB1xp67_ASAP7_75t_R c5833(
.A(net10531),
.Y(net5886)
);

HB2xp67_ASAP7_75t_R c5834(
.A(net9977),
.Y(net5887)
);

HB3xp67_ASAP7_75t_R c5835(
.A(net5818),
.Y(net5888)
);

HB4xp67_ASAP7_75t_R c5836(
.A(net4863),
.Y(net5889)
);

INVx11_ASAP7_75t_R c5837(
.A(net9948),
.Y(net5890)
);

XOR2x2_ASAP7_75t_R c5838(
.A(net5701),
.B(net5884),
.Y(net5891)
);

XOR2xp5_ASAP7_75t_R c5839(
.A(net5864),
.B(net5885),
.Y(net5892)
);

AND2x2_ASAP7_75t_R c5840(
.A(net5629),
.B(net5879),
.Y(net5893)
);

INVx13_ASAP7_75t_R c5841(
.A(net10555),
.Y(net5894)
);

AND2x4_ASAP7_75t_R c5842(
.A(net4964),
.B(net2034),
.Y(net5895)
);

AND2x6_ASAP7_75t_R c5843(
.A(net5860),
.B(net5892),
.Y(net5896)
);

HAxp5_ASAP7_75t_R c5844(
.A(net5871),
.B(net5896),
.CON(net5898),
.SN(net5897)
);

NAND2x1_ASAP7_75t_R c5845(
.A(net3936),
.B(net5786),
.Y(net5899)
);

NAND2x1p5_ASAP7_75t_R c5846(
.A(net4947),
.B(net5609),
.Y(net5900)
);

NAND2x2_ASAP7_75t_R c5847(
.A(net4996),
.B(net5824),
.Y(net5901)
);

NAND2xp33_ASAP7_75t_R c5848(
.A(net3079),
.B(net10240),
.Y(net5902)
);

NAND2xp5_ASAP7_75t_R c5849(
.A(net5863),
.B(net10224),
.Y(net5903)
);

NAND2xp67_ASAP7_75t_R c5850(
.A(net5827),
.B(net4911),
.Y(net5904)
);

NOR2x1_ASAP7_75t_R c5851(
.A(net3977),
.B(net4863),
.Y(net5905)
);

DFFASRHQNx1_ASAP7_75t_R c5852(
.D(net5870),
.RESETN(net5887),
.SETN(net5902),
.CLK(clk),
.QN(net5906)
);

NOR2x1p5_ASAP7_75t_R c5853(
.A(net5899),
.B(net5813),
.Y(net5907)
);

OAI21xp5_ASAP7_75t_R c5854(
.A1(net5874),
.A2(net5869),
.B(net5899),
.Y(net5908)
);

NOR2x2_ASAP7_75t_R c5855(
.A(net5878),
.B(net5899),
.Y(net5909)
);

OR3x1_ASAP7_75t_R c5856(
.A(net5875),
.B(net5903),
.C(net5905),
.Y(net5910)
);

NOR2xp33_ASAP7_75t_R c5857(
.A(net5877),
.B(net5905),
.Y(net5911)
);

INVx1_ASAP7_75t_R c5858(
.A(net10499),
.Y(net5912)
);

NOR2xp67_ASAP7_75t_R c5859(
.A(net5876),
.B(net5906),
.Y(net5913)
);

INVx2_ASAP7_75t_R c5860(
.A(net5703),
.Y(net5914)
);

INVx3_ASAP7_75t_R c5861(
.A(net5885),
.Y(net5915)
);

OR2x2_ASAP7_75t_R c5862(
.A(net5895),
.B(net5894),
.Y(net5916)
);

OR2x4_ASAP7_75t_R c5863(
.A(net3988),
.B(net5846),
.Y(net5917)
);

OR3x2_ASAP7_75t_R c5864(
.A(net5917),
.B(net5023),
.C(net5893),
.Y(net5918)
);

OR2x6_ASAP7_75t_R c5865(
.A(net5890),
.B(net5865),
.Y(net5919)
);

SDFHx1_ASAP7_75t_R c5866(
.D(net5916),
.SE(net5883),
.SI(net5910),
.CLK(clk),
.QN(net5920)
);

XNOR2x1_ASAP7_75t_R c5867(
.B(net5915),
.A(net5909),
.Y(net5921)
);

XNOR2x2_ASAP7_75t_R c5868(
.A(net5892),
.B(net3977),
.Y(net5922)
);

XNOR2xp5_ASAP7_75t_R c5869(
.A(net5896),
.B(net5884),
.Y(net5923)
);

OR3x4_ASAP7_75t_R c5870(
.A(net5859),
.B(net5921),
.C(net5890),
.Y(net5924)
);

AND3x1_ASAP7_75t_R c5871(
.A(net5869),
.B(net5906),
.C(net5015),
.Y(net5925)
);

AND3x2_ASAP7_75t_R c5872(
.A(net5902),
.B(net5920),
.C(net5911),
.Y(net5926)
);

XOR2x1_ASAP7_75t_R c5873(
.A(net5881),
.B(net5919),
.Y(net5927)
);

AND3x4_ASAP7_75t_R c5874(
.A(net5912),
.B(net5898),
.C(net5886),
.Y(net5928)
);

AO21x1_ASAP7_75t_R c5875(
.A1(net5911),
.A2(net5915),
.B(net4064),
.Y(net5929)
);

AO21x2_ASAP7_75t_R c5876(
.A1(net5919),
.A2(net5889),
.B(net5928),
.Y(net5930)
);

AOI21x1_ASAP7_75t_R c5877(
.A1(net5914),
.A2(net5906),
.B(net5876),
.Y(net5931)
);

AOI21xp33_ASAP7_75t_R c5878(
.A1(net5791),
.A2(net5931),
.B(net5915),
.Y(net5932)
);

INVx4_ASAP7_75t_R c5879(
.A(net10170),
.Y(net5933)
);

AOI21xp5_ASAP7_75t_R c5880(
.A1(net3939),
.A2(net5906),
.B(net5015),
.Y(net5934)
);

FAx1_ASAP7_75t_R c5881(
.A(net5927),
.B(net5829),
.CI(net10032),
.SN(net5936),
.CON(net5935)
);

MAJIxp5_ASAP7_75t_R c5882(
.A(net5905),
.B(net5935),
.C(net9977),
.Y(net5937)
);

XOR2x2_ASAP7_75t_R c5883(
.A(net5923),
.B(net5903),
.Y(net5938)
);

AND5x1_ASAP7_75t_R c5884(
.A(net5829),
.B(net5929),
.C(net5934),
.D(net5938),
.E(net5769),
.Y(net5939)
);

SDFHx2_ASAP7_75t_R c5885(
.D(net3846),
.SE(net5921),
.SI(net5932),
.CLK(clk),
.QN(net5940)
);

MAJx2_ASAP7_75t_R c5886(
.A(net5913),
.B(net5923),
.C(net10070),
.Y(net5941)
);

MAJx3_ASAP7_75t_R c5887(
.A(net4840),
.B(net5936),
.C(net5938),
.Y(net5942)
);

NAND3x1_ASAP7_75t_R c5888(
.A(net5937),
.B(net5910),
.C(net5933),
.Y(net5943)
);

NAND3x2_ASAP7_75t_R c5889(
.B(net3955),
.C(net5943),
.A(net5934),
.Y(net5944)
);

NAND3xp33_ASAP7_75t_R c5890(
.A(net5941),
.B(net5942),
.C(net5934),
.Y(net5945)
);

AND5x2_ASAP7_75t_R c5891(
.A(net4939),
.B(net5933),
.C(net4954),
.D(net5945),
.E(net5928),
.Y(net5946)
);

NOR3x1_ASAP7_75t_R c5892(
.A(net5945),
.B(net10013),
.C(net10270),
.Y(net5947)
);

INVx5_ASAP7_75t_R c5893(
.A(net10070),
.Y(net5948)
);

XOR2xp5_ASAP7_75t_R c5894(
.A(net5831),
.B(net1348),
.Y(net5949)
);

INVx6_ASAP7_75t_R c5895(
.A(net1337),
.Y(net5950)
);

INVx8_ASAP7_75t_R c5896(
.A(net9227),
.Y(net5951)
);

INVxp33_ASAP7_75t_R c5897(
.A(net9188),
.Y(net5952)
);

INVxp67_ASAP7_75t_R c5898(
.A(net5015),
.Y(net5953)
);

BUFx10_ASAP7_75t_R c5899(
.A(net5889),
.Y(net5954)
);

AND2x2_ASAP7_75t_R c5900(
.A(net5038),
.B(net5929),
.Y(net5955)
);

NOR3x2_ASAP7_75t_R c5901(
.B(net5951),
.C(net5894),
.A(net5900),
.Y(net5956)
);

SDFHx3_ASAP7_75t_R c5902(
.D(net5953),
.SE(net5843),
.SI(net5949),
.CLK(clk),
.QN(net5957)
);

BUFx12_ASAP7_75t_R c5903(
.A(net5938),
.Y(net5958)
);

AND2x4_ASAP7_75t_R c5904(
.A(net5094),
.B(net5769),
.Y(net5959)
);

AND2x6_ASAP7_75t_R c5905(
.A(net5938),
.B(net9811),
.Y(net5960)
);

BUFx12f_ASAP7_75t_R c5906(
.A(net5023),
.Y(net5961)
);

NOR3xp33_ASAP7_75t_R c5907(
.A(net5085),
.B(net4099),
.C(net4148),
.Y(net5962)
);

BUFx16f_ASAP7_75t_R c5908(
.A(net9188),
.Y(net5963)
);

ICGx5_ASAP7_75t_R c5909(
.ENA(net5880),
.SE(net5963),
.CLK(clk),
.GCLK(net5964)
);

BUFx24_ASAP7_75t_R c5910(
.A(net10127),
.Y(net5965)
);

BUFx2_ASAP7_75t_R c5911(
.A(net9208),
.Y(net5966)
);

HAxp5_ASAP7_75t_R c5912(
.A(net5963),
.B(net1196),
.CON(net5967)
);

BUFx3_ASAP7_75t_R c5913(
.A(net10465),
.Y(net5968)
);

BUFx4_ASAP7_75t_R c5914(
.A(net5033),
.Y(net5969)
);

BUFx4f_ASAP7_75t_R c5915(
.A(net5584),
.Y(net5970)
);

ICGx5p33DC_ASAP7_75t_R c5916(
.ENA(net5101),
.SE(net5959),
.CLK(clk),
.GCLK(net5971)
);

BUFx5_ASAP7_75t_R c5917(
.A(net5901),
.Y(net5972)
);

NAND2x1_ASAP7_75t_R c5918(
.A(net5036),
.B(net10127),
.Y(net5973)
);

NAND2x1p5_ASAP7_75t_R c5919(
.A(net4924),
.B(net5948),
.Y(net5974)
);

NAND2x2_ASAP7_75t_R c5920(
.A(net5965),
.B(net5889),
.Y(net5975)
);

BUFx6f_ASAP7_75t_R c5921(
.A(net9241),
.Y(net5976)
);

NAND2xp33_ASAP7_75t_R c5922(
.A(net5952),
.B(net5030),
.Y(net5977)
);

OA21x2_ASAP7_75t_R c5923(
.A1(net5966),
.A2(net5033),
.B(net5769),
.Y(net5978)
);

OAI21x1_ASAP7_75t_R c5924(
.A1(net5975),
.A2(net5951),
.B(net5971),
.Y(net5979)
);

ICGx6p67DC_ASAP7_75t_R c5925(
.ENA(net5004),
.SE(net5964),
.CLK(clk),
.GCLK(net5980)
);

NAND2xp5_ASAP7_75t_R c5926(
.A(net5012),
.B(net5833),
.Y(net5981)
);

NAND2xp67_ASAP7_75t_R c5927(
.A(net5964),
.B(net9690),
.Y(net5982)
);

NOR2x1_ASAP7_75t_R c5928(
.A(net5954),
.B(net5962),
.Y(net5983)
);

BUFx8_ASAP7_75t_R c5929(
.A(net4121),
.Y(net5984)
);

NOR2x1p5_ASAP7_75t_R c5930(
.A(net4148),
.B(net5982),
.Y(net5985)
);

ICGx8DC_ASAP7_75t_R c5931(
.ENA(net5955),
.SE(net5948),
.CLK(clk),
.GCLK(net5986)
);

NOR2x2_ASAP7_75t_R c5932(
.A(net5093),
.B(net3987),
.Y(net5987)
);

NOR2xp33_ASAP7_75t_R c5933(
.A(net5962),
.B(net4174),
.Y(net5988)
);

AOI31xp33_ASAP7_75t_R c5934(
.A1(net5970),
.A2(net5971),
.A3(net5087),
.B(net5929),
.Y(net5989)
);

AOI31xp67_ASAP7_75t_R c5935(
.A1(net5969),
.A2(net5975),
.A3(net5938),
.B(net5960),
.Y(net5990)
);

NOR2xp67_ASAP7_75t_R c5936(
.A(net3086),
.B(net5952),
.Y(net5991)
);

CKINVDCx10_ASAP7_75t_R c5937(
.A(net10441),
.Y(net5992)
);

OR2x2_ASAP7_75t_R c5938(
.A(net5957),
.B(net9690),
.Y(net5993)
);

OR2x4_ASAP7_75t_R c5939(
.A(net4128),
.B(net5948),
.Y(net5994)
);

CKINVDCx11_ASAP7_75t_R c5940(
.A(net5993),
.Y(net5995)
);

OAI21xp33_ASAP7_75t_R c5941(
.A1(net5951),
.A2(net5036),
.B(net10036),
.Y(net5996)
);

OR2x6_ASAP7_75t_R c5942(
.A(net5974),
.B(net4985),
.Y(net5997)
);

CKINVDCx12_ASAP7_75t_R c5943(
.A(net10166),
.Y(net5998)
);

XNOR2x1_ASAP7_75t_R c5944(
.B(net5981),
.A(net4962),
.Y(net5999)
);

XNOR2x2_ASAP7_75t_R c5945(
.A(net5972),
.B(net5982),
.Y(net6000)
);

CKINVDCx14_ASAP7_75t_R c5946(
.A(net10544),
.Y(net6001)
);

XNOR2xp5_ASAP7_75t_R c5947(
.A(net5976),
.B(net6000),
.Y(net6002)
);

XOR2x1_ASAP7_75t_R c5948(
.A(net5985),
.B(net5969),
.Y(net6003)
);

XOR2x2_ASAP7_75t_R c5949(
.A(net5961),
.B(net6003),
.Y(net6004)
);

XOR2xp5_ASAP7_75t_R c5950(
.A(net5044),
.B(net5833),
.Y(net6005)
);

ICGx1_ASAP7_75t_R c5951(
.ENA(net4140),
.SE(net5945),
.CLK(clk),
.GCLK(net6006)
);

AND2x2_ASAP7_75t_R c5952(
.A(net6005),
.B(net5975),
.Y(net6007)
);

AND2x4_ASAP7_75t_R c5953(
.A(net5100),
.B(net5986),
.Y(net6008)
);

AND2x6_ASAP7_75t_R c5954(
.A(net5995),
.B(net6006),
.Y(net6009)
);

AO221x1_ASAP7_75t_R c5955(
.A1(net6000),
.A2(net5786),
.B1(net5094),
.B2(net6007),
.C(net5077),
.Y(net6010)
);

NAND4xp25_ASAP7_75t_R c5956(
.A(net5894),
.B(net6006),
.C(net6007),
.D(net6010),
.Y(net6011)
);

CKINVDCx16_ASAP7_75t_R c5957(
.A(net6007),
.Y(net6012)
);

OAI21xp5_ASAP7_75t_R c5958(
.A1(net5958),
.A2(net6006),
.B(net5968),
.Y(net6013)
);

HAxp5_ASAP7_75t_R c5959(
.A(net6006),
.B(net5954),
.CON(net6014)
);

NAND2x1_ASAP7_75t_R c5960(
.A(net4116),
.B(net6002),
.Y(net6015)
);

NAND2x1p5_ASAP7_75t_R c5961(
.A(net6014),
.B(net5984),
.Y(net6016)
);

AOI321xp33_ASAP7_75t_R c5962(
.A1(net4125),
.A2(net5980),
.A3(net6010),
.B1(net5033),
.B2(net5105),
.C(net5996),
.Y(net6017)
);

NAND4xp75_ASAP7_75t_R c5963(
.A(net5631),
.B(net4177),
.C(net5974),
.D(net5833),
.Y(net6018)
);

NAND2x2_ASAP7_75t_R c5964(
.A(net4959),
.B(net5971),
.Y(net6019)
);

OR3x1_ASAP7_75t_R c5965(
.A(net5990),
.B(net5974),
.C(net6007),
.Y(net6020)
);

OR3x2_ASAP7_75t_R c5966(
.A(net6001),
.B(net6018),
.C(net6016),
.Y(net6021)
);

NOR4xp25_ASAP7_75t_R c5967(
.A(net6012),
.B(net5969),
.C(net6010),
.D(net5076),
.Y(net6022)
);

OR3x4_ASAP7_75t_R c5968(
.A(net6011),
.B(net6020),
.C(net5085),
.Y(net6023)
);

NAND2xp33_ASAP7_75t_R c5969(
.A(net5988),
.B(net10147),
.Y(net6024)
);

NAND2xp5_ASAP7_75t_R c5970(
.A(net6015),
.B(net6002),
.Y(net6025)
);

AND3x1_ASAP7_75t_R c5971(
.A(net6013),
.B(net6024),
.C(net9916),
.Y(net6026)
);

NAND2xp67_ASAP7_75t_R c5972(
.A(net5948),
.B(net6025),
.Y(net6027)
);

AND3x2_ASAP7_75t_R c5973(
.A(net6021),
.B(net6003),
.C(net6020),
.Y(net6028)
);

AND3x4_ASAP7_75t_R c5974(
.A(net6024),
.B(net6009),
.C(net6018),
.Y(net6029)
);

AO221x2_ASAP7_75t_R c5975(
.A1(net6010),
.A2(net3253),
.B1(net6029),
.B2(net5932),
.C(net10101),
.Y(net6030)
);

NOR2x1_ASAP7_75t_R c5976(
.A(net4897),
.B(net6013),
.Y(net6031)
);

CKINVDCx20_ASAP7_75t_R c5977(
.A(net10380),
.Y(net6032)
);

CKINVDCx5p33_ASAP7_75t_R c5978(
.A(net5979),
.Y(net6033)
);

CKINVDCx6p67_ASAP7_75t_R c5979(
.A(net9117),
.Y(net6034)
);

NOR2x1p5_ASAP7_75t_R c5980(
.A(net5124),
.B(net5964),
.Y(net6035)
);

NOR2x2_ASAP7_75t_R c5981(
.A(net5998),
.B(net5986),
.Y(net6036)
);

NOR2xp33_ASAP7_75t_R c5982(
.A(net6002),
.B(net5949),
.Y(net6037)
);

CKINVDCx8_ASAP7_75t_R c5983(
.A(net5949),
.Y(net6038)
);

NOR2xp67_ASAP7_75t_R c5984(
.A(net5076),
.B(net9884),
.Y(net6039)
);

CKINVDCx9p33_ASAP7_75t_R c5985(
.A(net10450),
.Y(net6040)
);

HB1xp67_ASAP7_75t_R c5986(
.A(net6037),
.Y(net6041)
);

HB2xp67_ASAP7_75t_R c5987(
.A(net5134),
.Y(net6042)
);

OR2x2_ASAP7_75t_R c5988(
.A(net5950),
.B(net5111),
.Y(net6043)
);

HB3xp67_ASAP7_75t_R c5989(
.A(net5185),
.Y(net6044)
);

HB4xp67_ASAP7_75t_R c5990(
.A(net6035),
.Y(net6045)
);

OR2x4_ASAP7_75t_R c5991(
.A(net5980),
.B(net6013),
.Y(net6046)
);

AO21x1_ASAP7_75t_R c5992(
.A1(net6010),
.A2(net6044),
.B(net10256),
.Y(net6047)
);

OR2x6_ASAP7_75t_R c5993(
.A(net5165),
.B(net6036),
.Y(net6048)
);

INVx11_ASAP7_75t_R c5994(
.A(net6034),
.Y(net6049)
);

XNOR2x1_ASAP7_75t_R c5995(
.B(net5645),
.A(net5059),
.Y(net6050)
);

XNOR2x2_ASAP7_75t_R c5996(
.A(net5113),
.B(net5824),
.Y(net6051)
);

XNOR2xp5_ASAP7_75t_R c5997(
.A(net5127),
.B(net5929),
.Y(net6052)
);

INVx13_ASAP7_75t_R c5998(
.A(net5929),
.Y(net6053)
);

AO21x2_ASAP7_75t_R c5999(
.A1(net6013),
.A2(net5996),
.B(net4962),
.Y(net6054)
);

INVx1_ASAP7_75t_R c6000(
.A(net5191),
.Y(net6055)
);

SDFHx4_ASAP7_75t_R c6001(
.D(net5647),
.SE(net6055),
.SI(net5130),
.CLK(clk),
.QN(net6056)
);

XOR2x1_ASAP7_75t_R c6002(
.A(net6043),
.B(net5047),
.Y(net6057)
);

INVx2_ASAP7_75t_R c6003(
.A(net10506),
.Y(net6058)
);

XOR2x2_ASAP7_75t_R c6004(
.A(net4195),
.B(net6045),
.Y(net6059)
);

XOR2xp5_ASAP7_75t_R c6005(
.A(net2381),
.B(net4222),
.Y(net6060)
);

INVx3_ASAP7_75t_R c6006(
.A(net9117),
.Y(net6061)
);

AND2x2_ASAP7_75t_R c6007(
.A(net5986),
.B(net5135),
.Y(net6062)
);

AND2x4_ASAP7_75t_R c6008(
.A(net6036),
.B(net6045),
.Y(net6063)
);

AND2x6_ASAP7_75t_R c6009(
.A(net6029),
.B(net4185),
.Y(net6064)
);

INVx4_ASAP7_75t_R c6010(
.A(net9802),
.Y(net6065)
);

INVx5_ASAP7_75t_R c6011(
.A(net10537),
.Y(net6066)
);

HAxp5_ASAP7_75t_R c6012(
.A(net5824),
.B(net6064),
.CON(net6068),
.SN(net6067)
);

INVx6_ASAP7_75t_R c6013(
.A(net6062),
.Y(net6069)
);

NAND2x1_ASAP7_75t_R c6014(
.A(net6061),
.B(net4195),
.Y(net6070)
);

NAND2x1p5_ASAP7_75t_R c6015(
.A(net6032),
.B(net5645),
.Y(net6071)
);

NAND2x2_ASAP7_75t_R c6016(
.A(net6063),
.B(net10270),
.Y(net6072)
);

NOR4xp75_ASAP7_75t_R c6017(
.A(net6038),
.B(net4953),
.C(net4960),
.D(net5968),
.Y(net6073)
);

NAND2xp33_ASAP7_75t_R c6018(
.A(net4249),
.B(net6029),
.Y(net6074)
);

NAND2xp5_ASAP7_75t_R c6019(
.A(net6004),
.B(net6010),
.Y(net6075)
);

NAND2xp67_ASAP7_75t_R c6020(
.A(net6070),
.B(net5047),
.Y(net6076)
);

NOR2x1_ASAP7_75t_R c6021(
.A(net5706),
.B(net6072),
.Y(net6077)
);

AOI21x1_ASAP7_75t_R c6022(
.A1(net5059),
.A2(net5121),
.B(net5191),
.Y(net6078)
);

INVx8_ASAP7_75t_R c6023(
.A(net10413),
.Y(net6079)
);

AOI21xp33_ASAP7_75t_R c6024(
.A1(net5164),
.A2(net6067),
.B(net5888),
.Y(net6080)
);

NOR2x1p5_ASAP7_75t_R c6025(
.A(net6061),
.B(net9936),
.Y(net6081)
);

NOR2x2_ASAP7_75t_R c6026(
.A(net5059),
.B(net9802),
.Y(net6082)
);

NOR2xp33_ASAP7_75t_R c6027(
.A(net6069),
.B(net9678),
.Y(net6083)
);

NOR2xp67_ASAP7_75t_R c6028(
.A(net5145),
.B(net6029),
.Y(net6084)
);

OR2x2_ASAP7_75t_R c6029(
.A(net5171),
.B(net6058),
.Y(net6085)
);

AOI21xp5_ASAP7_75t_R c6030(
.A1(net6068),
.A2(net6079),
.B(net6056),
.Y(net6086)
);

INVxp33_ASAP7_75t_R c6031(
.A(net10156),
.Y(net6087)
);

OR2x4_ASAP7_75t_R c6032(
.A(net6084),
.B(net5908),
.Y(net6088)
);

INVxp67_ASAP7_75t_R c6033(
.A(net10477),
.Y(net6089)
);

OR2x6_ASAP7_75t_R c6034(
.A(net6083),
.B(net4257),
.Y(net6090)
);

XNOR2x1_ASAP7_75t_R c6035(
.B(net5588),
.A(net5111),
.Y(net6091)
);

O2A1O1Ixp33_ASAP7_75t_R c6036(
.A1(net5888),
.A2(net6087),
.B(net5706),
.C(net4962),
.Y(net6092)
);

FAx1_ASAP7_75t_R c6037(
.A(net4222),
.B(net6082),
.CI(net6087),
.SN(net6094),
.CON(net6093)
);

XNOR2x2_ASAP7_75t_R c6038(
.A(net6030),
.B(net5185),
.Y(net6095)
);

XNOR2xp5_ASAP7_75t_R c6039(
.A(net6059),
.B(net6087),
.Y(net6096)
);

XOR2x1_ASAP7_75t_R c6040(
.A(net6047),
.B(net6038),
.Y(net6097)
);

XOR2x2_ASAP7_75t_R c6041(
.A(net6089),
.B(net6093),
.Y(net6098)
);

XOR2xp5_ASAP7_75t_R c6042(
.A(net5143),
.B(net5978),
.Y(net6099)
);

BUFx10_ASAP7_75t_R c6043(
.A(net10020),
.Y(net6100)
);

MAJIxp5_ASAP7_75t_R c6044(
.A(net6079),
.B(net6094),
.C(net6085),
.Y(net6101)
);

AND2x2_ASAP7_75t_R c6045(
.A(net6081),
.B(net6098),
.Y(net6102)
);

MAJx2_ASAP7_75t_R c6046(
.A(net6056),
.B(net5134),
.C(net6099),
.Y(net6103)
);

BUFx12_ASAP7_75t_R c6047(
.A(net10524),
.Y(net6104)
);

AO32x1_ASAP7_75t_R c6048(
.A1(net6091),
.A2(net6098),
.A3(net6102),
.B1(net6058),
.B2(net6099),
.Y(net6105)
);

AND2x4_ASAP7_75t_R c6049(
.A(net6090),
.B(net10271),
.Y(net6106)
);

AND2x6_ASAP7_75t_R c6050(
.A(net6078),
.B(net6094),
.Y(net6107)
);

AO32x2_ASAP7_75t_R c6051(
.A1(net6074),
.A2(net5165),
.A3(net6091),
.B1(net6087),
.B2(net6102),
.Y(net6108)
);

SDFLx1_ASAP7_75t_R c6052(
.D(net6108),
.SE(net6074),
.SI(net6102),
.CLK(clk),
.QN(net6109)
);

HAxp5_ASAP7_75t_R c6053(
.A(net6098),
.B(net6078),
.CON(net6110)
);

AOI221x1_ASAP7_75t_R c6054(
.A1(net6064),
.A2(net6100),
.B1(net6096),
.B2(net6109),
.C(net5996),
.Y(net6111)
);

NAND2x1_ASAP7_75t_R c6055(
.A(net6095),
.B(net6109),
.Y(net6112)
);

NAND2x1p5_ASAP7_75t_R c6056(
.A(net6106),
.B(net6059),
.Y(net6113)
);

BUFx12f_ASAP7_75t_R c6057(
.A(net10366),
.Y(net6114)
);

AOI221xp5_ASAP7_75t_R c6058(
.A1(net6086),
.A2(net6114),
.B1(net6040),
.B2(net6104),
.C(net5135),
.Y(net6115)
);

BUFx16f_ASAP7_75t_R c6059(
.A(net10448),
.Y(net6116)
);

BUFx24_ASAP7_75t_R c6060(
.A(net6107),
.Y(net6117)
);

BUFx2_ASAP7_75t_R c6061(
.A(net6042),
.Y(net6118)
);

NAND2x2_ASAP7_75t_R c6062(
.A(net5172),
.B(net5097),
.Y(net6119)
);

MAJx3_ASAP7_75t_R c6063(
.A(net4229),
.B(net5260),
.C(net9656),
.Y(net6120)
);

BUFx3_ASAP7_75t_R c6064(
.A(net9157),
.Y(net6121)
);

NAND2xp33_ASAP7_75t_R c6065(
.A(net5047),
.B(net5252),
.Y(net6122)
);

BUFx4_ASAP7_75t_R c6066(
.A(net3269),
.Y(net6123)
);

BUFx4f_ASAP7_75t_R c6067(
.A(net10502),
.Y(net6124)
);

NAND2xp5_ASAP7_75t_R c6068(
.A(net5934),
.B(net6100),
.Y(net6125)
);

NAND3x1_ASAP7_75t_R c6069(
.A(net6117),
.B(net6125),
.C(net6124),
.Y(net6126)
);

NAND2xp67_ASAP7_75t_R c6070(
.A(net4308),
.B(net4957),
.Y(net6127)
);

BUFx5_ASAP7_75t_R c6071(
.A(net3416),
.Y(net6128)
);

NOR2x1_ASAP7_75t_R c6072(
.A(net5223),
.B(net5211),
.Y(net6129)
);

BUFx6f_ASAP7_75t_R c6073(
.A(net6116),
.Y(net6130)
);

NAND3x2_ASAP7_75t_R c6074(
.B(net5242),
.C(net4329),
.A(net6123),
.Y(net6131)
);

BUFx8_ASAP7_75t_R c6075(
.A(net4960),
.Y(net6132)
);

CKINVDCx10_ASAP7_75t_R c6076(
.A(net10514),
.Y(net6133)
);

CKINVDCx11_ASAP7_75t_R c6077(
.A(net10443),
.Y(net6134)
);

NOR2x1p5_ASAP7_75t_R c6078(
.A(net6100),
.B(net6122),
.Y(net6135)
);

CKINVDCx12_ASAP7_75t_R c6079(
.A(net6041),
.Y(net6136)
);

NOR2x2_ASAP7_75t_R c6080(
.A(net6051),
.B(net6058),
.Y(net6137)
);

NOR2xp33_ASAP7_75t_R c6081(
.A(net6137),
.B(net5168),
.Y(net6138)
);

NOR2xp67_ASAP7_75t_R c6082(
.A(net6110),
.B(net6080),
.Y(net6139)
);

CKINVDCx14_ASAP7_75t_R c6083(
.A(net10468),
.Y(net6140)
);

CKINVDCx16_ASAP7_75t_R c6084(
.A(net6133),
.Y(net6141)
);

CKINVDCx20_ASAP7_75t_R c6085(
.A(net10540),
.Y(net6142)
);

CKINVDCx5p33_ASAP7_75t_R c6086(
.A(net9157),
.Y(net6143)
);

NAND3xp33_ASAP7_75t_R c6087(
.A(net4229),
.B(net6131),
.C(net4166),
.Y(net6144)
);

OR2x2_ASAP7_75t_R c6088(
.A(net5252),
.B(net4214),
.Y(net6145)
);

OR2x4_ASAP7_75t_R c6089(
.A(net6134),
.B(net6129),
.Y(net6146)
);

OR2x6_ASAP7_75t_R c6090(
.A(net6145),
.B(net10256),
.Y(net6147)
);

XNOR2x1_ASAP7_75t_R c6091(
.B(net5213),
.A(net6145),
.Y(net6148)
);

NOR3x1_ASAP7_75t_R c6092(
.A(net5251),
.B(net6119),
.C(net5218),
.Y(net6149)
);

CKINVDCx6p67_ASAP7_75t_R c6093(
.A(net10525),
.Y(net6150)
);

XNOR2x2_ASAP7_75t_R c6094(
.A(net6135),
.B(net6146),
.Y(net6151)
);

XNOR2xp5_ASAP7_75t_R c6095(
.A(net6118),
.B(net5898),
.Y(net6152)
);

XOR2x1_ASAP7_75t_R c6096(
.A(net6145),
.B(net6085),
.Y(net6153)
);

SDFLx2_ASAP7_75t_R c6097(
.D(net6082),
.SE(net6150),
.SI(net6144),
.CLK(clk),
.QN(net6154)
);

XOR2x2_ASAP7_75t_R c6098(
.A(net1526),
.B(net10104),
.Y(net6155)
);

CKINVDCx8_ASAP7_75t_R c6099(
.A(net10104),
.Y(net6156)
);

XOR2xp5_ASAP7_75t_R c6100(
.A(net6143),
.B(net5097),
.Y(net6157)
);

CKINVDCx9p33_ASAP7_75t_R c6101(
.A(net10442),
.Y(net6158)
);

AND2x2_ASAP7_75t_R c6102(
.A(net6155),
.B(net4957),
.Y(net6159)
);

AND2x4_ASAP7_75t_R c6103(
.A(net5218),
.B(net6155),
.Y(net6160)
);

AND2x6_ASAP7_75t_R c6104(
.A(net6065),
.B(net5147),
.Y(net6161)
);

NOR3x2_ASAP7_75t_R c6105(
.B(net5999),
.C(net6145),
.A(net9918),
.Y(net6162)
);

SDFLx3_ASAP7_75t_R c6106(
.D(net5217),
.SE(net6143),
.SI(net6159),
.CLK(clk),
.QN(net6163)
);

HAxp5_ASAP7_75t_R c6107(
.A(net6147),
.B(net9722),
.CON(net6165),
.SN(net6164)
);

NAND2x1_ASAP7_75t_R c6108(
.A(net6130),
.B(net10104),
.Y(net6166)
);

NAND2x1p5_ASAP7_75t_R c6109(
.A(net2498),
.B(net6166),
.Y(net6167)
);

NAND2x2_ASAP7_75t_R c6110(
.A(net4339),
.B(net6153),
.Y(net6168)
);

NAND2xp33_ASAP7_75t_R c6111(
.A(net6166),
.B(net9811),
.Y(net6169)
);

NAND2xp5_ASAP7_75t_R c6112(
.A(net6130),
.B(net5172),
.Y(net6170)
);

NAND2xp67_ASAP7_75t_R c6113(
.A(net6160),
.B(net6142),
.Y(net6171)
);

HB1xp67_ASAP7_75t_R c6114(
.A(net10452),
.Y(net6172)
);

NOR2x1_ASAP7_75t_R c6115(
.A(net6161),
.B(net6169),
.Y(net6173)
);

NOR2x1p5_ASAP7_75t_R c6116(
.A(net2452),
.B(net6107),
.Y(net6174)
);

NOR3xp33_ASAP7_75t_R c6117(
.A(net6170),
.B(net5223),
.C(net5833),
.Y(net6175)
);

AOI33xp33_ASAP7_75t_R c6118(
.A1(net6162),
.A2(net5833),
.A3(net6135),
.B1(net5135),
.B2(net6146),
.B3(net10256),
.Y(net6176)
);

NOR2x2_ASAP7_75t_R c6119(
.A(net6150),
.B(net6134),
.Y(net6177)
);

SDFLx4_ASAP7_75t_R c6120(
.D(net6171),
.SE(net6119),
.SI(net5225),
.CLK(clk),
.QN(net6178)
);

O2A1O1Ixp5_ASAP7_75t_R c6121(
.A1(net6125),
.A2(net6177),
.B(net6176),
.C(net6178),
.Y(net6179)
);

OA222x2_ASAP7_75t_R c6122(
.A1(net6177),
.A2(net6145),
.B1(net6163),
.B2(net6153),
.C1(net6085),
.C2(net10258),
.Y(net6180)
);

OA21x2_ASAP7_75t_R c6123(
.A1(net6166),
.A2(net9823),
.B(net10256),
.Y(net6181)
);

OAI21x1_ASAP7_75t_R c6124(
.A1(net6055),
.A2(net6144),
.B(net6169),
.Y(net6182)
);

HB2xp67_ASAP7_75t_R c6125(
.A(net10061),
.Y(net6183)
);

NOR2xp33_ASAP7_75t_R c6126(
.A(net6169),
.B(net6160),
.Y(net6184)
);

OA211x2_ASAP7_75t_R c6127(
.A1(net5111),
.A2(net3400),
.B(net10153),
.C(net10258),
.Y(net6185)
);

OAI21xp33_ASAP7_75t_R c6128(
.A1(net6184),
.A2(net6169),
.B(net9722),
.Y(net6186)
);

OAI21xp5_ASAP7_75t_R c6129(
.A1(net6176),
.A2(net6178),
.B(net6166),
.Y(net6187)
);

OR3x1_ASAP7_75t_R c6130(
.A(net6184),
.B(net4166),
.C(net9918),
.Y(net6188)
);

NOR2xp67_ASAP7_75t_R c6131(
.A(net6163),
.B(net9967),
.Y(net6189)
);

OR3x2_ASAP7_75t_R c6132(
.A(net6066),
.B(net6166),
.C(net6189),
.Y(net6190)
);

AOI311xp33_ASAP7_75t_R c6133(
.A1(net5769),
.A2(net6147),
.A3(net6169),
.B(net6189),
.C(net6122),
.Y(net6191)
);

OR2x2_ASAP7_75t_R c6134(
.A(net6163),
.B(net6117),
.Y(net6192)
);

HB3xp67_ASAP7_75t_R c6135(
.A(net10566),
.Y(net6193)
);

HB4xp67_ASAP7_75t_R c6136(
.A(net10423),
.Y(net6194)
);

OR3x4_ASAP7_75t_R c6137(
.A(net6147),
.B(net6189),
.C(net6169),
.Y(net6195)
);

DFFASRHQNx1_ASAP7_75t_R c6138(
.D(net6194),
.RESETN(net6195),
.SETN(net4310),
.CLK(clk),
.QN(net6196)
);

AND3x1_ASAP7_75t_R c6139(
.A(net6049),
.B(net6172),
.C(net6154),
.Y(net6197)
);

AND3x2_ASAP7_75t_R c6140(
.A(net6148),
.B(net6196),
.C(net6189),
.Y(net6198)
);

SDFHx1_ASAP7_75t_R c6141(
.D(net6197),
.SE(net6192),
.SI(net6189),
.CLK(clk),
.QN(net6199)
);

INVx11_ASAP7_75t_R c6142(
.A(net10127),
.Y(net6200)
);

INVx13_ASAP7_75t_R c6143(
.A(net5275),
.Y(net6201)
);

INVx1_ASAP7_75t_R c6144(
.A(net10546),
.Y(net6202)
);

INVx2_ASAP7_75t_R c6145(
.A(net10169),
.Y(net6203)
);

INVx3_ASAP7_75t_R c6146(
.A(net10357),
.Y(net6204)
);

OR2x4_ASAP7_75t_R c6147(
.A(net5077),
.B(net6203),
.Y(net6205)
);

INVx4_ASAP7_75t_R c6148(
.A(net5355),
.Y(net6206)
);

OR2x6_ASAP7_75t_R c6149(
.A(net4373),
.B(net5284),
.Y(net6207)
);

INVx5_ASAP7_75t_R c6150(
.A(net9914),
.Y(net6208)
);

XNOR2x1_ASAP7_75t_R c6151(
.B(net5147),
.A(net9882),
.Y(net6209)
);

INVx6_ASAP7_75t_R c6152(
.A(net5225),
.Y(net6210)
);

XNOR2x2_ASAP7_75t_R c6153(
.A(net4957),
.B(net6203),
.Y(net6211)
);

ICGx2_ASAP7_75t_R c6154(
.ENA(net5346),
.SE(net5296),
.CLK(clk),
.GCLK(net6212)
);

INVx8_ASAP7_75t_R c6155(
.A(net9155),
.Y(net6213)
);

XNOR2xp5_ASAP7_75t_R c6156(
.A(net6131),
.B(net10258),
.Y(net6214)
);

XOR2x1_ASAP7_75t_R c6157(
.A(net6212),
.B(net9901),
.Y(net6215)
);

XOR2x2_ASAP7_75t_R c6158(
.A(net5286),
.B(net4373),
.Y(net6216)
);

XOR2xp5_ASAP7_75t_R c6159(
.A(net6199),
.B(net4257),
.Y(net6217)
);

INVxp33_ASAP7_75t_R c6160(
.A(net10386),
.Y(net6218)
);

AND2x2_ASAP7_75t_R c6161(
.A(net5274),
.B(net10267),
.Y(net6219)
);

AND2x4_ASAP7_75t_R c6162(
.A(net5305),
.B(net4214),
.Y(net6220)
);

AND2x6_ASAP7_75t_R c6163(
.A(net6188),
.B(net5167),
.Y(net6221)
);

INVxp67_ASAP7_75t_R c6164(
.A(net10420),
.Y(net6222)
);

BUFx10_ASAP7_75t_R c6165(
.A(net9155),
.Y(net6223)
);

HAxp5_ASAP7_75t_R c6166(
.A(net5147),
.B(net6204),
.CON(net6225),
.SN(net6224)
);

NAND2x1_ASAP7_75t_R c6167(
.A(net6205),
.B(net5343),
.Y(net6226)
);

NAND2x1p5_ASAP7_75t_R c6168(
.A(net5291),
.B(net6212),
.Y(net6227)
);

NAND2x2_ASAP7_75t_R c6169(
.A(net6217),
.B(net6209),
.Y(net6228)
);

NAND2xp33_ASAP7_75t_R c6170(
.A(net5833),
.B(net5311),
.Y(net6229)
);

BUFx12_ASAP7_75t_R c6171(
.A(net5167),
.Y(net6230)
);

NAND2xp5_ASAP7_75t_R c6172(
.A(net4402),
.B(net6207),
.Y(net6231)
);

BUFx12f_ASAP7_75t_R c6173(
.A(net10118),
.Y(net6232)
);

BUFx16f_ASAP7_75t_R c6174(
.A(net4214),
.Y(net6233)
);

NAND2xp67_ASAP7_75t_R c6175(
.A(net6123),
.B(net5312),
.Y(net6234)
);

AOI32xp33_ASAP7_75t_R c6176(
.A1(net6202),
.A2(net6203),
.A3(net6204),
.B1(net6080),
.B2(net10127),
.Y(net6235)
);

NOR2x1_ASAP7_75t_R c6177(
.A(net3483),
.B(net6233),
.Y(net6236)
);

NOR2x1p5_ASAP7_75t_R c6178(
.A(net6232),
.B(net5275),
.Y(net6237)
);

NOR2x2_ASAP7_75t_R c6179(
.A(net5322),
.B(net3878),
.Y(net6238)
);

NOR2xp33_ASAP7_75t_R c6180(
.A(net6238),
.B(net5225),
.Y(net6239)
);

AND3x4_ASAP7_75t_R c6181(
.A(net6231),
.B(net6220),
.C(net5325),
.Y(net6240)
);

BUFx24_ASAP7_75t_R c6182(
.A(net6207),
.Y(net6241)
);

NOR2xp67_ASAP7_75t_R c6183(
.A(net6236),
.B(net4369),
.Y(net6242)
);

OR2x2_ASAP7_75t_R c6184(
.A(net4422),
.B(net6240),
.Y(net6243)
);

BUFx2_ASAP7_75t_R c6185(
.A(net6124),
.Y(net6244)
);

OR2x4_ASAP7_75t_R c6186(
.A(net6223),
.B(net5077),
.Y(net6245)
);

OR2x6_ASAP7_75t_R c6187(
.A(net3490),
.B(net6232),
.Y(net6246)
);

AO21x1_ASAP7_75t_R c6188(
.A1(net6234),
.A2(net6199),
.B(net6212),
.Y(net6247)
);

AO21x2_ASAP7_75t_R c6189(
.A1(net6200),
.A2(net6222),
.B(net10133),
.Y(net6248)
);

XNOR2x1_ASAP7_75t_R c6190(
.B(net6219),
.A(net6238),
.Y(net6249)
);

XNOR2x2_ASAP7_75t_R c6191(
.A(net6233),
.B(net6248),
.Y(net6250)
);

XNOR2xp5_ASAP7_75t_R c6192(
.A(net6241),
.B(net6248),
.Y(net6251)
);

XOR2x1_ASAP7_75t_R c6193(
.A(net6121),
.B(net5275),
.Y(net6252)
);

XOR2x2_ASAP7_75t_R c6194(
.A(net6167),
.B(net6224),
.Y(net6253)
);

BUFx3_ASAP7_75t_R c6195(
.A(net6218),
.Y(net6254)
);

BUFx4_ASAP7_75t_R c6196(
.A(net10432),
.Y(net6255)
);

XOR2xp5_ASAP7_75t_R c6197(
.A(net6245),
.B(net6227),
.Y(net6256)
);

AND2x2_ASAP7_75t_R c6198(
.A(net6228),
.B(net6196),
.Y(net6257)
);

BUFx4f_ASAP7_75t_R c6199(
.A(net10129),
.Y(net6258)
);

AOI21x1_ASAP7_75t_R c6200(
.A1(net6257),
.A2(net6258),
.B(net6146),
.Y(net6259)
);

AND2x4_ASAP7_75t_R c6201(
.A(net6237),
.B(net6258),
.Y(net6260)
);

AOI21xp33_ASAP7_75t_R c6202(
.A1(net6208),
.A2(net6245),
.B(net5346),
.Y(net6261)
);

BUFx5_ASAP7_75t_R c6203(
.A(net10122),
.Y(net6262)
);

AND2x6_ASAP7_75t_R c6204(
.A(net6244),
.B(net6200),
.Y(net6263)
);

HAxp5_ASAP7_75t_R c6205(
.A(net6250),
.B(net6058),
.CON(net6264)
);

AOI21xp5_ASAP7_75t_R c6206(
.A1(net6215),
.A2(net6256),
.B(net6234),
.Y(net6265)
);

NAND2x1_ASAP7_75t_R c6207(
.A(net6212),
.B(net6167),
.Y(net6266)
);

NAND2x1p5_ASAP7_75t_R c6208(
.A(net6253),
.B(net6207),
.Y(net6267)
);

NAND2x2_ASAP7_75t_R c6209(
.A(net6260),
.B(net6241),
.Y(net6268)
);

FAx1_ASAP7_75t_R c6210(
.A(net6254),
.B(net6256),
.CI(net6258),
.SN(net6270),
.CON(net6269)
);

NAND2xp33_ASAP7_75t_R c6211(
.A(net6262),
.B(net6253),
.Y(net6271)
);

MAJIxp5_ASAP7_75t_R c6212(
.A(net6269),
.B(net6258),
.C(net9815),
.Y(net6272)
);

MAJx2_ASAP7_75t_R c6213(
.A(net6196),
.B(net6263),
.C(net5726),
.Y(net6273)
);

OA33x2_ASAP7_75t_R c6214(
.A1(net6240),
.A2(net6270),
.A3(net6225),
.B1(net5833),
.B2(net2474),
.B3(net5325),
.Y(net6274)
);

MAJx3_ASAP7_75t_R c6215(
.A(net6270),
.B(net6272),
.C(net6256),
.Y(net6275)
);

NAND3x1_ASAP7_75t_R c6216(
.A(net6159),
.B(net6121),
.C(net6248),
.Y(net6276)
);

NAND3x2_ASAP7_75t_R c6217(
.B(net6033),
.C(net6245),
.A(net6221),
.Y(net6277)
);

NAND3xp33_ASAP7_75t_R c6218(
.A(net6266),
.B(net1652),
.C(net10172),
.Y(net6278)
);

NOR3x1_ASAP7_75t_R c6219(
.A(net6251),
.B(net6268),
.C(net6273),
.Y(net6279)
);

OAI222xp33_ASAP7_75t_R c6220(
.A1(net6275),
.A2(net6253),
.B1(net6272),
.B2(net6191),
.C1(net6263),
.C2(net6204),
.Y(net6280)
);

OAI321xp33_ASAP7_75t_R c6221(
.A1(net6277),
.A2(net6220),
.A3(net6146),
.B1(net6201),
.B2(net10172),
.C(net10273),
.Y(net6281)
);

NOR3x2_ASAP7_75t_R c6222(
.B(net6271),
.C(net6233),
.A(net10273),
.Y(net6282)
);

NOR3xp33_ASAP7_75t_R c6223(
.A(net6278),
.B(net6281),
.C(net10273),
.Y(net6283)
);

OA21x2_ASAP7_75t_R c6224(
.A1(net6258),
.A2(net6282),
.B(net10273),
.Y(net6284)
);

OAI21x1_ASAP7_75t_R c6225(
.A1(net5426),
.A2(net3564),
.B(net5412),
.Y(net6285)
);

NAND2xp5_ASAP7_75t_R c6226(
.A(net2578),
.B(net6285),
.Y(net6286)
);

NAND2xp67_ASAP7_75t_R c6227(
.A(net5352),
.B(net5135),
.Y(net6287)
);

BUFx6f_ASAP7_75t_R c6228(
.A(net10573),
.Y(net6288)
);

BUFx8_ASAP7_75t_R c6229(
.A(net5407),
.Y(net6289)
);

NOR2x1_ASAP7_75t_R c6230(
.A(net4431),
.B(net5274),
.Y(net6290)
);

CKINVDCx10_ASAP7_75t_R c6231(
.A(net9167),
.Y(net6291)
);

NOR2x1p5_ASAP7_75t_R c6232(
.A(net5274),
.B(out1),
.Y(net6292)
);

CKINVDCx11_ASAP7_75t_R c6233(
.A(net10042),
.Y(net6293)
);

CKINVDCx12_ASAP7_75t_R c6234(
.A(net10352),
.Y(net6294)
);

CKINVDCx14_ASAP7_75t_R c6235(
.A(net5726),
.Y(net6295)
);

NOR2x2_ASAP7_75t_R c6236(
.A(net6290),
.B(net6204),
.Y(net6296)
);

NOR2xp33_ASAP7_75t_R c6237(
.A(net5097),
.B(net6201),
.Y(net6297)
);

NOR2xp67_ASAP7_75t_R c6238(
.A(net6220),
.B(net5369),
.Y(net6298)
);

OR2x2_ASAP7_75t_R c6239(
.A(net6291),
.B(net6289),
.Y(net6299)
);

OR2x4_ASAP7_75t_R c6240(
.A(net4357),
.B(net10133),
.Y(net6300)
);

CKINVDCx16_ASAP7_75t_R c6241(
.A(net10371),
.Y(net6301)
);

CKINVDCx20_ASAP7_75t_R c6242(
.A(net3522),
.Y(net6302)
);

OR2x6_ASAP7_75t_R c6243(
.A(net3587),
.B(net4502),
.Y(net6303)
);

SDFHx2_ASAP7_75t_R c6244(
.D(net5315),
.SE(net5407),
.SI(net6122),
.CLK(clk),
.QN(net6304)
);

CKINVDCx5p33_ASAP7_75t_R c6245(
.A(net9167),
.Y(net6305)
);

CKINVDCx6p67_ASAP7_75t_R c6246(
.A(net6230),
.Y(net6306)
);

XNOR2x1_ASAP7_75t_R c6247(
.B(net6210),
.A(net6289),
.Y(net6307)
);

XNOR2x2_ASAP7_75t_R c6248(
.A(net6301),
.B(net4483),
.Y(net6308)
);

CKINVDCx8_ASAP7_75t_R c6249(
.A(net10455),
.Y(net6309)
);

XNOR2xp5_ASAP7_75t_R c6250(
.A(net5437),
.B(net6300),
.Y(net6310)
);

XOR2x1_ASAP7_75t_R c6251(
.A(net6291),
.B(out0),
.Y(net6311)
);

XOR2x2_ASAP7_75t_R c6252(
.A(net6278),
.B(net6201),
.Y(net6312)
);

CKINVDCx9p33_ASAP7_75t_R c6253(
.A(net10397),
.Y(net6313)
);

XOR2xp5_ASAP7_75t_R c6254(
.A(net5363),
.B(net6301),
.Y(net6314)
);

OAI21xp33_ASAP7_75t_R c6255(
.A1(net6312),
.A2(net6314),
.B(net6304),
.Y(net6315)
);

AND2x2_ASAP7_75t_R c6256(
.A(net6304),
.B(net10153),
.Y(net6316)
);

OAI21xp5_ASAP7_75t_R c6257(
.A1(net6315),
.A2(net6307),
.B(net5315),
.Y(net6317)
);

HB1xp67_ASAP7_75t_R c6258(
.A(net6248),
.Y(net6318)
);

AND2x4_ASAP7_75t_R c6259(
.A(net6308),
.B(net6213),
.Y(net6319)
);

NAND5xp2_ASAP7_75t_R c6260(
.A(net6019),
.B(net5377),
.C(net6296),
.D(net6301),
.E(net5411),
.Y(net6320)
);

AND2x6_ASAP7_75t_R c6261(
.A(net5387),
.B(net4467),
.Y(net6321)
);

HAxp5_ASAP7_75t_R c6262(
.A(net5312),
.B(net5407),
.CON(net6322)
);

HB2xp67_ASAP7_75t_R c6263(
.A(net6156),
.Y(net6323)
);

NAND2x1_ASAP7_75t_R c6264(
.A(net6306),
.B(net5414),
.Y(net6324)
);

HB3xp67_ASAP7_75t_R c6265(
.A(net6296),
.Y(net6325)
);

SDFHx3_ASAP7_75t_R c6266(
.D(net6319),
.SE(net6296),
.SI(net6201),
.CLK(clk),
.QN(net6326)
);

OR3x1_ASAP7_75t_R c6267(
.A(net5392),
.B(net3587),
.C(net5414),
.Y(net6327)
);

NAND2x1p5_ASAP7_75t_R c6268(
.A(net6255),
.B(net6292),
.Y(net6328)
);

NAND2x2_ASAP7_75t_R c6269(
.A(net6314),
.B(net6328),
.Y(net6329)
);

HB4xp67_ASAP7_75t_R c6270(
.A(net10350),
.Y(net6330)
);

INVx11_ASAP7_75t_R c6271(
.A(net6227),
.Y(net6331)
);

SDFHx4_ASAP7_75t_R c6272(
.D(net5401),
.SE(net6325),
.SI(net6331),
.CLK(clk),
.QN(net6332)
);

INVx13_ASAP7_75t_R c6273(
.A(net10155),
.Y(net6333)
);

NAND2xp33_ASAP7_75t_R c6274(
.A(net6321),
.B(net6301),
.Y(net6334)
);

INVx1_ASAP7_75t_R c6275(
.A(net10420),
.Y(net6335)
);

NAND2xp5_ASAP7_75t_R c6276(
.A(net6298),
.B(net6296),
.Y(net6336)
);

NOR5xp2_ASAP7_75t_R c6277(
.A(net4360),
.B(net6173),
.C(net5411),
.D(net4353),
.E(net6204),
.Y(net6337)
);

NAND2xp67_ASAP7_75t_R c6278(
.A(net6318),
.B(net6334),
.Y(net6338)
);

OR3x2_ASAP7_75t_R c6279(
.A(net4467),
.B(net6338),
.C(net5392),
.Y(net6339)
);

NOR2x1_ASAP7_75t_R c6280(
.A(net6322),
.B(net6221),
.Y(net6340)
);

NOR2x1p5_ASAP7_75t_R c6281(
.A(net2661),
.B(net9708),
.Y(net6341)
);

OR3x4_ASAP7_75t_R c6282(
.A(net6281),
.B(net6340),
.C(net5409),
.Y(net6342)
);

INVx2_ASAP7_75t_R c6283(
.A(net10467),
.Y(net6343)
);

NOR2x2_ASAP7_75t_R c6284(
.A(net4483),
.B(net6298),
.Y(net6344)
);

AND3x1_ASAP7_75t_R c6285(
.A(net6344),
.B(net6306),
.C(net6281),
.Y(net6345)
);

NOR2xp33_ASAP7_75t_R c6286(
.A(net9697),
.B(net10098),
.Y(net6346)
);

NOR2xp67_ASAP7_75t_R c6287(
.A(net6326),
.B(net9823),
.Y(net6347)
);

OA221x2_ASAP7_75t_R c6288(
.A1(net5400),
.A2(net6154),
.B1(net3587),
.B2(net6289),
.C(net6224),
.Y(net6348)
);

OR2x2_ASAP7_75t_R c6289(
.A(net5432),
.B(net9949),
.Y(net6349)
);

AND3x2_ASAP7_75t_R c6290(
.A(net6326),
.B(net6338),
.C(net6296),
.Y(net6350)
);

INVx3_ASAP7_75t_R c6291(
.A(net10362),
.Y(net6351)
);

AND3x4_ASAP7_75t_R c6292(
.A(net6294),
.B(net6332),
.C(net10098),
.Y(net6352)
);

INVx4_ASAP7_75t_R c6293(
.A(net10523),
.Y(net6353)
);

OR2x4_ASAP7_75t_R c6294(
.A(net6333),
.B(net6343),
.Y(net6354)
);

AO21x1_ASAP7_75t_R c6295(
.A1(net6284),
.A2(net6352),
.B(net6335),
.Y(net6355)
);

AO21x2_ASAP7_75t_R c6296(
.A1(net6352),
.A2(net5422),
.B(net10274),
.Y(net6356)
);

OAI221xp5_ASAP7_75t_R c6297(
.A1(net6309),
.A2(net6347),
.B1(net5443),
.B2(net5398),
.C(net10260),
.Y(net6357)
);

AOI21x1_ASAP7_75t_R c6298(
.A1(net4501),
.A2(net6321),
.B(net9987),
.Y(net6358)
);

SDFLx1_ASAP7_75t_R c6299(
.D(net6358),
.SE(net6350),
.SI(net6356),
.CLK(clk),
.QN(net6359)
);

OA22x2_ASAP7_75t_R c6300(
.A1(net6330),
.A2(net5392),
.B1(net5411),
.B2(net6319),
.Y(net6360)
);

SDFLx2_ASAP7_75t_R c6301(
.D(net6336),
.SE(net6359),
.SI(net6347),
.CLK(clk),
.QN(net6361)
);

AOI21xp33_ASAP7_75t_R c6302(
.A1(net6359),
.A2(net6343),
.B(net10151),
.Y(net6362)
);

AOI21xp5_ASAP7_75t_R c6303(
.A1(net6242),
.A2(net6346),
.B(net6362),
.Y(net6363)
);

FAx1_ASAP7_75t_R c6304(
.A(net6357),
.B(net6356),
.CI(net6361),
.SN(net6364)
);

MAJIxp5_ASAP7_75t_R c6305(
.A(net5369),
.B(net6364),
.C(net6359),
.Y(net6365)
);

INVx5_ASAP7_75t_R c6306(
.A(net10485),
.Y(net6366)
);

MAJx2_ASAP7_75t_R c6307(
.A(net6299),
.B(net6353),
.C(net4469),
.Y(net6367)
);

OR2x6_ASAP7_75t_R c6308(
.A(net5526),
.B(net6292),
.Y(net6368)
);

OA31x2_ASAP7_75t_R c6309(
.A1(net2719),
.A2(net5526),
.A3(net10230),
.B1(net10260),
.Y(net6369)
);

XNOR2x1_ASAP7_75t_R c6310(
.B(net5413),
.A(net9707),
.Y(net6370)
);

XNOR2x2_ASAP7_75t_R c6311(
.A(net5452),
.B(net4535),
.Y(net6371)
);

MAJx3_ASAP7_75t_R c6312(
.A(net4566),
.B(net6354),
.C(net5485),
.Y(net6372)
);

XNOR2xp5_ASAP7_75t_R c6313(
.A(net5516),
.B(net5526),
.Y(net6373)
);

NAND3x1_ASAP7_75t_R c6314(
.A(net4543),
.B(net5520),
.C(net10230),
.Y(net6374)
);

XOR2x1_ASAP7_75t_R c6315(
.A(net3639),
.B(net5516),
.Y(net6375)
);

XOR2x2_ASAP7_75t_R c6316(
.A(net5483),
.B(net5479),
.Y(net6376)
);

INVx6_ASAP7_75t_R c6317(
.A(net10348),
.Y(out3)
);

XOR2xp5_ASAP7_75t_R c6318(
.A(net5444),
.B(net10261),
.Y(net6377)
);

SDFLx3_ASAP7_75t_R c6319(
.D(net6216),
.SE(net6373),
.SI(net5461),
.CLK(clk),
.QN(net6378)
);

AND2x2_ASAP7_75t_R c6320(
.A(net6285),
.B(net6378),
.Y(net6379)
);

SDFLx4_ASAP7_75t_R c6321(
.D(net6372),
.SE(net6376),
.SI(net6328),
.CLK(clk),
.QN(net6380)
);

NAND3x2_ASAP7_75t_R c6322(
.B(net6292),
.C(net5325),
.A(net3662),
.Y(net6381)
);

AND2x4_ASAP7_75t_R c6323(
.A(net5496),
.B(net4543),
.Y(net6382)
);

INVx8_ASAP7_75t_R c6324(
.A(net10348),
.Y(net6383)
);

NAND3xp33_ASAP7_75t_R c6325(
.A(net6328),
.B(net5413),
.C(net5444),
.Y(net6384)
);

AND2x6_ASAP7_75t_R c6326(
.A(net5512),
.B(net6378),
.Y(net6385)
);

DFFASRHQNx1_ASAP7_75t_R c6327(
.D(net6374),
.RESETN(net6304),
.SETN(net6383),
.CLK(clk),
.QN(net6386)
);

NOR3x1_ASAP7_75t_R c6328(
.A(net5479),
.B(net6292),
.C(net4523),
.Y(net6387)
);

HAxp5_ASAP7_75t_R c6329(
.A(net5460),
.B(net9971),
.CON(net6389),
.SN(net6388)
);

SDFHx1_ASAP7_75t_R c6330(
.D(net3662),
.SE(net4589),
.SI(net5866),
.CLK(clk),
.QN(net6390)
);

NOR3x2_ASAP7_75t_R c6331(
.B(net5449),
.C(net1774),
.A(net5415),
.Y(net6391)
);

OAI211xp5_ASAP7_75t_R c6332(
.A1(net6375),
.A2(net6391),
.B(net5260),
.C(net10274),
.Y(net6392)
);

NOR3xp33_ASAP7_75t_R c6333(
.A(net5472),
.B(net6386),
.C(net6365),
.Y(net6393)
);

OA21x2_ASAP7_75t_R c6334(
.A1(net5300),
.A2(net3676),
.B(net6201),
.Y(net6394)
);

OAI21x1_ASAP7_75t_R c6335(
.A1(net6389),
.A2(net5525),
.B(net2703),
.Y(net6395)
);

NAND2x1_ASAP7_75t_R c6336(
.A(net4576),
.B(net4594),
.Y(net6396)
);

OAI21xp33_ASAP7_75t_R c6337(
.A1(net6390),
.A2(net6368),
.B(net4535),
.Y(net6397)
);

OAI21xp5_ASAP7_75t_R c6338(
.A1(net6331),
.A2(net4543),
.B(net5483),
.Y(net6398)
);

NAND2x1p5_ASAP7_75t_R c6339(
.A(net6122),
.B(net6390),
.Y(net6399)
);

OAI22x1_ASAP7_75t_R c6340(
.A1(net5415),
.A2(net6390),
.B1(net4523),
.B2(net6354),
.Y(net6400)
);

OR3x1_ASAP7_75t_R c6341(
.A(net6369),
.B(net6343),
.C(net5456),
.Y(net6401)
);

OR3x2_ASAP7_75t_R c6342(
.A(net5460),
.B(net5507),
.C(net5456),
.Y(net6402)
);

OAI22xp33_ASAP7_75t_R c6343(
.A1(net6386),
.A2(net4603),
.B1(net6396),
.B2(net5492),
.Y(net6403)
);

OR3x4_ASAP7_75t_R c6344(
.A(net6400),
.B(net6396),
.C(net9794),
.Y(net6404)
);

INVxp33_ASAP7_75t_R c6345(
.A(net10155),
.Y(net6405)
);

AND3x1_ASAP7_75t_R c6346(
.A(net4535),
.B(net6328),
.C(net5461),
.Y(net6406)
);

AND3x2_ASAP7_75t_R c6347(
.A(net6394),
.B(net6387),
.C(net5357),
.Y(net6407)
);

AND3x4_ASAP7_75t_R c6348(
.A(net5494),
.B(net6396),
.C(net3662),
.Y(net6408)
);

AO21x1_ASAP7_75t_R c6349(
.A1(net5463),
.A2(net6388),
.B(out5),
.Y(net6409)
);

INVxp67_ASAP7_75t_R c6350(
.A(net10394),
.Y(net6410)
);

AO21x2_ASAP7_75t_R c6351(
.A1(net5518),
.A2(net6354),
.B(net6381),
.Y(net6411)
);

AOI21x1_ASAP7_75t_R c6352(
.A1(net5507),
.A2(net6404),
.B(net5357),
.Y(net6412)
);

AOI21xp33_ASAP7_75t_R c6353(
.A1(net6324),
.A2(net6396),
.B(net4593),
.Y(net6413)
);

NAND2x2_ASAP7_75t_R c6354(
.A(net3628),
.B(net6396),
.Y(net6414)
);

AOI21xp5_ASAP7_75t_R c6355(
.A1(net6408),
.A2(net6376),
.B(net6409),
.Y(net6415)
);

NAND2xp33_ASAP7_75t_R c6356(
.A(net6239),
.B(net5520),
.Y(net6416)
);

FAx1_ASAP7_75t_R c6357(
.A(net6408),
.B(net6416),
.CI(net9897),
.SN(net6417)
);

NAND2xp5_ASAP7_75t_R c6358(
.A(net6287),
.B(net6386),
.Y(net6418)
);

MAJIxp5_ASAP7_75t_R c6359(
.A(net5464),
.B(net6324),
.C(net9852),
.Y(net6419)
);

OAI311xp33_ASAP7_75t_R c6360(
.A1(net6418),
.A2(net5415),
.A3(net6263),
.B1(net6409),
.C1(net9736),
.Y(net6420)
);

MAJx2_ASAP7_75t_R c6361(
.A(net5485),
.B(net6400),
.C(net5290),
.Y(net6421)
);

MAJx3_ASAP7_75t_R c6362(
.A(net6414),
.B(net6402),
.C(net4468),
.Y(net6422)
);

NAND3x1_ASAP7_75t_R c6363(
.A(net6377),
.B(net5520),
.C(net6390),
.Y(net6423)
);

NAND3x2_ASAP7_75t_R c6364(
.B(net6373),
.C(net6403),
.A(net4593),
.Y(net6424)
);

NAND3xp33_ASAP7_75t_R c6365(
.A(net6420),
.B(net5496),
.C(net6324),
.Y(net6425)
);

NOR3x1_ASAP7_75t_R c6366(
.A(net6421),
.B(net6400),
.C(net6380),
.Y(net6426)
);

NOR3x2_ASAP7_75t_R c6367(
.B(net6423),
.C(net6370),
.A(net5300),
.Y(net6427)
);

NOR3xp33_ASAP7_75t_R c6368(
.A(net5514),
.B(net6426),
.C(net6379),
.Y(net6428)
);

OA21x2_ASAP7_75t_R c6369(
.A1(net6354),
.A2(net6426),
.B(net6409),
.Y(net6429)
);

OAI22xp5_ASAP7_75t_R c6370(
.A1(net2703),
.A2(net5512),
.B1(net6390),
.B2(net6408),
.Y(net6430)
);

OAI21x1_ASAP7_75t_R c6371(
.A1(net6410),
.A2(net6428),
.B(net6416),
.Y(net6431)
);

SDFHx2_ASAP7_75t_R c6372(
.D(net6428),
.SE(net5415),
.SI(net6365),
.CLK(clk),
.QN(net6432)
);

OAI21xp33_ASAP7_75t_R c6373(
.A1(net4593),
.A2(net6389),
.B(net9893),
.Y(net6433)
);

SDFHx3_ASAP7_75t_R c6374(
.D(net6379),
.SE(net6411),
.SI(net10275),
.CLK(clk),
.QN(net6434)
);

OAI21xp5_ASAP7_75t_R c6375(
.A1(net6348),
.A2(net6408),
.B(net4523),
.Y(net6435)
);

OR3x1_ASAP7_75t_R c6376(
.A(net6201),
.B(net6419),
.C(net6426),
.Y(net6436)
);

OR3x2_ASAP7_75t_R c6377(
.A(net6433),
.B(net6416),
.C(net6422),
.Y(net6437)
);

OR3x4_ASAP7_75t_R c6378(
.A(net6398),
.B(net5267),
.C(net6416),
.Y(net6438)
);

AND3x1_ASAP7_75t_R c6379(
.A(net6422),
.B(net6396),
.C(net6432),
.Y(net6439)
);

AND3x2_ASAP7_75t_R c6380(
.A(net6439),
.B(net5452),
.C(net9893),
.Y(net6440)
);

SDFHx4_ASAP7_75t_R c6381(
.D(net6376),
.SE(net6437),
.SI(net6421),
.CLK(clk),
.QN(net6441)
);

AND3x4_ASAP7_75t_R c6382(
.A(net5467),
.B(net6331),
.C(net10274),
.Y(net6442)
);

AO21x1_ASAP7_75t_R c6383(
.A1(net6432),
.A2(net6436),
.B(net9960),
.Y(net6443)
);

SDFLx1_ASAP7_75t_R c6384(
.D(net6441),
.SE(net6443),
.SI(net9736),
.CLK(clk),
.QN(net6444)
);

OAI31xp33_ASAP7_75t_R c6385(
.A1(net6436),
.A2(net6424),
.A3(net6441),
.B(net4589),
.Y(net6445)
);

OAI31xp67_ASAP7_75t_R c6386(
.A1(net6442),
.A2(net6410),
.A3(net6381),
.B(net10275),
.Y(net6446)
);

OAI32xp33_ASAP7_75t_R c6387(
.A1(net6385),
.A2(net6446),
.A3(net6347),
.B1(net9943),
.B2(net10275),
.Y(net6447)
);

OR4x1_ASAP7_75t_R c6388(
.A(net6365),
.B(net6439),
.C(net6408),
.D(net9779),
.Y(net6448)
);

OR4x2_ASAP7_75t_R c6389(
.A(net6443),
.B(net6405),
.C(net3635),
.D(net6446),
.Y(net6449)
);

OR5x1_ASAP7_75t_R c6390(
.A(net4523),
.B(net6418),
.C(net6388),
.D(net1653),
.E(net9831),
.Y(net6450)
);

BUFx10_ASAP7_75t_R c6391(
.A(net3728),
.Y(net6451)
);

BUFx12_ASAP7_75t_R c6392(
.A(net9147),
.Y(net6452)
);

BUFx12f_ASAP7_75t_R c6393(
.A(net4681),
.Y(net6453)
);

NAND2xp67_ASAP7_75t_R c6394(
.A(net5560),
.B(net4657),
.Y(net6454)
);

BUFx16f_ASAP7_75t_R c6395(
.A(net3759),
.Y(net6455)
);

BUFx24_ASAP7_75t_R c6396(
.A(net4657),
.Y(net6456)
);

BUFx2_ASAP7_75t_R c6397(
.A(net3710),
.Y(net6457)
);

ICGx2p67DC_ASAP7_75t_R c6398(
.ENA(net6451),
.SE(net5531),
.CLK(clk),
.GCLK(net6458)
);

NOR2x1_ASAP7_75t_R c6399(
.A(net4642),
.B(net5532),
.Y(net6459)
);

BUFx3_ASAP7_75t_R c6400(
.A(net968),
.Y(net6460)
);

BUFx4_ASAP7_75t_R c6401(
.A(net4616),
.Y(net6461)
);

BUFx4f_ASAP7_75t_R c6402(
.A(net1861),
.Y(net6462)
);

BUFx5_ASAP7_75t_R c6403(
.A(net5549),
.Y(net6463)
);

BUFx6f_ASAP7_75t_R c6404(
.A(net6461),
.Y(net6464)
);

BUFx8_ASAP7_75t_R c6405(
.A(net4642),
.Y(net6465)
);

CKINVDCx10_ASAP7_75t_R c6406(
.A(net5533),
.Y(net6466)
);

CKINVDCx11_ASAP7_75t_R c6407(
.A(net3747),
.Y(net6467)
);

CKINVDCx12_ASAP7_75t_R c6408(
.A(net6457),
.Y(net6468)
);

CKINVDCx14_ASAP7_75t_R c6409(
.A(net5539),
.Y(net6469)
);

CKINVDCx16_ASAP7_75t_R c6410(
.A(net4610),
.Y(net6470)
);

NOR2x1p5_ASAP7_75t_R c6411(
.A(net3707),
.B(net10264),
.Y(net6471)
);

CKINVDCx20_ASAP7_75t_R c6412(
.A(net6462),
.Y(net6472)
);

CKINVDCx5p33_ASAP7_75t_R c6413(
.A(net2811),
.Y(net6473)
);

NOR2x2_ASAP7_75t_R c6414(
.A(net5561),
.B(net5549),
.Y(net6474)
);

CKINVDCx6p67_ASAP7_75t_R c6415(
.A(net6469),
.Y(net6475)
);

CKINVDCx8_ASAP7_75t_R c6416(
.A(net9147),
.Y(net6476)
);

CKINVDCx9p33_ASAP7_75t_R c6417(
.A(net9211),
.Y(net6477)
);

NOR2xp33_ASAP7_75t_R c6418(
.A(net6476),
.B(net6460),
.Y(net6478)
);

HB1xp67_ASAP7_75t_R c6419(
.A(net9226),
.Y(net6479)
);

HB2xp67_ASAP7_75t_R c6420(
.A(net6478),
.Y(net6480)
);

NOR2xp67_ASAP7_75t_R c6421(
.A(net6465),
.B(net5609),
.Y(net6481)
);

OR2x2_ASAP7_75t_R c6422(
.A(net3759),
.B(net5597),
.Y(net6482)
);

OR2x4_ASAP7_75t_R c6423(
.A(net5581),
.B(net3728),
.Y(net6483)
);

OR2x6_ASAP7_75t_R c6424(
.A(net6455),
.B(net6458),
.Y(net6484)
);

XNOR2x1_ASAP7_75t_R c6425(
.B(net6471),
.A(net4616),
.Y(net6485)
);

HB3xp67_ASAP7_75t_R c6426(
.A(net6484),
.Y(net6486)
);

HB4xp67_ASAP7_75t_R c6427(
.A(net6460),
.Y(net6487)
);

XNOR2x2_ASAP7_75t_R c6428(
.A(net6487),
.B(net6484),
.Y(net6488)
);

XNOR2xp5_ASAP7_75t_R c6429(
.A(net6488),
.B(net3759),
.Y(net6489)
);

XOR2x1_ASAP7_75t_R c6430(
.A(net6485),
.B(net6486),
.Y(net6490)
);

INVx11_ASAP7_75t_R c6431(
.A(net9226),
.Y(net6491)
);

XOR2x2_ASAP7_75t_R c6432(
.A(net4618),
.B(net6488),
.Y(net6492)
);

ICGx3_ASAP7_75t_R c6433(
.ENA(net5600),
.SE(net10263),
.CLK(clk),
.GCLK(net6493)
);

INVx13_ASAP7_75t_R c6434(
.A(net4660),
.Y(net6494)
);

INVx1_ASAP7_75t_R c6435(
.A(net9282),
.Y(net6495)
);

INVx2_ASAP7_75t_R c6436(
.A(net9207),
.Y(net6496)
);

SDFLx2_ASAP7_75t_R c6437(
.D(net4610),
.SE(net6468),
.SI(net6451),
.CLK(clk),
.QN(net6497)
);

INVx3_ASAP7_75t_R c6438(
.A(net9660),
.Y(net6498)
);

INVx4_ASAP7_75t_R c6439(
.A(net6496),
.Y(net6499)
);

ICGx4DC_ASAP7_75t_R c6440(
.ENA(net6492),
.SE(net10219),
.CLK(clk),
.GCLK(net6500)
);

ICGx4_ASAP7_75t_R c6441(
.ENA(net6481),
.SE(net5593),
.CLK(clk),
.GCLK(net6501)
);

INVx5_ASAP7_75t_R c6442(
.A(net6498),
.Y(net6502)
);

XOR2xp5_ASAP7_75t_R c6443(
.A(net6459),
.B(net6500),
.Y(net6503)
);

AO21x2_ASAP7_75t_R c6444(
.A1(net6462),
.A2(net6496),
.B(net6499),
.Y(net6504)
);

AND2x2_ASAP7_75t_R c6445(
.A(net6468),
.B(net6503),
.Y(net6505)
);

AND2x4_ASAP7_75t_R c6446(
.A(net6476),
.B(net6504),
.Y(net6506)
);

AND2x6_ASAP7_75t_R c6447(
.A(net6472),
.B(net6504),
.Y(net6507)
);

A2O1A1Ixp33_ASAP7_75t_R c6448(
.A1(net6500),
.A2(net6499),
.B(net6470),
.C(net5609),
.Y(net6508)
);

AOI21x1_ASAP7_75t_R c6449(
.A1(net5581),
.A2(net6504),
.B(net5532),
.Y(net6509)
);

ICGx5_ASAP7_75t_R c6450(
.ENA(net4656),
.SE(net6508),
.CLK(clk),
.GCLK(net6510)
);

ICGx5p33DC_ASAP7_75t_R c6451(
.ENA(net6494),
.SE(net6505),
.CLK(clk),
.GCLK(net6511)
);

HAxp5_ASAP7_75t_R c6452(
.A(net6497),
.B(net10263),
.CON(net6513),
.SN(net6512)
);

NAND2x1_ASAP7_75t_R c6453(
.A(net6479),
.B(net6512),
.Y(net6514)
);

SDFLx3_ASAP7_75t_R c6454(
.D(net6456),
.SE(net6505),
.SI(net6488),
.CLK(clk),
.QN(net6515)
);

NAND2x1p5_ASAP7_75t_R c6455(
.A(net6502),
.B(net6515),
.Y(net6516)
);

NAND2x2_ASAP7_75t_R c6456(
.A(net6470),
.B(net6502),
.Y(net6517)
);

NAND2xp33_ASAP7_75t_R c6457(
.A(net5560),
.B(net6492),
.Y(net6518)
);

NAND2xp5_ASAP7_75t_R c6458(
.A(net5597),
.B(net6516),
.Y(net6519)
);

AOI21xp33_ASAP7_75t_R c6459(
.A1(net6515),
.A2(net4621),
.B(net9660),
.Y(net6520)
);

NAND2xp67_ASAP7_75t_R c6460(
.A(net6515),
.B(net6500),
.Y(net6521)
);

NOR2x1_ASAP7_75t_R c6461(
.A(net6499),
.B(net5605),
.Y(net6522)
);

SDFLx4_ASAP7_75t_R c6462(
.D(net6517),
.SE(net6474),
.SI(net6510),
.CLK(clk),
.QN(net6523)
);

OAI33xp33_ASAP7_75t_R c6463(
.A1(net6509),
.A2(net6475),
.A3(net6523),
.B1(net6451),
.B2(net6508),
.B3(net5609),
.Y(net6524)
);

AOI21xp5_ASAP7_75t_R c6464(
.A1(net6467),
.A2(net6470),
.B(net6514),
.Y(net6525)
);

FAx1_ASAP7_75t_R c6465(
.A(net6516),
.B(net5551),
.CI(net6519),
.SN(net6526)
);

MAJIxp5_ASAP7_75t_R c6466(
.A(net6495),
.B(net6523),
.C(net5532),
.Y(net6527)
);

MAJx2_ASAP7_75t_R c6467(
.A(net6507),
.B(net6478),
.C(net6501),
.Y(net6528)
);

MAJx3_ASAP7_75t_R c6468(
.A(net6528),
.B(net6525),
.C(net10276),
.Y(net6529)
);

AO222x2_ASAP7_75t_R c6469(
.A1(net6503),
.A2(net6529),
.B1(net6508),
.B2(net6510),
.C1(net5609),
.C2(net6455),
.Y(net6530)
);

DFFASRHQNx1_ASAP7_75t_R c6470(
.D(net6463),
.RESETN(net6527),
.SETN(net10277),
.CLK(clk),
.QN(net6531)
);

AND4x1_ASAP7_75t_R c6471(
.A(net6527),
.B(net6514),
.C(net6525),
.D(net10276),
.Y(net6532)
);

NAND3x1_ASAP7_75t_R c6472(
.A(net6529),
.B(net6525),
.C(net10277),
.Y(net6533)
);

AND4x2_ASAP7_75t_R c6473(
.A(net6531),
.B(net6520),
.C(net10276),
.D(net10277),
.Y(net6534)
);

INVx6_ASAP7_75t_R c6474(
.A(net6525),
.Y(net6535)
);

INVx8_ASAP7_75t_R c6475(
.A(net9114),
.Y(net6536)
);

INVxp33_ASAP7_75t_R c6476(
.A(net4756),
.Y(net6537)
);

INVxp67_ASAP7_75t_R c6477(
.A(net5668),
.Y(net6538)
);

NAND3x2_ASAP7_75t_R c6478(
.B(net5614),
.C(net4749),
.A(net3747),
.Y(net6539)
);

BUFx10_ASAP7_75t_R c6479(
.A(net4661),
.Y(net6540)
);

BUFx12_ASAP7_75t_R c6480(
.A(net5691),
.Y(net6541)
);

BUFx12f_ASAP7_75t_R c6481(
.A(net4697),
.Y(net6542)
);

BUFx16f_ASAP7_75t_R c6482(
.A(net9114),
.Y(net6543)
);

AO211x2_ASAP7_75t_R c6483(
.A1(net6531),
.A2(net5691),
.B(net5574),
.C(net3825),
.Y(net6544)
);

BUFx24_ASAP7_75t_R c6484(
.A(net6485),
.Y(net6545)
);

BUFx2_ASAP7_75t_R c6485(
.A(net10576),
.Y(net6546)
);

BUFx3_ASAP7_75t_R c6486(
.A(net6537),
.Y(net6547)
);

NOR2x1p5_ASAP7_75t_R c6487(
.A(net6460),
.B(net6506),
.Y(net6548)
);

NOR2x2_ASAP7_75t_R c6488(
.A(net4716),
.B(net5576),
.Y(net6549)
);

BUFx4_ASAP7_75t_R c6489(
.A(net5681),
.Y(net6550)
);

BUFx4f_ASAP7_75t_R c6490(
.A(net6455),
.Y(net6551)
);

BUFx5_ASAP7_75t_R c6491(
.A(net5670),
.Y(net6552)
);

BUFx6f_ASAP7_75t_R c6492(
.A(net6541),
.Y(net6553)
);

BUFx8_ASAP7_75t_R c6493(
.A(net6548),
.Y(net6554)
);

CKINVDCx10_ASAP7_75t_R c6494(
.A(net6536),
.Y(net6555)
);

CKINVDCx11_ASAP7_75t_R c6495(
.A(net6540),
.Y(net6556)
);

CKINVDCx12_ASAP7_75t_R c6496(
.A(net6546),
.Y(net6557)
);

NOR2xp33_ASAP7_75t_R c6497(
.A(net5551),
.B(net5541),
.Y(net6558)
);

CKINVDCx14_ASAP7_75t_R c6498(
.A(net6538),
.Y(net6559)
);

CKINVDCx16_ASAP7_75t_R c6499(
.A(net6491),
.Y(net6560)
);

NOR2xp67_ASAP7_75t_R c6500(
.A(net4740),
.B(net5638),
.Y(net6561)
);

OR2x2_ASAP7_75t_R c6501(
.A(net6558),
.B(net5618),
.Y(net6562)
);

NAND3xp33_ASAP7_75t_R c6502(
.A(net6466),
.B(net6536),
.C(net6534),
.Y(net6563)
);

CKINVDCx20_ASAP7_75t_R c6503(
.A(net6553),
.Y(net6564)
);

CKINVDCx5p33_ASAP7_75t_R c6504(
.A(net6543),
.Y(net6565)
);

CKINVDCx6p67_ASAP7_75t_R c6505(
.A(net6534),
.Y(net6566)
);

NOR3x1_ASAP7_75t_R c6506(
.A(net6514),
.B(net4724),
.C(net6550),
.Y(net6567)
);

OR2x4_ASAP7_75t_R c6507(
.A(net6545),
.B(net5551),
.Y(net6568)
);

CKINVDCx8_ASAP7_75t_R c6508(
.A(net6497),
.Y(net6569)
);

NOR3x2_ASAP7_75t_R c6509(
.B(net6551),
.C(net6567),
.A(net6563),
.Y(net6570)
);

CKINVDCx9p33_ASAP7_75t_R c6510(
.A(net6556),
.Y(net6571)
);

OR2x6_ASAP7_75t_R c6511(
.A(net3728),
.B(net4692),
.Y(net6572)
);

HB1xp67_ASAP7_75t_R c6512(
.A(net9253),
.Y(net6573)
);

NOR3xp33_ASAP7_75t_R c6513(
.A(net6541),
.B(net6558),
.C(net6554),
.Y(net6574)
);

AO22x1_ASAP7_75t_R c6514(
.A1(net6564),
.A2(net5638),
.B1(net6565),
.B2(net10219),
.Y(net6575)
);

HB2xp67_ASAP7_75t_R c6515(
.A(net6552),
.Y(net6576)
);

XNOR2x1_ASAP7_75t_R c6516(
.B(net6570),
.A(net6561),
.Y(net6577)
);

HB3xp67_ASAP7_75t_R c6517(
.A(net6539),
.Y(net6578)
);

XNOR2x2_ASAP7_75t_R c6518(
.A(net968),
.B(net9698),
.Y(net6579)
);

HB4xp67_ASAP7_75t_R c6519(
.A(net6551),
.Y(net6580)
);

XNOR2xp5_ASAP7_75t_R c6520(
.A(net4616),
.B(net6565),
.Y(net6581)
);

XOR2x1_ASAP7_75t_R c6521(
.A(net4692),
.B(net6553),
.Y(net6582)
);

INVx11_ASAP7_75t_R c6522(
.A(net9963),
.Y(net6583)
);

INVx13_ASAP7_75t_R c6523(
.A(net10557),
.Y(net6584)
);

OA21x2_ASAP7_75t_R c6524(
.A1(net6582),
.A2(net5620),
.B(net6581),
.Y(net6585)
);

INVx1_ASAP7_75t_R c6525(
.A(net6573),
.Y(net6586)
);

OAI21x1_ASAP7_75t_R c6526(
.A1(net6458),
.A2(net4732),
.B(net6583),
.Y(net6587)
);

XOR2x2_ASAP7_75t_R c6527(
.A(net6506),
.B(net9818),
.Y(net6588)
);

XOR2xp5_ASAP7_75t_R c6528(
.A(net5615),
.B(net6565),
.Y(net6589)
);

AND2x2_ASAP7_75t_R c6529(
.A(net6566),
.B(net6560),
.Y(net6590)
);

INVx2_ASAP7_75t_R c6530(
.A(net10501),
.Y(net6591)
);

AND2x4_ASAP7_75t_R c6531(
.A(net6565),
.B(net6583),
.Y(net6592)
);

AO22x2_ASAP7_75t_R c6532(
.A1(net6591),
.A2(net6575),
.B1(net6590),
.B2(net2811),
.Y(net6593)
);

AND2x6_ASAP7_75t_R c6533(
.A(net6590),
.B(net10277),
.Y(net6594)
);

INVx3_ASAP7_75t_R c6534(
.A(net10278),
.Y(net6595)
);

HAxp5_ASAP7_75t_R c6535(
.A(net6579),
.B(net6594),
.CON(net6597),
.SN(net6596)
);

INVx4_ASAP7_75t_R c6536(
.A(net6583),
.Y(net6598)
);

NAND2x1_ASAP7_75t_R c6537(
.A(net6594),
.B(net4661),
.Y(net6599)
);

NAND2x1p5_ASAP7_75t_R c6538(
.A(net6571),
.B(net6596),
.Y(net6600)
);

NAND2x2_ASAP7_75t_R c6539(
.A(net6587),
.B(net6491),
.Y(net6601)
);

AO31x2_ASAP7_75t_R c6540(
.A1(net6588),
.A2(net6545),
.A3(net6600),
.B(net10279),
.Y(net6602)
);

OR5x2_ASAP7_75t_R c6541(
.A(net6597),
.B(net6553),
.C(net6583),
.D(net6600),
.E(net10279),
.Y(net6603)
);

OAI21xp33_ASAP7_75t_R c6542(
.A1(net6580),
.A2(net5618),
.B(net6601),
.Y(net6604)
);

INVx5_ASAP7_75t_R c6543(
.A(net10405),
.Y(net6605)
);

A2O1A1O1Ixp25_ASAP7_75t_R c6544(
.A1(net6603),
.A2(net6599),
.B(net6548),
.C(net6600),
.D(net5689),
.Y(net6606)
);

SDFHx1_ASAP7_75t_R c6545(
.D(net6604),
.SE(net4692),
.SI(net6561),
.CLK(clk),
.QN(net6607)
);

OAI21xp5_ASAP7_75t_R c6546(
.A1(net6584),
.A2(net6607),
.B(net6592),
.Y(net6608)
);

OR3x1_ASAP7_75t_R c6547(
.A(net5610),
.B(net6535),
.C(net9698),
.Y(net6609)
);

INVx6_ASAP7_75t_R c6548(
.A(net10412),
.Y(net6610)
);

NAND2xp33_ASAP7_75t_R c6549(
.A(net5676),
.B(net6595),
.Y(net6611)
);

NAND2xp5_ASAP7_75t_R c6550(
.A(net6607),
.B(net6537),
.Y(net6612)
);

NAND2xp67_ASAP7_75t_R c6551(
.A(net6599),
.B(net9830),
.Y(net6613)
);

OR3x2_ASAP7_75t_R c6552(
.A(net6559),
.B(net6582),
.C(net6569),
.Y(net6614)
);

ICGx6p67DC_ASAP7_75t_R c6553(
.ENA(net6614),
.SE(net9766),
.CLK(clk),
.GCLK(net6615)
);

NOR2x1_ASAP7_75t_R c6554(
.A(net6608),
.B(net6615),
.Y(net6616)
);

AND5x1_ASAP7_75t_R c6555(
.A(net6592),
.B(net6610),
.C(net6614),
.D(net6569),
.E(net6608),
.Y(net6617)
);

AO33x2_ASAP7_75t_R c6556(
.A1(net6610),
.A2(net6565),
.A3(net6608),
.B1(net6616),
.B2(net6612),
.B3(net4738),
.Y(net6618)
);

INVx8_ASAP7_75t_R c6557(
.A(net5735),
.Y(net6619)
);

INVxp33_ASAP7_75t_R c6558(
.A(net4650),
.Y(net6620)
);

INVxp67_ASAP7_75t_R c6559(
.A(net10096),
.Y(net6621)
);

BUFx10_ASAP7_75t_R c6560(
.A(net6555),
.Y(net6622)
);

BUFx12_ASAP7_75t_R c6561(
.A(net9719),
.Y(net6623)
);

NOR2x1p5_ASAP7_75t_R c6562(
.A(net6473),
.B(net6600),
.Y(net6624)
);

NOR2x2_ASAP7_75t_R c6563(
.A(net6586),
.B(net6569),
.Y(net6625)
);

NOR2xp33_ASAP7_75t_R c6564(
.A(net6611),
.B(net4681),
.Y(net6626)
);

NOR2xp67_ASAP7_75t_R c6565(
.A(net6589),
.B(net5763),
.Y(net6627)
);

BUFx12f_ASAP7_75t_R c6566(
.A(net5751),
.Y(net6628)
);

BUFx16f_ASAP7_75t_R c6567(
.A(net9186),
.Y(net6629)
);

OR2x2_ASAP7_75t_R c6568(
.A(net4846),
.B(net6629),
.Y(net6630)
);

BUFx24_ASAP7_75t_R c6569(
.A(net10093),
.Y(net6631)
);

BUFx2_ASAP7_75t_R c6570(
.A(net6628),
.Y(net6632)
);

OR2x4_ASAP7_75t_R c6571(
.A(net6619),
.B(net6625),
.Y(net6633)
);

BUFx3_ASAP7_75t_R c6572(
.A(net5638),
.Y(net6634)
);

OR2x6_ASAP7_75t_R c6573(
.A(net6634),
.B(net9800),
.Y(net6635)
);

XNOR2x1_ASAP7_75t_R c6574(
.B(net5625),
.A(net2963),
.Y(net6636)
);

OR3x4_ASAP7_75t_R c6575(
.A(net6636),
.B(net6634),
.C(net4849),
.Y(net6637)
);

XNOR2x2_ASAP7_75t_R c6576(
.A(net5770),
.B(net6561),
.Y(net6638)
);

BUFx4_ASAP7_75t_R c6577(
.A(net4856),
.Y(net6639)
);

AND3x1_ASAP7_75t_R c6578(
.A(net6637),
.B(net6620),
.C(net10279),
.Y(net6640)
);

BUFx4f_ASAP7_75t_R c6579(
.A(net9186),
.Y(net6641)
);

AND3x2_ASAP7_75t_R c6580(
.A(net4849),
.B(net6634),
.C(net6542),
.Y(net6642)
);

ICGx8DC_ASAP7_75t_R c6581(
.ENA(net6624),
.SE(net10052),
.CLK(clk),
.GCLK(net6643)
);

AND3x4_ASAP7_75t_R c6582(
.A(net2754),
.B(net3767),
.C(net6601),
.Y(net6644)
);

BUFx5_ASAP7_75t_R c6583(
.A(net5742),
.Y(net6645)
);

XNOR2xp5_ASAP7_75t_R c6584(
.A(net3804),
.B(net5775),
.Y(net6646)
);

XOR2x1_ASAP7_75t_R c6585(
.A(net6590),
.B(net6589),
.Y(net6647)
);

BUFx6f_ASAP7_75t_R c6586(
.A(net10449),
.Y(net6648)
);

XOR2x2_ASAP7_75t_R c6587(
.A(net6601),
.B(net3804),
.Y(net6649)
);

XOR2xp5_ASAP7_75t_R c6588(
.A(net5766),
.B(net6646),
.Y(net6650)
);

BUFx8_ASAP7_75t_R c6589(
.A(net9207),
.Y(net6651)
);

CKINVDCx10_ASAP7_75t_R c6590(
.A(net6632),
.Y(net6652)
);

AND2x2_ASAP7_75t_R c6591(
.A(net5696),
.B(net5772),
.Y(net6653)
);

SDFHx2_ASAP7_75t_R c6592(
.D(net5704),
.SE(net6600),
.SI(net5638),
.CLK(clk),
.QN(net6654)
);

AND2x4_ASAP7_75t_R c6593(
.A(net6563),
.B(net6625),
.Y(net6655)
);

AND2x6_ASAP7_75t_R c6594(
.A(net6654),
.B(net6631),
.Y(net6656)
);

AO21x1_ASAP7_75t_R c6595(
.A1(net5741),
.A2(net6616),
.B(net2754),
.Y(net6657)
);

CKINVDCx11_ASAP7_75t_R c6596(
.A(net10165),
.Y(net6658)
);

HAxp5_ASAP7_75t_R c6597(
.A(net6576),
.B(net6652),
.CON(net6659)
);

CKINVDCx12_ASAP7_75t_R c6598(
.A(net6581),
.Y(net6660)
);

AO21x2_ASAP7_75t_R c6599(
.A1(net5774),
.A2(net6627),
.B(net6654),
.Y(net6661)
);

AOI21x1_ASAP7_75t_R c6600(
.A1(net6653),
.A2(net6625),
.B(net10052),
.Y(net6662)
);

CKINVDCx14_ASAP7_75t_R c6601(
.A(net10404),
.Y(net6663)
);

AOI21xp33_ASAP7_75t_R c6602(
.A1(net6648),
.A2(net5766),
.B(net6618),
.Y(net6664)
);

NAND2x1_ASAP7_75t_R c6603(
.A(net6642),
.B(net9675),
.Y(net6665)
);

NAND2x1p5_ASAP7_75t_R c6604(
.A(net6613),
.B(net6635),
.Y(net6666)
);

SDFHx3_ASAP7_75t_R c6605(
.D(net6627),
.SE(net6629),
.SI(net6660),
.CLK(clk),
.QN(net6667)
);

CKINVDCx16_ASAP7_75t_R c6606(
.A(net6634),
.Y(net6668)
);

CKINVDCx20_ASAP7_75t_R c6607(
.A(net10116),
.Y(net6669)
);

CKINVDCx5p33_ASAP7_75t_R c6608(
.A(net9193),
.Y(net6670)
);

NAND2x2_ASAP7_75t_R c6609(
.A(net6659),
.B(net6655),
.Y(net6671)
);

NAND2xp33_ASAP7_75t_R c6610(
.A(net6662),
.B(net6669),
.Y(net6672)
);

CKINVDCx6p67_ASAP7_75t_R c6611(
.A(net6655),
.Y(net6673)
);

AOI21xp5_ASAP7_75t_R c6612(
.A1(net6452),
.A2(net6667),
.B(net6669),
.Y(net6674)
);

CKINVDCx8_ASAP7_75t_R c6613(
.A(net6664),
.Y(net6675)
);

NAND2xp5_ASAP7_75t_R c6614(
.A(net6648),
.B(net9827),
.Y(net6676)
);

NAND2xp67_ASAP7_75t_R c6615(
.A(net6622),
.B(net5770),
.Y(net6677)
);

FAx1_ASAP7_75t_R c6616(
.A(net6675),
.B(net3878),
.CI(net6646),
.SN(net6679),
.CON(net6678)
);

CKINVDCx9p33_ASAP7_75t_R c6617(
.A(net10093),
.Y(net6680)
);

MAJIxp5_ASAP7_75t_R c6618(
.A(net5767),
.B(net6654),
.C(net5718),
.Y(net6681)
);

MAJx2_ASAP7_75t_R c6619(
.A(net6674),
.B(net6655),
.C(net6669),
.Y(net6682)
);

NOR2x1_ASAP7_75t_R c6620(
.A(net6626),
.B(net6677),
.Y(net6683)
);

NOR2x1p5_ASAP7_75t_R c6621(
.A(net6672),
.B(net6595),
.Y(net6684)
);

NOR2x2_ASAP7_75t_R c6622(
.A(net6677),
.B(net6664),
.Y(net6685)
);

NOR2xp33_ASAP7_75t_R c6623(
.A(net6660),
.B(net5770),
.Y(net6686)
);

AOI211x1_ASAP7_75t_R c6624(
.A1(net6656),
.A2(net6679),
.B(net6577),
.C(net6508),
.Y(net6687)
);

HB1xp67_ASAP7_75t_R c6625(
.A(net10458),
.Y(net6688)
);

HB2xp67_ASAP7_75t_R c6626(
.A(net10464),
.Y(net6689)
);

MAJx3_ASAP7_75t_R c6627(
.A(net6671),
.B(net6674),
.C(net6636),
.Y(net6690)
);

HB3xp67_ASAP7_75t_R c6628(
.A(net10449),
.Y(net6691)
);

ICGx1_ASAP7_75t_R c6629(
.ENA(net6683),
.SE(net6667),
.CLK(clk),
.GCLK(net6692)
);

HB4xp67_ASAP7_75t_R c6630(
.A(net10507),
.Y(net6693)
);

NAND3x1_ASAP7_75t_R c6631(
.A(net6631),
.B(net6692),
.C(net5660),
.Y(net6694)
);

NAND3x2_ASAP7_75t_R c6632(
.B(net6650),
.C(net6673),
.A(net6681),
.Y(net6695)
);

NOR2xp67_ASAP7_75t_R c6633(
.A(net4783),
.B(net6695),
.Y(net6696)
);

INVx11_ASAP7_75t_R c6634(
.A(net10434),
.Y(net6697)
);

NAND3xp33_ASAP7_75t_R c6635(
.A(net6689),
.B(net6684),
.C(net5657),
.Y(net6698)
);

OR2x2_ASAP7_75t_R c6636(
.A(net6697),
.B(net6663),
.Y(net6699)
);

SDFHx4_ASAP7_75t_R c6637(
.D(net6699),
.SE(net6665),
.SI(net6651),
.CLK(clk),
.QN(net6700)
);

OR2x4_ASAP7_75t_R c6638(
.A(net6673),
.B(net6700),
.Y(net6701)
);

AOI222xp33_ASAP7_75t_R c6639(
.A1(net6693),
.A2(net6690),
.B1(net6699),
.B2(net6700),
.C1(net6701),
.C2(net6643),
.Y(net6702)
);

INVx13_ASAP7_75t_R c6640(
.A(net10474),
.Y(net6703)
);

OR2x6_ASAP7_75t_R c6641(
.A(net5807),
.B(net5819),
.Y(net6704)
);

XNOR2x1_ASAP7_75t_R c6642(
.B(net6641),
.A(net5848),
.Y(net6705)
);

XNOR2x2_ASAP7_75t_R c6643(
.A(net5802),
.B(net6685),
.Y(net6706)
);

XNOR2xp5_ASAP7_75t_R c6644(
.A(net6658),
.B(net10164),
.Y(net6707)
);

XOR2x1_ASAP7_75t_R c6645(
.A(net5776),
.B(net6482),
.Y(net6708)
);

XOR2x2_ASAP7_75t_R c6646(
.A(net5839),
.B(net5775),
.Y(net6709)
);

XOR2xp5_ASAP7_75t_R c6647(
.A(net4933),
.B(net6618),
.Y(net6710)
);

INVx1_ASAP7_75t_R c6648(
.A(net10164),
.Y(net6711)
);

AND2x2_ASAP7_75t_R c6649(
.A(net4905),
.B(net5796),
.Y(net6712)
);

INVx2_ASAP7_75t_R c6650(
.A(net6623),
.Y(net6713)
);

ICGx2_ASAP7_75t_R c6651(
.ENA(net6704),
.SE(net5780),
.CLK(clk),
.GCLK(net6714)
);

INVx3_ASAP7_75t_R c6652(
.A(net3054),
.Y(net6715)
);

AND2x4_ASAP7_75t_R c6653(
.A(net5757),
.B(net3984),
.Y(net6716)
);

INVx4_ASAP7_75t_R c6654(
.A(net10379),
.Y(net6717)
);

NOR3x1_ASAP7_75t_R c6655(
.A(net4788),
.B(net6695),
.C(net3015),
.Y(net6718)
);

AND2x6_ASAP7_75t_R c6656(
.A(net5836),
.B(net10028),
.Y(net6719)
);

HAxp5_ASAP7_75t_R c6657(
.A(net5819),
.B(net6706),
.CON(net6720)
);

SDFLx1_ASAP7_75t_R c6658(
.D(net6578),
.SE(net6577),
.SI(net5775),
.CLK(clk),
.QN(net6721)
);

NAND2x1_ASAP7_75t_R c6659(
.A(net6713),
.B(net5793),
.Y(net6722)
);

NAND2x1p5_ASAP7_75t_R c6660(
.A(net4877),
.B(net6642),
.Y(net6723)
);

NAND2x2_ASAP7_75t_R c6661(
.A(net6504),
.B(net6621),
.Y(net6724)
);

NAND2xp33_ASAP7_75t_R c6662(
.A(net5779),
.B(net10085),
.Y(net6725)
);

NAND2xp5_ASAP7_75t_R c6663(
.A(net6577),
.B(net6451),
.Y(net6726)
);

INVx5_ASAP7_75t_R c6664(
.A(net10164),
.Y(net6727)
);

INVx6_ASAP7_75t_R c6665(
.A(net10431),
.Y(net6728)
);

NOR3x2_ASAP7_75t_R c6666(
.B(net6621),
.C(net6723),
.A(net6658),
.Y(net6729)
);

INVx8_ASAP7_75t_R c6667(
.A(net10020),
.Y(net6730)
);

INVxp33_ASAP7_75t_R c6668(
.A(net5810),
.Y(net6731)
);

NAND2xp67_ASAP7_75t_R c6669(
.A(net3059),
.B(net3942),
.Y(net6732)
);

INVxp67_ASAP7_75t_R c6670(
.A(net10128),
.Y(net6733)
);

NOR2x1_ASAP7_75t_R c6671(
.A(net6695),
.B(net4905),
.Y(net6734)
);

NOR2x1p5_ASAP7_75t_R c6672(
.A(net6577),
.B(net9841),
.Y(net6735)
);

NOR2x2_ASAP7_75t_R c6673(
.A(net5763),
.B(net6598),
.Y(net6736)
);

NOR2xp33_ASAP7_75t_R c6674(
.A(net6717),
.B(net6730),
.Y(net6737)
);

NOR2xp67_ASAP7_75t_R c6675(
.A(net6727),
.B(net5839),
.Y(net6738)
);

OR2x2_ASAP7_75t_R c6676(
.A(net6700),
.B(net5788),
.Y(net6739)
);

NOR3xp33_ASAP7_75t_R c6677(
.A(net6652),
.B(net6705),
.C(net6733),
.Y(net6740)
);

OR2x4_ASAP7_75t_R c6678(
.A(net5541),
.B(net6723),
.Y(net6741)
);

OR2x6_ASAP7_75t_R c6679(
.A(net5748),
.B(net6708),
.Y(net6742)
);

OA21x2_ASAP7_75t_R c6680(
.A1(net5810),
.A2(net6649),
.B(net10269),
.Y(net6743)
);

BUFx10_ASAP7_75t_R c6681(
.A(net10410),
.Y(net6744)
);

OAI21x1_ASAP7_75t_R c6682(
.A1(net6731),
.A2(net6709),
.B(net6700),
.Y(net6745)
);

XNOR2x1_ASAP7_75t_R c6683(
.B(net5780),
.A(net4788),
.Y(net6746)
);

XNOR2x2_ASAP7_75t_R c6684(
.A(net5711),
.B(net6707),
.Y(net6747)
);

OAI21xp33_ASAP7_75t_R c6685(
.A1(net6715),
.A2(net6621),
.B(net9881),
.Y(net6748)
);

BUFx12_ASAP7_75t_R c6686(
.A(net10474),
.Y(net6749)
);

XNOR2xp5_ASAP7_75t_R c6687(
.A(net6651),
.B(net950),
.Y(net6750)
);

ICGx2p67DC_ASAP7_75t_R c6688(
.ENA(net6598),
.SE(net6679),
.CLK(clk),
.GCLK(net6751)
);

BUFx12f_ASAP7_75t_R c6689(
.A(net10379),
.Y(net6752)
);

XOR2x1_ASAP7_75t_R c6690(
.A(net6744),
.B(net6732),
.Y(net6753)
);

SDFLx2_ASAP7_75t_R c6691(
.D(net6752),
.SE(net6747),
.SI(net10264),
.CLK(clk),
.QN(net6754)
);

XOR2x2_ASAP7_75t_R c6692(
.A(net6638),
.B(net6692),
.Y(net6755)
);

XOR2xp5_ASAP7_75t_R c6693(
.A(net6754),
.B(net6714),
.Y(net6756)
);

AND2x2_ASAP7_75t_R c6694(
.A(net6733),
.B(net9769),
.Y(net6757)
);

AND2x4_ASAP7_75t_R c6695(
.A(net6639),
.B(net6755),
.Y(net6758)
);

AND2x6_ASAP7_75t_R c6696(
.A(net6748),
.B(net10134),
.Y(net6759)
);

HAxp5_ASAP7_75t_R c6697(
.A(net6757),
.B(net6710),
.CON(net6761),
.SN(net6760)
);

AOI211xp5_ASAP7_75t_R c6698(
.A1(net5804),
.A2(net6752),
.B(net3984),
.C(net4911),
.Y(net6762)
);

NAND2x1_ASAP7_75t_R c6699(
.A(net6746),
.B(net10280),
.Y(net6763)
);

NAND2x1p5_ASAP7_75t_R c6700(
.A(net6756),
.B(net9845),
.Y(net6764)
);

OAI21xp5_ASAP7_75t_R c6701(
.A1(net6750),
.A2(net6709),
.B(net9826),
.Y(net6765)
);

NAND2x2_ASAP7_75t_R c6702(
.A(net5853),
.B(net6748),
.Y(net6766)
);

NAND2xp33_ASAP7_75t_R c6703(
.A(net6722),
.B(net5772),
.Y(net6767)
);

OR3x1_ASAP7_75t_R c6704(
.A(net6645),
.B(net6763),
.C(net6747),
.Y(net6768)
);

NAND2xp5_ASAP7_75t_R c6705(
.A(net5796),
.B(net6742),
.Y(net6769)
);

NAND2xp67_ASAP7_75t_R c6706(
.A(net9867),
.B(net10280),
.Y(net6770)
);

NOR2x1_ASAP7_75t_R c6707(
.A(net6769),
.B(net4732),
.Y(net6771)
);

NOR2x1p5_ASAP7_75t_R c6708(
.A(net6770),
.B(net5839),
.Y(net6772)
);

NOR2x2_ASAP7_75t_R c6709(
.A(net6703),
.B(net4940),
.Y(net6773)
);

NOR2xp33_ASAP7_75t_R c6710(
.A(net5656),
.B(net6767),
.Y(net6774)
);

AOI22x1_ASAP7_75t_R c6711(
.A1(net6740),
.A2(net6767),
.B1(net6748),
.B2(net5839),
.Y(net6775)
);

NOR2xp67_ASAP7_75t_R c6712(
.A(net6750),
.B(net6703),
.Y(net6776)
);

SDFLx3_ASAP7_75t_R c6713(
.D(net6776),
.SE(net6732),
.SI(net6755),
.CLK(clk),
.QN(net6777)
);

OR3x2_ASAP7_75t_R c6714(
.A(net5793),
.B(net6721),
.C(net10158),
.Y(net6778)
);

OR2x2_ASAP7_75t_R c6715(
.A(net3942),
.B(net6748),
.Y(net6779)
);

OR3x4_ASAP7_75t_R c6716(
.A(net6756),
.B(net6779),
.C(net10158),
.Y(net6780)
);

AND3x1_ASAP7_75t_R c6717(
.A(net6778),
.B(net6749),
.C(net9881),
.Y(net6781)
);

OR2x4_ASAP7_75t_R c6718(
.A(net6712),
.B(net6700),
.Y(net6782)
);

OR2x6_ASAP7_75t_R c6719(
.A(net5660),
.B(net6778),
.Y(net6783)
);

AND3x2_ASAP7_75t_R c6720(
.A(net6779),
.B(net6765),
.C(net6774),
.Y(net6784)
);

AOI321xp33_ASAP7_75t_R c6721(
.A1(net6778),
.A2(net6754),
.A3(net6666),
.B1(net6748),
.B2(net5657),
.C(net9769),
.Y(net6785)
);

XNOR2x1_ASAP7_75t_R c6722(
.B(net6783),
.A(net9932),
.Y(net6786)
);

BUFx16f_ASAP7_75t_R c6723(
.A(net6736),
.Y(net6787)
);

BUFx24_ASAP7_75t_R c6724(
.A(net6786),
.Y(net6788)
);

XNOR2x2_ASAP7_75t_R c6725(
.A(net6725),
.B(net5006),
.Y(net6789)
);

AOI22xp33_ASAP7_75t_R c6726(
.A1(net6670),
.A2(net6701),
.B1(net5006),
.B2(net5931),
.Y(net6790)
);

XNOR2xp5_ASAP7_75t_R c6727(
.A(net6774),
.B(net5942),
.Y(net6791)
);

BUFx2_ASAP7_75t_R c6728(
.A(net6692),
.Y(net6792)
);

AOI22xp5_ASAP7_75t_R c6729(
.A1(net5747),
.A2(net4951),
.B1(net6791),
.B2(net10130),
.Y(net6793)
);

SDFLx4_ASAP7_75t_R c6730(
.D(net5925),
.SE(net6763),
.SI(net5866),
.CLK(clk),
.QN(net6794)
);

XOR2x1_ASAP7_75t_R c6731(
.A(net5891),
.B(net6670),
.Y(net6795)
);

XOR2x2_ASAP7_75t_R c6732(
.A(net6685),
.B(net5942),
.Y(net6796)
);

BUFx3_ASAP7_75t_R c6733(
.A(net4971),
.Y(net6797)
);

BUFx4_ASAP7_75t_R c6734(
.A(net10475),
.Y(net6798)
);

XOR2xp5_ASAP7_75t_R c6735(
.A(net5618),
.B(net6791),
.Y(net6799)
);

BUFx4f_ASAP7_75t_R c6736(
.A(net10280),
.Y(net6800)
);

AND2x2_ASAP7_75t_R c6737(
.A(net5920),
.B(net10254),
.Y(net6801)
);

BUFx5_ASAP7_75t_R c6738(
.A(net6763),
.Y(net6802)
);

BUFx6f_ASAP7_75t_R c6739(
.A(net9097),
.Y(net6803)
);

BUFx8_ASAP7_75t_R c6740(
.A(net10574),
.Y(net6804)
);

AND2x4_ASAP7_75t_R c6741(
.A(net6797),
.B(net6721),
.Y(net6805)
);

AND2x6_ASAP7_75t_R c6742(
.A(net5006),
.B(net5926),
.Y(net6806)
);

ICGx3_ASAP7_75t_R c6743(
.ENA(net6752),
.SE(net6791),
.CLK(clk),
.GCLK(net6807)
);

AND3x4_ASAP7_75t_R c6744(
.A(net6759),
.B(net4835),
.C(net10281),
.Y(net6808)
);

HAxp5_ASAP7_75t_R c6745(
.A(net6618),
.B(net10255),
.CON(net6809)
);

CKINVDCx10_ASAP7_75t_R c6746(
.A(net10145),
.Y(net6810)
);

CKINVDCx11_ASAP7_75t_R c6747(
.A(net10391),
.Y(net6811)
);

NAND2x1_ASAP7_75t_R c6748(
.A(net5932),
.B(net10032),
.Y(net6812)
);

NAND2x1p5_ASAP7_75t_R c6749(
.A(net5918),
.B(net10281),
.Y(net6813)
);

AO21x1_ASAP7_75t_R c6750(
.A1(net6724),
.A2(net5879),
.B(net6794),
.Y(net6814)
);

CKINVDCx12_ASAP7_75t_R c6751(
.A(net6767),
.Y(net6815)
);

NAND2x2_ASAP7_75t_R c6752(
.A(net6800),
.B(net10190),
.Y(net6816)
);

CKINVDCx14_ASAP7_75t_R c6753(
.A(net10531),
.Y(net6817)
);

CKINVDCx16_ASAP7_75t_R c6754(
.A(net10555),
.Y(net6818)
);

CKINVDCx20_ASAP7_75t_R c6755(
.A(net6807),
.Y(net6819)
);

NAND2xp33_ASAP7_75t_R c6756(
.A(net6805),
.B(net5891),
.Y(net6820)
);

CKINVDCx5p33_ASAP7_75t_R c6757(
.A(net5797),
.Y(net6821)
);

NAND2xp5_ASAP7_75t_R c6758(
.A(net6721),
.B(net6815),
.Y(net6822)
);

CKINVDCx6p67_ASAP7_75t_R c6759(
.A(net10103),
.Y(net6823)
);

NAND2xp67_ASAP7_75t_R c6760(
.A(net6821),
.B(net6814),
.Y(net6824)
);

CKINVDCx8_ASAP7_75t_R c6761(
.A(net6817),
.Y(net6825)
);

NOR2x1_ASAP7_75t_R c6762(
.A(net4032),
.B(net1078),
.Y(net6826)
);

CKINVDCx9p33_ASAP7_75t_R c6763(
.A(net10266),
.Y(net6827)
);

HB1xp67_ASAP7_75t_R c6764(
.A(net6826),
.Y(net6828)
);

HB2xp67_ASAP7_75t_R c6765(
.A(net4064),
.Y(net6829)
);

HB3xp67_ASAP7_75t_R c6766(
.A(net6775),
.Y(net6830)
);

NOR2x1p5_ASAP7_75t_R c6767(
.A(net6812),
.B(net6817),
.Y(net6831)
);

DFFASRHQNx1_ASAP7_75t_R c6768(
.D(net6819),
.RESETN(net6815),
.SETN(net6791),
.CLK(clk),
.QN(net6832)
);

NOR2x2_ASAP7_75t_R c6769(
.A(net5922),
.B(net3707),
.Y(net6833)
);

NOR2xp33_ASAP7_75t_R c6770(
.A(net6818),
.B(net5858),
.Y(net6834)
);

NOR2xp67_ASAP7_75t_R c6771(
.A(net6824),
.B(net6710),
.Y(net6835)
);

OR2x2_ASAP7_75t_R c6772(
.A(net5931),
.B(net6751),
.Y(net6836)
);

OR2x4_ASAP7_75t_R c6773(
.A(net6833),
.B(net5797),
.Y(net6837)
);

AO21x2_ASAP7_75t_R c6774(
.A1(net6810),
.A2(net5940),
.B(net6692),
.Y(net6838)
);

HB4xp67_ASAP7_75t_R c6775(
.A(net4911),
.Y(net6839)
);

INVx11_ASAP7_75t_R c6776(
.A(net9097),
.Y(net6840)
);

AOI21x1_ASAP7_75t_R c6777(
.A1(net6823),
.A2(net6789),
.B(net6802),
.Y(net6841)
);

AOI21xp33_ASAP7_75t_R c6778(
.A1(net6834),
.A2(net6833),
.B(net6774),
.Y(net6842)
);

OR2x6_ASAP7_75t_R c6779(
.A(net6839),
.B(net6707),
.Y(net6843)
);

XNOR2x1_ASAP7_75t_R c6780(
.B(net6685),
.A(net9936),
.Y(net6844)
);

XNOR2x2_ASAP7_75t_R c6781(
.A(net6787),
.B(net9731),
.Y(net6845)
);

XNOR2xp5_ASAP7_75t_R c6782(
.A(net5893),
.B(net6839),
.Y(net6846)
);

INVx13_ASAP7_75t_R c6783(
.A(net10369),
.Y(net6847)
);

INVx1_ASAP7_75t_R c6784(
.A(net10094),
.Y(net6848)
);

INVx2_ASAP7_75t_R c6785(
.A(net6813),
.Y(net6849)
);

XOR2x1_ASAP7_75t_R c6786(
.A(net6828),
.B(net4953),
.Y(net6850)
);

SDFHx1_ASAP7_75t_R c6787(
.D(net6820),
.SE(net6807),
.SI(net6789),
.CLK(clk),
.QN(net6851)
);

INVx3_ASAP7_75t_R c6788(
.A(net10401),
.Y(net6852)
);

INVx4_ASAP7_75t_R c6789(
.A(net10359),
.Y(net6853)
);

AOI21xp5_ASAP7_75t_R c6790(
.A1(net6822),
.A2(net6844),
.B(net5618),
.Y(net6854)
);

XOR2x2_ASAP7_75t_R c6791(
.A(net6839),
.B(net9778),
.Y(net6855)
);

FAx1_ASAP7_75t_R c6792(
.A(net6829),
.B(net6835),
.CI(net4930),
.SN(net6857),
.CON(net6856)
);

XOR2xp5_ASAP7_75t_R c6793(
.A(net6848),
.B(net6787),
.Y(net6858)
);

INVx5_ASAP7_75t_R c6794(
.A(net10565),
.Y(net6859)
);

AND5x2_ASAP7_75t_R c6795(
.A(net6842),
.B(net6858),
.C(net6848),
.D(net6791),
.E(net10281),
.Y(net6860)
);

INVx6_ASAP7_75t_R c6796(
.A(net9193),
.Y(net6861)
);

AOI33xp33_ASAP7_75t_R c6797(
.A1(net6858),
.A2(net6857),
.A3(net6836),
.B1(net5609),
.B2(net4962),
.B3(net6791),
.Y(net6862)
);

AOI31xp33_ASAP7_75t_R c6798(
.A1(net5882),
.A2(net6821),
.A3(net6839),
.B(net10283),
.Y(net6863)
);

AND2x2_ASAP7_75t_R c6799(
.A(net5907),
.B(net6846),
.Y(net6864)
);

MAJIxp5_ASAP7_75t_R c6800(
.A(net6811),
.B(net6861),
.C(net6858),
.Y(net6865)
);

AND2x4_ASAP7_75t_R c6801(
.A(net6849),
.B(net6851),
.Y(net6866)
);

MAJx2_ASAP7_75t_R c6802(
.A(net5940),
.B(net6866),
.C(net6864),
.Y(net6867)
);

MAJx3_ASAP7_75t_R c6803(
.A(net6865),
.B(net6861),
.C(net10282),
.Y(net6868)
);

NAND3x1_ASAP7_75t_R c6804(
.A(net6831),
.B(net6865),
.C(net6832),
.Y(net6869)
);

OA222x2_ASAP7_75t_R c6805(
.A1(net6853),
.A2(net6827),
.B1(net6869),
.B2(net6868),
.C1(net6832),
.C2(net6749),
.Y(net6870)
);

INVx8_ASAP7_75t_R c6806(
.A(net5697),
.Y(net6871)
);

AND2x6_ASAP7_75t_R c6807(
.A(net5992),
.B(net6852),
.Y(net6872)
);

INVxp33_ASAP7_75t_R c6808(
.A(net4104),
.Y(net6873)
);

INVxp67_ASAP7_75t_R c6809(
.A(net10464),
.Y(net6874)
);

BUFx10_ASAP7_75t_R c6810(
.A(net9132),
.Y(net6875)
);

HAxp5_ASAP7_75t_R c6811(
.A(net4143),
.B(net6794),
.CON(net6877),
.SN(net6876)
);

NAND2x1_ASAP7_75t_R c6812(
.A(net5927),
.B(net5697),
.Y(net6878)
);

BUFx12_ASAP7_75t_R c6813(
.A(net6009),
.Y(net6879)
);

BUFx12f_ASAP7_75t_R c6814(
.A(net5775),
.Y(net6880)
);

BUFx16f_ASAP7_75t_R c6815(
.A(net6879),
.Y(net6881)
);

BUFx24_ASAP7_75t_R c6816(
.A(net5786),
.Y(net6882)
);

NAND2x1p5_ASAP7_75t_R c6817(
.A(net6880),
.B(net5982),
.Y(net6883)
);

BUFx2_ASAP7_75t_R c6818(
.A(net9132),
.Y(net6884)
);

NAND3x2_ASAP7_75t_R c6819(
.B(net6875),
.C(net5957),
.A(net5983),
.Y(net6885)
);

BUFx3_ASAP7_75t_R c6820(
.A(net10119),
.Y(net6886)
);

BUFx4_ASAP7_75t_R c6821(
.A(net6881),
.Y(net6887)
);

BUFx4f_ASAP7_75t_R c6822(
.A(net5039),
.Y(net6888)
);

BUFx5_ASAP7_75t_R c6823(
.A(net6883),
.Y(net6889)
);

BUFx6f_ASAP7_75t_R c6824(
.A(net6851),
.Y(net6890)
);

NAND3xp33_ASAP7_75t_R c6825(
.A(net2990),
.B(net6876),
.C(net5964),
.Y(net6891)
);

BUFx8_ASAP7_75t_R c6826(
.A(net6801),
.Y(net6892)
);

CKINVDCx10_ASAP7_75t_R c6827(
.A(net10282),
.Y(net6893)
);

NAND2x2_ASAP7_75t_R c6828(
.A(net6873),
.B(net6864),
.Y(net6894)
);

CKINVDCx11_ASAP7_75t_R c6829(
.A(net4174),
.Y(net6895)
);

NOR3x1_ASAP7_75t_R c6830(
.A(net6840),
.B(net6790),
.C(net6855),
.Y(net6896)
);

CKINVDCx12_ASAP7_75t_R c6831(
.A(net10548),
.Y(net6897)
);

NAND2xp33_ASAP7_75t_R c6832(
.A(net6886),
.B(net6016),
.Y(net6898)
);

CKINVDCx14_ASAP7_75t_R c6833(
.A(net6008),
.Y(net6899)
);

NAND2xp5_ASAP7_75t_R c6834(
.A(net6861),
.B(net6875),
.Y(net6900)
);

NAND2xp67_ASAP7_75t_R c6835(
.A(net6888),
.B(net6008),
.Y(net6901)
);

CKINVDCx16_ASAP7_75t_R c6836(
.A(net6893),
.Y(net6902)
);

NOR2x1_ASAP7_75t_R c6837(
.A(net6814),
.B(net6667),
.Y(net6903)
);

CKINVDCx20_ASAP7_75t_R c6838(
.A(net3872),
.Y(net6904)
);

CKINVDCx5p33_ASAP7_75t_R c6839(
.A(net5982),
.Y(net6905)
);

CKINVDCx6p67_ASAP7_75t_R c6840(
.A(net5977),
.Y(net6906)
);

NOR2x1p5_ASAP7_75t_R c6841(
.A(net6874),
.B(net10081),
.Y(net6907)
);

NOR2x2_ASAP7_75t_R c6842(
.A(net5080),
.B(net6851),
.Y(net6908)
);

CKINVDCx8_ASAP7_75t_R c6843(
.A(net6872),
.Y(net6909)
);

CKINVDCx9p33_ASAP7_75t_R c6844(
.A(net3253),
.Y(net6910)
);

NOR2xp33_ASAP7_75t_R c6845(
.A(net6910),
.B(net6861),
.Y(net6911)
);

HB1xp67_ASAP7_75t_R c6846(
.A(net10372),
.Y(net6912)
);

NOR2xp67_ASAP7_75t_R c6847(
.A(net6836),
.B(net5933),
.Y(net6913)
);

OR2x2_ASAP7_75t_R c6848(
.A(net6884),
.B(net6883),
.Y(net6914)
);

AO221x1_ASAP7_75t_R c6849(
.A1(net4931),
.A2(net6851),
.B1(net6832),
.B2(net10281),
.C(net10282),
.Y(net6915)
);

OR2x4_ASAP7_75t_R c6850(
.A(net6790),
.B(net6832),
.Y(net6916)
);

SDFHx2_ASAP7_75t_R c6851(
.D(net4138),
.SE(net5928),
.SI(net6892),
.CLK(clk),
.QN(net6917)
);

OR2x6_ASAP7_75t_R c6852(
.A(net6894),
.B(net6883),
.Y(net6918)
);

SDFHx3_ASAP7_75t_R c6853(
.D(net6794),
.SE(net5933),
.SI(net6891),
.CLK(clk),
.QN(net6919)
);

XNOR2x1_ASAP7_75t_R c6854(
.B(net6892),
.A(net6906),
.Y(net6920)
);

NOR3x2_ASAP7_75t_R c6855(
.B(net6877),
.C(net6791),
.A(net6884),
.Y(net6921)
);

HB2xp67_ASAP7_75t_R c6856(
.A(net9731),
.Y(net6922)
);

NOR3xp33_ASAP7_75t_R c6857(
.A(net6915),
.B(net5996),
.C(net6895),
.Y(net6923)
);

HB3xp67_ASAP7_75t_R c6858(
.A(net6889),
.Y(net6924)
);

XNOR2x2_ASAP7_75t_R c6859(
.A(net10099),
.B(net10281),
.Y(net6925)
);

XNOR2xp5_ASAP7_75t_R c6860(
.A(net5069),
.B(net6864),
.Y(net6926)
);

XOR2x1_ASAP7_75t_R c6861(
.A(net6707),
.B(net5968),
.Y(net6927)
);

XOR2x2_ASAP7_75t_R c6862(
.A(net6912),
.B(net3872),
.Y(net6928)
);

AO221x2_ASAP7_75t_R c6863(
.A1(net6890),
.A2(net5080),
.B1(net6925),
.B2(net6869),
.C(net6832),
.Y(net6929)
);

OA21x2_ASAP7_75t_R c6864(
.A1(net6755),
.A2(net6927),
.B(net6905),
.Y(net6930)
);

HB4xp67_ASAP7_75t_R c6865(
.A(net9241),
.Y(net6931)
);

OAI21x1_ASAP7_75t_R c6866(
.A1(net6907),
.A2(net6836),
.B(net5932),
.Y(net6932)
);

OAI21xp33_ASAP7_75t_R c6867(
.A1(net6927),
.A2(net6906),
.B(net5039),
.Y(net6933)
);

XOR2xp5_ASAP7_75t_R c6868(
.A(net6922),
.B(net10048),
.Y(net6934)
);

AND2x2_ASAP7_75t_R c6869(
.A(net6911),
.B(net6701),
.Y(net6935)
);

AND2x4_ASAP7_75t_R c6870(
.A(net4173),
.B(net6009),
.Y(net6936)
);

AND2x6_ASAP7_75t_R c6871(
.A(net6927),
.B(net9711),
.Y(net6937)
);

HAxp5_ASAP7_75t_R c6872(
.A(net6903),
.B(net6935),
.CON(net6938)
);

NAND2x1_ASAP7_75t_R c6873(
.A(net6929),
.B(net10146),
.Y(net6939)
);

NAND2x1p5_ASAP7_75t_R c6874(
.A(net6918),
.B(net6914),
.Y(net6940)
);

INVx11_ASAP7_75t_R c6875(
.A(net10036),
.Y(net6941)
);

OAI21xp5_ASAP7_75t_R c6876(
.A1(net6941),
.A2(net6749),
.B(net6737),
.Y(net6942)
);

OR3x1_ASAP7_75t_R c6877(
.A(net6018),
.B(net6942),
.C(net6881),
.Y(net6943)
);

NAND2x2_ASAP7_75t_R c6878(
.A(net6934),
.B(net6794),
.Y(net6944)
);

INVx13_ASAP7_75t_R c6879(
.A(net9970),
.Y(net6945)
);

OR3x2_ASAP7_75t_R c6880(
.A(net6902),
.B(net6940),
.C(net6945),
.Y(net6946)
);

OR3x4_ASAP7_75t_R c6881(
.A(net5983),
.B(net6942),
.C(net6928),
.Y(net6947)
);

AOI31xp67_ASAP7_75t_R c6882(
.A1(net6871),
.A2(net6937),
.A3(net6942),
.B(net6928),
.Y(net6948)
);

NAND2xp33_ASAP7_75t_R c6883(
.A(net6932),
.B(net6927),
.Y(net6949)
);

AND3x1_ASAP7_75t_R c6884(
.A(net6949),
.B(net6936),
.C(net6947),
.Y(net6950)
);

NAND4xp25_ASAP7_75t_R c6885(
.A(net6667),
.B(net6895),
.C(net6947),
.D(net6927),
.Y(net6951)
);

NAND4xp75_ASAP7_75t_R c6886(
.A(net6944),
.B(net6942),
.C(net6947),
.D(net6906),
.Y(net6952)
);

AO32x1_ASAP7_75t_R c6887(
.A1(net6951),
.A2(net6816),
.A3(net6942),
.B1(net6027),
.B2(net6914),
.Y(net6953)
);

AO32x2_ASAP7_75t_R c6888(
.A1(net6950),
.A2(net6737),
.A3(net6917),
.B1(net9760),
.B2(net10144),
.Y(net6954)
);

NAND2xp5_ASAP7_75t_R c6889(
.A(net5848),
.B(net6869),
.Y(net6955)
);

NAND2xp67_ASAP7_75t_R c6890(
.A(net4845),
.B(net5848),
.Y(net6956)
);

NOR2x1_ASAP7_75t_R c6891(
.A(net5121),
.B(net5184),
.Y(net6957)
);

NOR2x1p5_ASAP7_75t_R c6892(
.A(net2262),
.B(net10271),
.Y(net6958)
);

INVx1_ASAP7_75t_R c6893(
.A(net5747),
.Y(net6959)
);

NOR2x2_ASAP7_75t_R c6894(
.A(net6897),
.B(net6048),
.Y(net6960)
);

INVx2_ASAP7_75t_R c6895(
.A(net6102),
.Y(net6961)
);

NOR2xp33_ASAP7_75t_R c6896(
.A(net3339),
.B(net6914),
.Y(net6962)
);

NOR2xp67_ASAP7_75t_R c6897(
.A(net6864),
.B(net6815),
.Y(net6963)
);

OR2x2_ASAP7_75t_R c6898(
.A(net5978),
.B(net6016),
.Y(net6964)
);

OR2x4_ASAP7_75t_R c6899(
.A(net6962),
.B(net6895),
.Y(net6965)
);

OR2x6_ASAP7_75t_R c6900(
.A(net6109),
.B(net6102),
.Y(net6966)
);

XNOR2x1_ASAP7_75t_R c6901(
.B(net5932),
.A(net5971),
.Y(net6967)
);

XNOR2x2_ASAP7_75t_R c6902(
.A(net6956),
.B(net6101),
.Y(net6968)
);

XNOR2xp5_ASAP7_75t_R c6903(
.A(net6933),
.B(net6737),
.Y(net6969)
);

AND3x2_ASAP7_75t_R c6904(
.A(net6960),
.B(net6950),
.C(net10272),
.Y(net6970)
);

XOR2x1_ASAP7_75t_R c6905(
.A(net6926),
.B(net6968),
.Y(net6971)
);

INVx3_ASAP7_75t_R c6906(
.A(net6963),
.Y(net6972)
);

INVx4_ASAP7_75t_R c6907(
.A(net10523),
.Y(net6973)
);

XOR2x2_ASAP7_75t_R c6908(
.A(net6815),
.B(net6960),
.Y(net6974)
);

XOR2xp5_ASAP7_75t_R c6909(
.A(net6737),
.B(net6972),
.Y(net6975)
);

INVx5_ASAP7_75t_R c6910(
.A(net10346),
.Y(net6976)
);

AND2x2_ASAP7_75t_R c6911(
.A(net6968),
.B(net6919),
.Y(net6977)
);

INVx6_ASAP7_75t_R c6912(
.A(net10128),
.Y(net6978)
);

AND2x4_ASAP7_75t_R c6913(
.A(net6758),
.B(net10081),
.Y(net6979)
);

AND2x6_ASAP7_75t_R c6914(
.A(net5184),
.B(net5926),
.Y(net6980)
);

HAxp5_ASAP7_75t_R c6915(
.A(net6048),
.B(net6109),
.CON(net6981)
);

AND3x4_ASAP7_75t_R c6916(
.A(net6855),
.B(net6968),
.C(net10272),
.Y(net6982)
);

INVx8_ASAP7_75t_R c6917(
.A(net10416),
.Y(net6983)
);

NAND2x1_ASAP7_75t_R c6918(
.A(net6791),
.B(net6102),
.Y(net6984)
);

NAND2x1p5_ASAP7_75t_R c6919(
.A(net6959),
.B(net6027),
.Y(net6985)
);

NAND2x2_ASAP7_75t_R c6920(
.A(net6045),
.B(net6968),
.Y(net6986)
);

INVxp33_ASAP7_75t_R c6921(
.A(net10366),
.Y(net6987)
);

NAND2xp33_ASAP7_75t_R c6922(
.A(net6978),
.B(net9678),
.Y(net6988)
);

NAND2xp5_ASAP7_75t_R c6923(
.A(net6493),
.B(net6978),
.Y(net6989)
);

INVxp67_ASAP7_75t_R c6924(
.A(net10488),
.Y(net6990)
);

NAND2xp67_ASAP7_75t_R c6925(
.A(net6519),
.B(net6974),
.Y(net6991)
);

NOR4xp25_ASAP7_75t_R c6926(
.A(net6977),
.B(net6987),
.C(net6031),
.D(net6016),
.Y(net6992)
);

NOR2x1_ASAP7_75t_R c6927(
.A(net6981),
.B(net6104),
.Y(net6993)
);

NOR2x1p5_ASAP7_75t_R c6928(
.A(net6990),
.B(net6102),
.Y(net6994)
);

AO21x1_ASAP7_75t_R c6929(
.A1(net6087),
.A2(net6967),
.B(net6988),
.Y(net6995)
);

NOR2x2_ASAP7_75t_R c6930(
.A(net6965),
.B(net6948),
.Y(net6996)
);

NOR2xp33_ASAP7_75t_R c6931(
.A(net6057),
.B(net6987),
.Y(net6997)
);

NOR2xp67_ASAP7_75t_R c6932(
.A(net6104),
.B(net6905),
.Y(net6998)
);

OR2x2_ASAP7_75t_R c6933(
.A(net6983),
.B(net6987),
.Y(net6999)
);

BUFx10_ASAP7_75t_R c6934(
.A(net10370),
.Y(net7000)
);

OR2x4_ASAP7_75t_R c6935(
.A(net6974),
.B(net7000),
.Y(net7001)
);

BUFx12_ASAP7_75t_R c6936(
.A(net10156),
.Y(net7002)
);

OR2x6_ASAP7_75t_R c6937(
.A(net6998),
.B(net6887),
.Y(net7003)
);

XNOR2x1_ASAP7_75t_R c6938(
.B(net6919),
.A(net6928),
.Y(net7004)
);

BUFx12f_ASAP7_75t_R c6939(
.A(net10551),
.Y(net7005)
);

OA33x2_ASAP7_75t_R c6940(
.A1(net6999),
.A2(net7005),
.A3(net6069),
.B1(net5932),
.B2(net6972),
.B3(net5726),
.Y(net7006)
);

XNOR2x2_ASAP7_75t_R c6941(
.A(net7002),
.B(net6904),
.Y(net7007)
);

BUFx16f_ASAP7_75t_R c6942(
.A(net10384),
.Y(net7008)
);

AO21x2_ASAP7_75t_R c6943(
.A1(net6991),
.A2(net10149),
.B(net10284),
.Y(net7009)
);

XNOR2xp5_ASAP7_75t_R c6944(
.A(net7009),
.B(net7005),
.Y(net7010)
);

XOR2x1_ASAP7_75t_R c6945(
.A(net7004),
.B(net10081),
.Y(net7011)
);

XOR2x2_ASAP7_75t_R c6946(
.A(net5181),
.B(net6968),
.Y(net7012)
);

XOR2xp5_ASAP7_75t_R c6947(
.A(net6904),
.B(net6960),
.Y(net7013)
);

BUFx24_ASAP7_75t_R c6948(
.A(net9973),
.Y(net7014)
);

AND2x2_ASAP7_75t_R c6949(
.A(net6989),
.B(net6967),
.Y(net7015)
);

AND2x4_ASAP7_75t_R c6950(
.A(net7011),
.B(net5848),
.Y(net7016)
);

AOI21x1_ASAP7_75t_R c6951(
.A1(net7001),
.A2(net7004),
.B(net7016),
.Y(net7017)
);

SDFHx4_ASAP7_75t_R c6952(
.D(net5163),
.SE(net7015),
.SI(net6898),
.CLK(clk),
.QN(net7018)
);

BUFx2_ASAP7_75t_R c6953(
.A(net10346),
.Y(net7019)
);

NOR4xp75_ASAP7_75t_R c6954(
.A(net6978),
.B(net5968),
.C(net6104),
.D(net6979),
.Y(net7020)
);

AOI221x1_ASAP7_75t_R c6955(
.A1(net6999),
.A2(net7015),
.B1(net6972),
.B2(net7019),
.C(net10149),
.Y(net7021)
);

AND2x6_ASAP7_75t_R c6956(
.A(net6995),
.B(net7018),
.Y(net7022)
);

HAxp5_ASAP7_75t_R c6957(
.A(net6987),
.B(net7017),
.CON(net7023)
);

AOI21xp33_ASAP7_75t_R c6958(
.A1(net6920),
.A2(net6026),
.B(net7021),
.Y(net7024)
);

SDFLx1_ASAP7_75t_R c6959(
.D(net6980),
.SE(net6979),
.SI(net7009),
.CLK(clk),
.QN(net7025)
);

SDFLx2_ASAP7_75t_R c6960(
.D(net7021),
.SE(net7025),
.SI(net5076),
.CLK(clk),
.QN(net7026)
);

OAI222xp33_ASAP7_75t_R c6961(
.A1(net7022),
.A2(net7013),
.B1(net7021),
.B2(net5076),
.C1(net7026),
.C2(net6791),
.Y(net7027)
);

AOI21xp5_ASAP7_75t_R c6962(
.A1(net7016),
.A2(net10167),
.B(net10254),
.Y(net7028)
);

FAx1_ASAP7_75t_R c6963(
.A(net5130),
.B(net7000),
.CI(net10167),
.SN(net7029)
);

MAJIxp5_ASAP7_75t_R c6964(
.A(net7029),
.B(net7014),
.C(net7020),
.Y(net7030)
);

MAJx2_ASAP7_75t_R c6965(
.A(net7018),
.B(net7021),
.C(net6917),
.Y(net7031)
);

MAJx3_ASAP7_75t_R c6966(
.A(net6996),
.B(net6950),
.C(net7019),
.Y(net7032)
);

NAND3x1_ASAP7_75t_R c6967(
.A(net6991),
.B(net6976),
.C(net10167),
.Y(net7033)
);

NAND3x2_ASAP7_75t_R c6968(
.B(net7020),
.C(net7025),
.A(net7033),
.Y(net7034)
);

O2A1O1Ixp33_ASAP7_75t_R c6969(
.A1(net6971),
.A2(net7016),
.B(net6972),
.C(net9972),
.Y(net7035)
);

OAI321xp33_ASAP7_75t_R c6970(
.A1(net4185),
.A2(net7025),
.A3(net4953),
.B1(net6960),
.B2(net7026),
.C(net10284),
.Y(net7036)
);

O2A1O1Ixp5_ASAP7_75t_R c6971(
.A1(net7000),
.A2(net7006),
.B(net5115),
.C(net6058),
.Y(net7037)
);

SDFLx3_ASAP7_75t_R c6972(
.D(net4349),
.SE(net6027),
.SI(net6643),
.CLK(clk),
.QN(net7038)
);

NAND3xp33_ASAP7_75t_R c6973(
.A(net6993),
.B(net3404),
.C(net6808),
.Y(net7039)
);

NAND2x1_ASAP7_75t_R c6974(
.A(net6128),
.B(net10254),
.Y(net7040)
);

BUFx3_ASAP7_75t_R c6975(
.A(net6178),
.Y(net7041)
);

BUFx4_ASAP7_75t_R c6976(
.A(net6878),
.Y(net7042)
);

BUFx4f_ASAP7_75t_R c6977(
.A(net9122),
.Y(net7043)
);

BUFx5_ASAP7_75t_R c6978(
.A(net9122),
.Y(net7044)
);

BUFx6f_ASAP7_75t_R c6979(
.A(net10467),
.Y(net7045)
);

NAND2x1p5_ASAP7_75t_R c6980(
.A(net3366),
.B(net6887),
.Y(net7046)
);

BUFx8_ASAP7_75t_R c6981(
.A(net6758),
.Y(net7047)
);

NAND2x2_ASAP7_75t_R c6982(
.A(net6898),
.B(net10135),
.Y(net7048)
);

CKINVDCx10_ASAP7_75t_R c6983(
.A(net10135),
.Y(net7049)
);

SDFLx4_ASAP7_75t_R c6984(
.D(net5926),
.SE(net6863),
.SI(net6198),
.CLK(clk),
.QN(net7050)
);

CKINVDCx11_ASAP7_75t_R c6985(
.A(net10368),
.Y(net7051)
);

CKINVDCx12_ASAP7_75t_R c6986(
.A(net10382),
.Y(net7052)
);

DFFASRHQNx1_ASAP7_75t_R c6987(
.D(net6863),
.RESETN(net6136),
.SETN(net5726),
.CLK(clk),
.QN(net7053)
);

CKINVDCx14_ASAP7_75t_R c6988(
.A(net10493),
.Y(net7054)
);

CKINVDCx16_ASAP7_75t_R c6989(
.A(net10094),
.Y(net7055)
);

NAND2xp33_ASAP7_75t_R c6990(
.A(net6040),
.B(net7045),
.Y(net7056)
);

NAND2xp5_ASAP7_75t_R c6991(
.A(net6140),
.B(net7053),
.Y(net7057)
);

CKINVDCx20_ASAP7_75t_R c6992(
.A(net6931),
.Y(net7058)
);

CKINVDCx5p33_ASAP7_75t_R c6993(
.A(net10148),
.Y(net7059)
);

CKINVDCx6p67_ASAP7_75t_R c6994(
.A(net6158),
.Y(net7060)
);

NAND2xp67_ASAP7_75t_R c6995(
.A(net7003),
.B(net5971),
.Y(net7061)
);

NOR2x1_ASAP7_75t_R c6996(
.A(net6072),
.B(net7044),
.Y(net7062)
);

CKINVDCx8_ASAP7_75t_R c6997(
.A(net7007),
.Y(net7063)
);

NOR2x1p5_ASAP7_75t_R c6998(
.A(net7062),
.B(net5266),
.Y(net7064)
);

NOR2x2_ASAP7_75t_R c6999(
.A(net5110),
.B(net7056),
.Y(net7065)
);

NOR2xp33_ASAP7_75t_R c7000(
.A(net7049),
.B(net6154),
.Y(net7066)
);

NOR3x1_ASAP7_75t_R c7001(
.A(net6193),
.B(net7066),
.C(net6837),
.Y(net7067)
);

NOR2xp67_ASAP7_75t_R c7002(
.A(net6901),
.B(net7044),
.Y(net7068)
);

OR2x2_ASAP7_75t_R c7003(
.A(net7065),
.B(net6178),
.Y(net7069)
);

OR2x4_ASAP7_75t_R c7004(
.A(net6071),
.B(net7061),
.Y(net7070)
);

CKINVDCx9p33_ASAP7_75t_R c7005(
.A(net9204),
.Y(net7071)
);

HB1xp67_ASAP7_75t_R c7006(
.A(net10423),
.Y(net7072)
);

OR2x6_ASAP7_75t_R c7007(
.A(net6181),
.B(net7052),
.Y(net7073)
);

XNOR2x1_ASAP7_75t_R c7008(
.B(net7070),
.A(net7053),
.Y(net7074)
);

NOR3x2_ASAP7_75t_R c7009(
.B(net7071),
.C(net6991),
.A(net7073),
.Y(net7075)
);

HB2xp67_ASAP7_75t_R c7010(
.A(net6097),
.Y(net7076)
);

XNOR2x2_ASAP7_75t_R c7011(
.A(net6808),
.B(net6931),
.Y(net7077)
);

XNOR2xp5_ASAP7_75t_R c7012(
.A(net6969),
.B(net7054),
.Y(net7078)
);

XOR2x1_ASAP7_75t_R c7013(
.A(net7072),
.B(net6146),
.Y(net7079)
);

ICGx4DC_ASAP7_75t_R c7014(
.ENA(net6929),
.SE(net6979),
.CLK(clk),
.GCLK(net7080)
);

XOR2x2_ASAP7_75t_R c7015(
.A(net6976),
.B(net7050),
.Y(net7081)
);

NOR3xp33_ASAP7_75t_R c7016(
.A(net7081),
.B(net7067),
.C(net5110),
.Y(net7082)
);

OA21x2_ASAP7_75t_R c7017(
.A1(net7055),
.A2(net7082),
.B(net7057),
.Y(net7083)
);

HB3xp67_ASAP7_75t_R c7018(
.A(net10375),
.Y(net7084)
);

XOR2xp5_ASAP7_75t_R c7019(
.A(net1490),
.B(net5964),
.Y(net7085)
);

OAI21x1_ASAP7_75t_R c7020(
.A1(net7080),
.A2(net7071),
.B(net5110),
.Y(net7086)
);

AND2x2_ASAP7_75t_R c7021(
.A(net7077),
.B(net6166),
.Y(net7087)
);

HB4xp67_ASAP7_75t_R c7022(
.A(net10368),
.Y(net7088)
);

AND2x4_ASAP7_75t_R c7023(
.A(net7078),
.B(net6136),
.Y(net7089)
);

ICGx4_ASAP7_75t_R c7024(
.ENA(net6961),
.SE(net7080),
.CLK(clk),
.GCLK(net7090)
);

OAI21xp33_ASAP7_75t_R c7025(
.A1(net6174),
.A2(net7085),
.B(net7087),
.Y(net7091)
);

AND2x6_ASAP7_75t_R c7026(
.A(net6097),
.B(net10142),
.Y(net7092)
);

HAxp5_ASAP7_75t_R c7027(
.A(net4099),
.B(net10254),
.CON(net7094),
.SN(net7093)
);

NAND2x1_ASAP7_75t_R c7028(
.A(net4310),
.B(net7083),
.Y(net7095)
);

SDFHx1_ASAP7_75t_R c7029(
.D(net7092),
.SE(net7053),
.SI(net7060),
.CLK(clk),
.QN(net7096)
);

INVx11_ASAP7_75t_R c7030(
.A(net10003),
.Y(net7097)
);

NAND2x1p5_ASAP7_75t_R c7031(
.A(net7097),
.B(net7054),
.Y(net7098)
);

INVx13_ASAP7_75t_R c7032(
.A(net7044),
.Y(net7099)
);

OAI33xp33_ASAP7_75t_R c7033(
.A1(net7082),
.A2(net6859),
.A3(net6097),
.B1(net6979),
.B2(net7026),
.B3(net7054),
.Y(net7100)
);

NAND2x2_ASAP7_75t_R c7034(
.A(net7098),
.B(net7087),
.Y(net7101)
);

NAND2xp33_ASAP7_75t_R c7035(
.A(net6153),
.B(net7082),
.Y(net7102)
);

OAI21xp5_ASAP7_75t_R c7036(
.A1(net7079),
.A2(net7050),
.B(net10135),
.Y(net7103)
);

NAND2xp5_ASAP7_75t_R c7037(
.A(net7086),
.B(net6072),
.Y(net7104)
);

OR3x1_ASAP7_75t_R c7038(
.A(net2474),
.B(net6146),
.C(net7050),
.Y(net7105)
);

NAND2xp67_ASAP7_75t_R c7039(
.A(net7104),
.B(net6154),
.Y(net7106)
);

NOR2x1_ASAP7_75t_R c7040(
.A(net7088),
.B(net6863),
.Y(net7107)
);

OR3x2_ASAP7_75t_R c7041(
.A(net7004),
.B(net5110),
.C(net6140),
.Y(net7108)
);

NOR2x1p5_ASAP7_75t_R c7042(
.A(net7094),
.B(net7103),
.Y(net7109)
);

NOR2x2_ASAP7_75t_R c7043(
.A(net7107),
.B(net7106),
.Y(net7110)
);

NOR2xp33_ASAP7_75t_R c7044(
.A(net6859),
.B(net5255),
.Y(net7111)
);

OR3x4_ASAP7_75t_R c7045(
.A(net3267),
.B(net6972),
.C(net7066),
.Y(net7112)
);

NOR2xp67_ASAP7_75t_R c7046(
.A(net7099),
.B(net7104),
.Y(net7113)
);

INVx1_ASAP7_75t_R c7047(
.A(net10452),
.Y(net7114)
);

OR2x2_ASAP7_75t_R c7048(
.A(net7103),
.B(net7093),
.Y(net7115)
);

INVx2_ASAP7_75t_R c7049(
.A(net10442),
.Y(net7116)
);

INVx3_ASAP7_75t_R c7050(
.A(net10142),
.Y(net7117)
);

SDFHx2_ASAP7_75t_R c7051(
.D(net7109),
.SE(net7095),
.SI(net7085),
.CLK(clk),
.QN(net7118)
);

SDFHx3_ASAP7_75t_R c7052(
.D(net3404),
.SE(net6859),
.SI(net7060),
.CLK(clk),
.QN(net7119)
);

AND3x1_ASAP7_75t_R c7053(
.A(net7117),
.B(net7114),
.C(net7119),
.Y(net7120)
);

AND3x2_ASAP7_75t_R c7054(
.A(net7120),
.B(net7092),
.C(net7118),
.Y(net7121)
);

INVx4_ASAP7_75t_R c7055(
.A(net10398),
.Y(net7122)
);

OR2x4_ASAP7_75t_R c7056(
.A(net2459),
.B(net5325),
.Y(net7123)
);

OR2x6_ASAP7_75t_R c7057(
.A(net4419),
.B(net10284),
.Y(net7124)
);

INVx5_ASAP7_75t_R c7058(
.A(net10331),
.Y(net7125)
);

XNOR2x1_ASAP7_75t_R c7059(
.B(net3460),
.A(net6129),
.Y(net7126)
);

INVx6_ASAP7_75t_R c7060(
.A(net10374),
.Y(net7127)
);

INVx8_ASAP7_75t_R c7061(
.A(net10396),
.Y(net7128)
);

OA211x2_ASAP7_75t_R c7062(
.A1(net7123),
.A2(net7083),
.B(net6816),
.C(net5260),
.Y(net7129)
);

XNOR2x2_ASAP7_75t_R c7063(
.A(net6247),
.B(net6272),
.Y(net7130)
);

SDFHx4_ASAP7_75t_R c7064(
.D(net5336),
.SE(net6247),
.SI(net7043),
.CLK(clk),
.QN(net7131)
);

XNOR2xp5_ASAP7_75t_R c7065(
.A(net6265),
.B(net10284),
.Y(net7132)
);

XOR2x1_ASAP7_75t_R c7066(
.A(net7110),
.B(net5349),
.Y(net7133)
);

XOR2x2_ASAP7_75t_R c7067(
.A(net7087),
.B(net7038),
.Y(net7134)
);

SDFLx1_ASAP7_75t_R c7068(
.D(net4377),
.SE(net7124),
.SI(net6204),
.CLK(clk),
.QN(net7135)
);

INVxp33_ASAP7_75t_R c7069(
.A(net10394),
.Y(net7136)
);

INVxp67_ASAP7_75t_R c7070(
.A(out0),
.Y(net7137)
);

XOR2xp5_ASAP7_75t_R c7071(
.A(net7135),
.B(net10198),
.Y(net7138)
);

AND2x2_ASAP7_75t_R c7072(
.A(net4419),
.B(net6058),
.Y(net7139)
);

BUFx10_ASAP7_75t_R c7073(
.A(net10118),
.Y(net7140)
);

AND2x4_ASAP7_75t_R c7074(
.A(net6246),
.B(net7069),
.Y(net7141)
);

AND2x6_ASAP7_75t_R c7075(
.A(net7073),
.B(net6885),
.Y(net7142)
);

AOI221xp5_ASAP7_75t_R c7076(
.A1(net6249),
.A2(net4310),
.B1(net6183),
.B2(net5883),
.C(net3443),
.Y(net7143)
);

OA22x2_ASAP7_75t_R c7077(
.A1(net7137),
.A2(net6214),
.B1(net5336),
.B2(net7138),
.Y(net7144)
);

HAxp5_ASAP7_75t_R c7078(
.A(net7059),
.B(net7064),
.CON(net7146),
.SN(net7145)
);

AND3x4_ASAP7_75t_R c7079(
.A(net7127),
.B(net7131),
.C(net7064),
.Y(net7147)
);

BUFx12_ASAP7_75t_R c7080(
.A(net10375),
.Y(net7148)
);

NAND2x1_ASAP7_75t_R c7081(
.A(net609),
.B(net7073),
.Y(net7149)
);

NAND2x1p5_ASAP7_75t_R c7082(
.A(net6222),
.B(net10284),
.Y(net7150)
);

NAND2x2_ASAP7_75t_R c7083(
.A(net5237),
.B(net7079),
.Y(net7151)
);

NAND2xp33_ASAP7_75t_R c7084(
.A(net7016),
.B(net6885),
.Y(net7152)
);

BUFx12f_ASAP7_75t_R c7085(
.A(net10447),
.Y(net7153)
);

NAND2xp5_ASAP7_75t_R c7086(
.A(net6885),
.B(net7016),
.Y(net7154)
);

AO21x1_ASAP7_75t_R c7087(
.A1(net5349),
.A2(net6204),
.B(net7136),
.Y(net7155)
);

OA31x2_ASAP7_75t_R c7088(
.A1(net6243),
.A2(net1653),
.A3(net7138),
.B1(net10286),
.Y(net7156)
);

BUFx16f_ASAP7_75t_R c7089(
.A(net10570),
.Y(net7157)
);

AO222x2_ASAP7_75t_R c7090(
.A1(net5267),
.A2(net6222),
.B1(net6267),
.B2(net7148),
.C1(net6265),
.C2(net10287),
.Y(net7158)
);

AO21x2_ASAP7_75t_R c7091(
.A1(net7133),
.A2(net5237),
.B(net7127),
.Y(net7159)
);

NAND2xp67_ASAP7_75t_R c7092(
.A(net7154),
.B(net7026),
.Y(net7160)
);

NOR2x1_ASAP7_75t_R c7093(
.A(net7079),
.B(net7123),
.Y(net7161)
);

NOR2x1p5_ASAP7_75t_R c7094(
.A(net6252),
.B(net10287),
.Y(net7162)
);

BUFx24_ASAP7_75t_R c7095(
.A(net10558),
.Y(net7163)
);

NOR2x2_ASAP7_75t_R c7096(
.A(net7155),
.B(net7108),
.Y(net7164)
);

NOR2xp33_ASAP7_75t_R c7097(
.A(net7063),
.B(net6267),
.Y(net7165)
);

BUFx2_ASAP7_75t_R c7098(
.A(net10447),
.Y(net7166)
);

NOR2xp67_ASAP7_75t_R c7099(
.A(net7140),
.B(net7155),
.Y(net7167)
);

BUFx3_ASAP7_75t_R c7100(
.A(net10119),
.Y(net7168)
);

SDFLx2_ASAP7_75t_R c7101(
.D(net6283),
.SE(net7152),
.SI(net7162),
.CLK(clk),
.QN(net7169)
);

OR2x2_ASAP7_75t_R c7102(
.A(net5266),
.B(net7152),
.Y(net7170)
);

OR2x4_ASAP7_75t_R c7103(
.A(net7150),
.B(net7161),
.Y(net7171)
);

OR2x6_ASAP7_75t_R c7104(
.A(net7166),
.B(net7170),
.Y(net7172)
);

XNOR2x1_ASAP7_75t_R c7105(
.B(net7132),
.A(net7171),
.Y(net7173)
);

XNOR2x2_ASAP7_75t_R c7106(
.A(net6267),
.B(net7111),
.Y(net7174)
);

XNOR2xp5_ASAP7_75t_R c7107(
.A(net7173),
.B(net7172),
.Y(net7175)
);

AOI21x1_ASAP7_75t_R c7108(
.A1(net7169),
.A2(net6209),
.B(net9902),
.Y(net7176)
);

XOR2x1_ASAP7_75t_R c7109(
.A(net7152),
.B(net7167),
.Y(net7177)
);

XOR2x2_ASAP7_75t_R c7110(
.A(net6203),
.B(net7168),
.Y(net7178)
);

XOR2xp5_ASAP7_75t_R c7111(
.A(net7174),
.B(net9671),
.Y(net7179)
);

AND2x2_ASAP7_75t_R c7112(
.A(net7167),
.B(net7054),
.Y(net7180)
);

AND2x4_ASAP7_75t_R c7113(
.A(net7171),
.B(net7169),
.Y(net7181)
);

AND2x6_ASAP7_75t_R c7114(
.A(net7176),
.B(net6267),
.Y(net7182)
);

HAxp5_ASAP7_75t_R c7115(
.A(net7084),
.B(net7147),
.CON(net7184),
.SN(net7183)
);

OAI211xp5_ASAP7_75t_R c7116(
.A1(net7131),
.A2(net7178),
.B(net4369),
.C(net7026),
.Y(net7185)
);

AOI21xp33_ASAP7_75t_R c7117(
.A1(net7066),
.A2(net6146),
.B(net7161),
.Y(net7186)
);

NAND2x1_ASAP7_75t_R c7118(
.A(net677),
.B(net7033),
.Y(net7187)
);

NAND2x1p5_ASAP7_75t_R c7119(
.A(net7149),
.B(net7168),
.Y(net7188)
);

AOI21xp5_ASAP7_75t_R c7120(
.A1(net7187),
.A2(net7155),
.B(net7182),
.Y(net7189)
);

SDFLx3_ASAP7_75t_R c7121(
.D(net4302),
.SE(net7152),
.SI(net7189),
.CLK(clk),
.QN(net7190)
);

FAx1_ASAP7_75t_R c7122(
.A(net7177),
.B(out25),
.CI(net7176),
.SN(net7191)
);

NAND2x2_ASAP7_75t_R c7123(
.A(net6991),
.B(net4363),
.Y(net7192)
);

MAJIxp5_ASAP7_75t_R c7124(
.A(net7186),
.B(net7190),
.C(net7183),
.Y(net7193)
);

NAND2xp33_ASAP7_75t_R c7125(
.A(net7180),
.B(net7168),
.Y(net7194)
);

MAJx2_ASAP7_75t_R c7126(
.A(net7010),
.B(net7181),
.C(net7187),
.Y(net7195)
);

NAND2xp5_ASAP7_75t_R c7127(
.A(net7194),
.B(net7193),
.Y(net7196)
);

MAJx3_ASAP7_75t_R c7128(
.A(net6891),
.B(net7196),
.C(net7187),
.Y(net7197)
);

NAND3x1_ASAP7_75t_R c7129(
.A(net7182),
.B(net7173),
.C(net7187),
.Y(net7198)
);

NAND3x2_ASAP7_75t_R c7130(
.B(net7042),
.C(net7123),
.A(net7113),
.Y(net7199)
);

SDFLx4_ASAP7_75t_R c7131(
.D(net7195),
.SE(net7176),
.SI(net6191),
.CLK(clk),
.QN(net7200)
);

NAND3xp33_ASAP7_75t_R c7132(
.A(net7188),
.B(net7133),
.C(net7199),
.Y(net7201)
);

OAI22x1_ASAP7_75t_R c7133(
.A1(net7128),
.A2(net7138),
.B1(net5236),
.B2(net10242),
.Y(net7202)
);

DFFASRHQNx1_ASAP7_75t_R c7134(
.D(net7199),
.RESETN(net7194),
.SETN(net7200),
.CLK(clk),
.QN(net7203)
);

AO33x2_ASAP7_75t_R c7135(
.A1(net7174),
.A2(net7200),
.A3(net7176),
.B1(net6267),
.B2(net7178),
.B3(net7179),
.Y(net7204)
);

NOR3x1_ASAP7_75t_R c7136(
.A(net9914),
.B(net10114),
.C(net10288),
.Y(net7205)
);

BUFx4_ASAP7_75t_R c7137(
.A(net10331),
.Y(net7206)
);

NAND2xp67_ASAP7_75t_R c7138(
.A(net6957),
.B(net6347),
.Y(net7207)
);

NOR2x1_ASAP7_75t_R c7139(
.A(net7130),
.B(net6225),
.Y(net7208)
);

NOR2x1p5_ASAP7_75t_R c7140(
.A(net6305),
.B(net6887),
.Y(net7209)
);

NOR2x2_ASAP7_75t_R c7141(
.A(net7203),
.B(net3564),
.Y(net7210)
);

NOR2xp33_ASAP7_75t_R c7142(
.A(net2642),
.B(net7185),
.Y(net7211)
);

NOR2xp67_ASAP7_75t_R c7143(
.A(net7125),
.B(net6362),
.Y(net7212)
);

BUFx4f_ASAP7_75t_R c7144(
.A(net10353),
.Y(net7213)
);

OR2x2_ASAP7_75t_R c7145(
.A(net4099),
.B(net6347),
.Y(net7214)
);

OR2x4_ASAP7_75t_R c7146(
.A(net6341),
.B(net6323),
.Y(net7215)
);

BUFx5_ASAP7_75t_R c7147(
.A(net10332),
.Y(net7216)
);

OR2x6_ASAP7_75t_R c7148(
.A(net6225),
.B(net7148),
.Y(net7217)
);

XNOR2x1_ASAP7_75t_R c7149(
.B(net7141),
.A(net7192),
.Y(net7218)
);

XNOR2x2_ASAP7_75t_R c7150(
.A(net6349),
.B(net7214),
.Y(net7219)
);

XNOR2xp5_ASAP7_75t_R c7151(
.A(net7185),
.B(net7203),
.Y(net7220)
);

XOR2x1_ASAP7_75t_R c7152(
.A(net7209),
.B(net7213),
.Y(net7221)
);

NOR3x2_ASAP7_75t_R c7153(
.B(net4492),
.C(net5726),
.A(net10288),
.Y(net7222)
);

NOR3xp33_ASAP7_75t_R c7154(
.A(net7214),
.B(net7057),
.C(net3557),
.Y(net7223)
);

XOR2x2_ASAP7_75t_R c7155(
.A(net7113),
.B(net4502),
.Y(net7224)
);

AOI311xp33_ASAP7_75t_R c7156(
.A1(net2617),
.A2(net5409),
.A3(net2578),
.B(net6342),
.C(net10228),
.Y(net7225)
);

XOR2xp5_ASAP7_75t_R c7157(
.A(net6310),
.B(net6204),
.Y(net7226)
);

AND2x2_ASAP7_75t_R c7158(
.A(net5398),
.B(net686),
.Y(net7227)
);

AND2x4_ASAP7_75t_R c7159(
.A(net4502),
.B(net7214),
.Y(net7228)
);

AND2x6_ASAP7_75t_R c7160(
.A(net6351),
.B(net6225),
.Y(net7229)
);

BUFx6f_ASAP7_75t_R c7161(
.A(net10332),
.Y(net7230)
);

HAxp5_ASAP7_75t_R c7162(
.A(net4469),
.B(net10242),
.CON(net7231)
);

NAND2x1_ASAP7_75t_R c7163(
.A(net6316),
.B(net7208),
.Y(net7232)
);

NAND2x1p5_ASAP7_75t_R c7164(
.A(net7213),
.B(net7217),
.Y(net7233)
);

NAND2x2_ASAP7_75t_R c7165(
.A(net7219),
.B(net7214),
.Y(net7234)
);

NAND2xp33_ASAP7_75t_R c7166(
.A(net7038),
.B(net7208),
.Y(net7235)
);

NAND2xp5_ASAP7_75t_R c7167(
.A(net7135),
.B(net5398),
.Y(net7236)
);

BUFx8_ASAP7_75t_R c7168(
.A(net10382),
.Y(net7237)
);

NAND2xp67_ASAP7_75t_R c7169(
.A(net7208),
.B(net3557),
.Y(net7238)
);

OA21x2_ASAP7_75t_R c7170(
.A1(net7170),
.A2(net7125),
.B(net10288),
.Y(net7239)
);

NOR2x1_ASAP7_75t_R c7171(
.A(net7234),
.B(net7141),
.Y(net7240)
);

OAI21x1_ASAP7_75t_R c7172(
.A1(net5402),
.A2(net4492),
.B(net7207),
.Y(net7241)
);

OAI21xp33_ASAP7_75t_R c7173(
.A1(net7102),
.A2(net7220),
.B(net7208),
.Y(net7242)
);

OAI21xp5_ASAP7_75t_R c7174(
.A1(net7220),
.A2(net7113),
.B(net7096),
.Y(net7243)
);

NOR2x1p5_ASAP7_75t_R c7175(
.A(net7235),
.B(net6342),
.Y(net7244)
);

OR3x1_ASAP7_75t_R c7176(
.A(net7231),
.B(net7220),
.C(net5414),
.Y(net7245)
);

NOR2x2_ASAP7_75t_R c7177(
.A(net7211),
.B(net7178),
.Y(net7246)
);

SDFHx1_ASAP7_75t_R c7178(
.D(net7221),
.SE(net7239),
.SI(net5443),
.CLK(clk),
.QN(net7247)
);

SDFHx2_ASAP7_75t_R c7179(
.D(net6361),
.SE(net6310),
.SI(net6342),
.CLK(clk),
.QN(net7248)
);

NOR2xp33_ASAP7_75t_R c7180(
.A(net7238),
.B(net9720),
.Y(net7249)
);

OR3x2_ASAP7_75t_R c7181(
.A(net7096),
.B(net5354),
.C(net6213),
.Y(net7250)
);

SDFHx3_ASAP7_75t_R c7182(
.D(net6226),
.SE(net7235),
.SI(net5385),
.CLK(clk),
.QN(net7251)
);

OR3x4_ASAP7_75t_R c7183(
.A(net7250),
.B(net7247),
.C(net10122),
.Y(net7252)
);

CKINVDCx10_ASAP7_75t_R c7184(
.A(net10500),
.Y(net7253)
);

AND3x1_ASAP7_75t_R c7185(
.A(net7218),
.B(net7161),
.C(net6224),
.Y(net7254)
);

NOR2xp67_ASAP7_75t_R c7186(
.A(net7228),
.B(net7215),
.Y(net7255)
);

AND3x2_ASAP7_75t_R c7187(
.A(net6289),
.B(net7251),
.C(net7239),
.Y(net7256)
);

AND3x4_ASAP7_75t_R c7188(
.A(net6288),
.B(net7251),
.C(net7229),
.Y(net7257)
);

OR2x2_ASAP7_75t_R c7189(
.A(net4484),
.B(net7247),
.Y(net7258)
);

AO21x1_ASAP7_75t_R c7190(
.A1(net7238),
.A2(net7258),
.B(net5377),
.Y(net7259)
);

OR2x4_ASAP7_75t_R c7191(
.A(net7142),
.B(net7210),
.Y(net7260)
);

AO21x2_ASAP7_75t_R c7192(
.A1(net7251),
.A2(net6293),
.B(net7248),
.Y(net7261)
);

OR2x6_ASAP7_75t_R c7193(
.A(net7261),
.B(net7223),
.Y(net7262)
);

XNOR2x1_ASAP7_75t_R c7194(
.B(net7249),
.A(net7230),
.Y(net7263)
);

AOI32xp33_ASAP7_75t_R c7195(
.A1(net7222),
.A2(net7207),
.A3(net7179),
.B1(net4502),
.B2(net7232),
.Y(net7264)
);

SDFHx4_ASAP7_75t_R c7196(
.D(net5296),
.SE(net7258),
.SI(net7179),
.CLK(clk),
.QN(net7265)
);

XNOR2x2_ASAP7_75t_R c7197(
.A(net7253),
.B(net7255),
.Y(net7266)
);

AOI21x1_ASAP7_75t_R c7198(
.A1(net7266),
.A2(net7178),
.B(net9831),
.Y(net7267)
);

AOI21xp33_ASAP7_75t_R c7199(
.A1(net7229),
.A2(net7215),
.B(net6335),
.Y(net7268)
);

XNOR2xp5_ASAP7_75t_R c7200(
.A(net7243),
.B(net7262),
.Y(net7269)
);

XOR2x1_ASAP7_75t_R c7201(
.A(net7246),
.B(net7265),
.Y(net7270)
);

CKINVDCx11_ASAP7_75t_R c7202(
.A(net10371),
.Y(net7271)
);

XOR2x2_ASAP7_75t_R c7203(
.A(net7266),
.B(net7265),
.Y(net7272)
);

AOI21xp5_ASAP7_75t_R c7204(
.A1(net7262),
.A2(net6332),
.B(net9720),
.Y(net7273)
);

FAx1_ASAP7_75t_R c7205(
.A(net5397),
.B(net7272),
.CI(net7179),
.SN(net7274)
);

AOI222xp33_ASAP7_75t_R c7206(
.A1(net7157),
.A2(net6362),
.B1(net7268),
.B2(net7251),
.C1(net7161),
.C2(net7265),
.Y(net7275)
);

MAJIxp5_ASAP7_75t_R c7207(
.A(net6272),
.B(net7232),
.C(net9847),
.Y(net7276)
);

CKINVDCx12_ASAP7_75t_R c7208(
.A(net10042),
.Y(net7277)
);

MAJx2_ASAP7_75t_R c7209(
.A(net7236),
.B(net7179),
.C(net7240),
.Y(net7278)
);

OAI22xp33_ASAP7_75t_R c7210(
.A1(net7275),
.A2(net7214),
.B1(net7268),
.B2(net10041),
.Y(net7279)
);

NAND5xp2_ASAP7_75t_R c7211(
.A(net2661),
.B(net7229),
.C(net7268),
.D(net5267),
.E(net10030),
.Y(net7280)
);

XOR2xp5_ASAP7_75t_R c7212(
.A(net5284),
.B(net4484),
.Y(net7281)
);

MAJx3_ASAP7_75t_R c7213(
.A(net5354),
.B(net7248),
.C(net7135),
.Y(net7282)
);

AND2x2_ASAP7_75t_R c7214(
.A(net7276),
.B(net7273),
.Y(net7283)
);

NAND3x1_ASAP7_75t_R c7215(
.A(net7281),
.B(net7258),
.C(net9773),
.Y(net7284)
);

NAND3x2_ASAP7_75t_R c7216(
.B(net5414),
.C(net7248),
.A(net7238),
.Y(net7285)
);

AND2x4_ASAP7_75t_R c7217(
.A(net7212),
.B(net7270),
.Y(net7286)
);

AND2x6_ASAP7_75t_R c7218(
.A(net7285),
.B(net9971),
.Y(net7287)
);

AOI321xp33_ASAP7_75t_R c7219(
.A1(net7252),
.A2(net6303),
.A3(net7229),
.B1(net6347),
.B2(net7287),
.C(net7268),
.Y(net7288)
);

NAND3xp33_ASAP7_75t_R c7220(
.A(net7224),
.B(net7248),
.C(net9999),
.Y(net7289)
);

NOR3x1_ASAP7_75t_R c7221(
.A(net5502),
.B(net7237),
.C(net10289),
.Y(out19)
);

SDFLx1_ASAP7_75t_R c7222(
.D(net4594),
.SE(net6446),
.SI(net7233),
.CLK(clk),
.QN(net7290)
);

HAxp5_ASAP7_75t_R c7223(
.A(net6343),
.B(net7233),
.CON(net7291)
);

NOR3x2_ASAP7_75t_R c7224(
.B(net3674),
.C(net5332),
.A(net5461),
.Y(net7292)
);

NOR3xp33_ASAP7_75t_R c7225(
.A(net7147),
.B(net6391),
.C(net10260),
.Y(net7293)
);

OA21x2_ASAP7_75t_R c7226(
.A1(net6429),
.A2(net7271),
.B(net6419),
.Y(net7294)
);

OAI21x1_ASAP7_75t_R c7227(
.A1(net1774),
.A2(net7217),
.B(net5492),
.Y(net7295)
);

OAI21xp33_ASAP7_75t_R c7228(
.A1(net4469),
.A2(net7293),
.B(net6381),
.Y(net7296)
);

SDFLx2_ASAP7_75t_R c7229(
.D(net5513),
.SE(net7240),
.SI(net6887),
.CLK(clk),
.QN(net7297)
);

CKINVDCx14_ASAP7_75t_R c7230(
.A(net10339),
.Y(net7298)
);

OAI21xp5_ASAP7_75t_R c7231(
.A1(net7216),
.A2(net7136),
.B(net7237),
.Y(net7299)
);

OR3x1_ASAP7_75t_R c7232(
.A(net6303),
.B(net5443),
.C(net3316),
.Y(net7300)
);

OR3x2_ASAP7_75t_R c7233(
.A(net4573),
.B(net7290),
.C(net6391),
.Y(net7301)
);

SDFLx3_ASAP7_75t_R c7234(
.D(net6409),
.SE(net6300),
.SI(net6446),
.CLK(clk),
.QN(net7302)
);

OR3x4_ASAP7_75t_R c7235(
.A(net6427),
.B(net6384),
.C(net10289),
.Y(net7303)
);

AND3x1_ASAP7_75t_R c7236(
.A(net6391),
.B(net7232),
.C(net9773),
.Y(out8)
);

AND3x2_ASAP7_75t_R c7237(
.A(net7301),
.B(net6391),
.C(net10289),
.Y(net7304)
);

AND3x4_ASAP7_75t_R c7238(
.A(net4584),
.B(net6409),
.C(net5422),
.Y(net7305)
);

AO21x1_ASAP7_75t_R c7239(
.A1(net3655),
.A2(net7302),
.B(net4357),
.Y(net7306)
);

AO21x2_ASAP7_75t_R c7240(
.A1(net6347),
.A2(net6391),
.B(net7265),
.Y(out9)
);

AOI21x1_ASAP7_75t_R c7241(
.A1(net7217),
.A2(net6300),
.B(net6412),
.Y(net7307)
);

AOI21xp33_ASAP7_75t_R c7242(
.A1(net7043),
.A2(net5267),
.B(net7290),
.Y(net7308)
);

AOI21xp5_ASAP7_75t_R c7243(
.A1(net7237),
.A2(net7216),
.B(out9),
.Y(net7309)
);

FAx1_ASAP7_75t_R c7244(
.A(net7306),
.B(net5443),
.CI(net7183),
.SN(net7310)
);

MAJIxp5_ASAP7_75t_R c7245(
.A(net5456),
.B(net7147),
.C(net6383),
.Y(net7311)
);

MAJx2_ASAP7_75t_R c7246(
.A(net6399),
.B(net2578),
.C(net7307),
.Y(net7312)
);

MAJx3_ASAP7_75t_R c7247(
.A(net7302),
.B(net6382),
.C(net10260),
.Y(net7313)
);

NAND2x1_ASAP7_75t_R c7248(
.A(net6393),
.B(net6413),
.Y(net7314)
);

NAND3x1_ASAP7_75t_R c7249(
.A(net7291),
.B(net6409),
.C(net7311),
.Y(net7315)
);

NAND3x2_ASAP7_75t_R c7250(
.B(net6146),
.C(net7148),
.A(net6343),
.Y(net7316)
);

NOR5xp2_ASAP7_75t_R c7251(
.A(net7223),
.B(net7271),
.C(net6427),
.D(net6380),
.E(net6434),
.Y(net7317)
);

SDFLx4_ASAP7_75t_R c7252(
.D(net5198),
.SE(net7136),
.SI(net7232),
.CLK(clk),
.QN(net7318)
);

NAND3xp33_ASAP7_75t_R c7253(
.A(net7316),
.B(net3644),
.C(net10228),
.Y(net7319)
);

NOR3x1_ASAP7_75t_R c7254(
.A(net6380),
.B(net4600),
.C(net4594),
.Y(net7320)
);

NOR3x2_ASAP7_75t_R c7255(
.B(net5495),
.C(net7290),
.A(net10260),
.Y(net7321)
);

NOR3xp33_ASAP7_75t_R c7256(
.A(net6450),
.B(net7318),
.C(net10010),
.Y(net7322)
);

OA21x2_ASAP7_75t_R c7257(
.A1(net5409),
.A2(net9976),
.B(net10290),
.Y(net7323)
);

OA221x2_ASAP7_75t_R c7258(
.A1(net7322),
.A2(net6263),
.B1(net6429),
.B2(net7183),
.C(net6380),
.Y(net7324)
);

OAI21x1_ASAP7_75t_R c7259(
.A1(net5448),
.A2(net4549),
.B(net7223),
.Y(net7325)
);

OAI21xp33_ASAP7_75t_R c7260(
.A1(net7320),
.A2(net7233),
.B(net6303),
.Y(net7326)
);

OAI21xp5_ASAP7_75t_R c7261(
.A1(net7298),
.A2(net7307),
.B(net3635),
.Y(net7327)
);

OR3x1_ASAP7_75t_R c7262(
.A(net7297),
.B(net6401),
.C(net7318),
.Y(net7328)
);

DFFASRHQNx1_ASAP7_75t_R c7263(
.D(net7323),
.RESETN(net7312),
.SETN(net1774),
.CLK(clk),
.QN(net7329)
);

OAI221xp5_ASAP7_75t_R c7264(
.A1(net7296),
.A2(net7043),
.B1(net1526),
.B2(out9),
.C(net5461),
.Y(net7330)
);

OR3x2_ASAP7_75t_R c7265(
.A(net7277),
.B(net10246),
.C(net10290),
.Y(net7331)
);

OR3x4_ASAP7_75t_R c7266(
.A(net7329),
.B(net7311),
.C(net9921),
.Y(net7332)
);

AND3x1_ASAP7_75t_R c7267(
.A(net7192),
.B(net7326),
.C(net7307),
.Y(net7333)
);

AND3x2_ASAP7_75t_R c7268(
.A(net6450),
.B(net7329),
.C(net6401),
.Y(net7334)
);

AND3x4_ASAP7_75t_R c7269(
.A(net2707),
.B(net7314),
.C(out1),
.Y(net7335)
);

AO21x1_ASAP7_75t_R c7270(
.A1(net7318),
.A2(net7333),
.B(net10290),
.Y(net7336)
);

AO21x2_ASAP7_75t_R c7271(
.A1(net5422),
.A2(net7331),
.B(net4573),
.Y(net7337)
);

CKINVDCx16_ASAP7_75t_R c7272(
.A(net10339),
.Y(net7338)
);

SDFHx1_ASAP7_75t_R c7273(
.D(net6191),
.SE(net7329),
.SI(net7318),
.CLK(clk),
.QN(net7339)
);

NAND2x1p5_ASAP7_75t_R c7274(
.A(net7277),
.B(net7339),
.Y(net7340)
);

AOI21x1_ASAP7_75t_R c7275(
.A1(net3635),
.A2(net7295),
.B(net7329),
.Y(net7341)
);

AOI21xp33_ASAP7_75t_R c7276(
.A1(net6384),
.A2(net7299),
.B(net10246),
.Y(net7342)
);

AOI21xp5_ASAP7_75t_R c7277(
.A1(net7315),
.A2(net7339),
.B(net4357),
.Y(net7343)
);

FAx1_ASAP7_75t_R c7278(
.A(net6304),
.B(net5456),
.CI(net6399),
.SN(net7344)
);

MAJIxp5_ASAP7_75t_R c7279(
.A(net7305),
.B(net3644),
.C(net6434),
.Y(net7345)
);

MAJx2_ASAP7_75t_R c7280(
.A(net6304),
.B(net10005),
.C(net10008),
.Y(net7346)
);

MAJx3_ASAP7_75t_R c7281(
.A(net7346),
.B(net5527),
.C(net5513),
.Y(net7347)
);

SDFHx2_ASAP7_75t_R c7282(
.D(net6380),
.SE(net2747),
.SI(net10027),
.CLK(clk),
.QN(net7348)
);

NAND3x1_ASAP7_75t_R c7283(
.A(net4600),
.B(net6434),
.C(out9),
.Y(net7349)
);

SDFHx3_ASAP7_75t_R c7284(
.D(net7319),
.SE(net7348),
.SI(net10291),
.CLK(clk),
.QN(net7350)
);

NAND3x2_ASAP7_75t_R c7285(
.B(net5461),
.C(net6381),
.A(net9762),
.Y(net7351)
);

NAND2x2_ASAP7_75t_R c7286(
.A(net7337),
.B(net7347),
.Y(net7352)
);

NAND3xp33_ASAP7_75t_R c7287(
.A(net7350),
.B(net7340),
.C(net10041),
.Y(net7353)
);

NOR3x1_ASAP7_75t_R c7288(
.A(net7309),
.B(net7348),
.C(net9921),
.Y(net7354)
);

NOR3x2_ASAP7_75t_R c7289(
.B(net7352),
.C(net7354),
.A(net7350),
.Y(net7355)
);

OAI22xp5_ASAP7_75t_R c7290(
.A1(net7300),
.A2(net7334),
.B1(net7354),
.B2(net7318),
.Y(net7356)
);

OAI311xp33_ASAP7_75t_R c7291(
.A1(net7344),
.A2(net7350),
.A3(net7354),
.B1(out9),
.C1(net9637),
.Y(net7357)
);

OAI32xp33_ASAP7_75t_R c7292(
.A1(net5461),
.A2(net7318),
.A3(net7354),
.B1(net7232),
.B2(net9637),
.Y(net7358)
);

NOR3xp33_ASAP7_75t_R c7293(
.A(net7353),
.B(net6429),
.C(net9988),
.Y(net7359)
);

OA21x2_ASAP7_75t_R c7294(
.A1(net7348),
.A2(net7332),
.B(net7329),
.Y(net7360)
);

OAI21x1_ASAP7_75t_R c7295(
.A1(net7307),
.A2(net5866),
.B(net9983),
.Y(net7361)
);

OAI21xp33_ASAP7_75t_R c7296(
.A1(net6380),
.A2(net9901),
.B(net10072),
.Y(net7362)
);

OAI21xp5_ASAP7_75t_R c7297(
.A1(net7338),
.A2(net7297),
.B(net10060),
.Y(net7363)
);

OR3x1_ASAP7_75t_R c7298(
.A(net7327),
.B(net7329),
.C(net10049),
.Y(net7364)
);

SDFHx4_ASAP7_75t_R c7299(
.D(net7360),
.SE(net7348),
.SI(net10261),
.CLK(clk),
.QN(net7365)
);

OAI31xp33_ASAP7_75t_R c7300(
.A1(net4580),
.A2(net7342),
.A3(net7322),
.B(net7329),
.Y(net7366)
);

AOI33xp33_ASAP7_75t_R c7301(
.A1(net7290),
.A2(net6426),
.A3(net6347),
.B1(net6446),
.B2(net10010),
.B3(net10292),
.Y(net7367)
);

OR3x2_ASAP7_75t_R c7302(
.A(net7349),
.B(net5198),
.C(net10027),
.Y(net7368)
);

OR5x1_ASAP7_75t_R c7303(
.A(net6380),
.B(net7232),
.C(net10011),
.D(net10072),
.E(net10246),
.Y(net7369)
);

NAND2xp33_ASAP7_75t_R c7304(
.A(net6484),
.B(net6501),
.Y(net7370)
);

CKINVDCx20_ASAP7_75t_R c7305(
.A(net4621),
.Y(net7371)
);

CKINVDCx5p33_ASAP7_75t_R c7306(
.A(net6493),
.Y(net7372)
);

CKINVDCx6p67_ASAP7_75t_R c7307(
.A(net6477),
.Y(net7373)
);

NAND2xp5_ASAP7_75t_R c7308(
.A(net7371),
.B(net2779),
.Y(net7374)
);

CKINVDCx8_ASAP7_75t_R c7309(
.A(net6513),
.Y(net7375)
);

NAND2xp67_ASAP7_75t_R c7310(
.A(net6527),
.B(net5576),
.Y(net7376)
);

NOR2x1_ASAP7_75t_R c7311(
.A(net7370),
.B(net6465),
.Y(net7377)
);

NOR2x1p5_ASAP7_75t_R c7312(
.A(net5588),
.B(net6461),
.Y(net7378)
);

CKINVDCx9p33_ASAP7_75t_R c7313(
.A(net7375),
.Y(net7379)
);

HB1xp67_ASAP7_75t_R c7314(
.A(net6486),
.Y(net7380)
);

OR3x4_ASAP7_75t_R c7315(
.A(net6454),
.B(net6453),
.C(net7378),
.Y(net7381)
);

HB2xp67_ASAP7_75t_R c7316(
.A(net9148),
.Y(net7382)
);

HB3xp67_ASAP7_75t_R c7317(
.A(net6478),
.Y(net7383)
);

HB4xp67_ASAP7_75t_R c7318(
.A(net6453),
.Y(net7384)
);

INVx11_ASAP7_75t_R c7319(
.A(net5593),
.Y(net7385)
);

INVx13_ASAP7_75t_R c7320(
.A(net4650),
.Y(net7386)
);

INVx1_ASAP7_75t_R c7321(
.A(net6523),
.Y(net7387)
);

NOR2x2_ASAP7_75t_R c7322(
.A(net5605),
.B(net6453),
.Y(net7388)
);

NOR2xp33_ASAP7_75t_R c7323(
.A(net4652),
.B(net6505),
.Y(net7389)
);

NOR2xp67_ASAP7_75t_R c7324(
.A(net7383),
.B(net6511),
.Y(net7390)
);

INVx2_ASAP7_75t_R c7325(
.A(net9203),
.Y(net7391)
);

SDFLx1_ASAP7_75t_R c7326(
.D(net6511),
.SE(net5546),
.SI(net1833),
.CLK(clk),
.QN(net7392)
);

OR2x2_ASAP7_75t_R c7327(
.A(net2779),
.B(net4609),
.Y(net7393)
);

INVx3_ASAP7_75t_R c7328(
.A(net9658),
.Y(net7394)
);

OR2x4_ASAP7_75t_R c7329(
.A(net6501),
.B(net4650),
.Y(net7395)
);

INVx4_ASAP7_75t_R c7330(
.A(net7373),
.Y(net7396)
);

ICGx5_ASAP7_75t_R c7331(
.ENA(net6454),
.SE(net6464),
.CLK(clk),
.GCLK(net7397)
);

INVx5_ASAP7_75t_R c7332(
.A(net7394),
.Y(net7398)
);

SDFLx2_ASAP7_75t_R c7333(
.D(net7370),
.SE(net6471),
.SI(net7378),
.CLK(clk),
.QN(net7399)
);

OR2x6_ASAP7_75t_R c7334(
.A(net7379),
.B(net7383),
.Y(net7400)
);

XNOR2x1_ASAP7_75t_R c7335(
.B(net5530),
.A(net7384),
.Y(net7401)
);

INVx6_ASAP7_75t_R c7336(
.A(net9217),
.Y(net7402)
);

INVx8_ASAP7_75t_R c7337(
.A(net9288),
.Y(net7403)
);

XNOR2x2_ASAP7_75t_R c7338(
.A(net6523),
.B(net7373),
.Y(net7404)
);

INVxp33_ASAP7_75t_R c7339(
.A(net9658),
.Y(net7405)
);

INVxp67_ASAP7_75t_R c7340(
.A(net7376),
.Y(net7406)
);

BUFx10_ASAP7_75t_R c7341(
.A(net5561),
.Y(net7407)
);

BUFx12_ASAP7_75t_R c7342(
.A(net7405),
.Y(net7408)
);

AND3x1_ASAP7_75t_R c7343(
.A(net7394),
.B(net7399),
.C(net6484),
.Y(net7409)
);

BUFx12f_ASAP7_75t_R c7344(
.A(net7402),
.Y(net7410)
);

BUFx16f_ASAP7_75t_R c7345(
.A(net7376),
.Y(net7411)
);

BUFx24_ASAP7_75t_R c7346(
.A(net9288),
.Y(net7412)
);

XNOR2xp5_ASAP7_75t_R c7347(
.A(net7388),
.B(net6532),
.Y(net7413)
);

XOR2x1_ASAP7_75t_R c7348(
.A(net6456),
.B(net6521),
.Y(net7414)
);

BUFx2_ASAP7_75t_R c7349(
.A(net7391),
.Y(net7415)
);

ICGx5p33DC_ASAP7_75t_R c7350(
.ENA(net7401),
.SE(net6493),
.CLK(clk),
.GCLK(net7416)
);

ICGx6p67DC_ASAP7_75t_R c7351(
.ENA(net7415),
.SE(net7413),
.CLK(clk),
.GCLK(net7417)
);

OAI31xp67_ASAP7_75t_R c7352(
.A1(net7417),
.A2(net7370),
.A3(net7398),
.B(net6510),
.Y(net7418)
);

XOR2x2_ASAP7_75t_R c7353(
.A(net5549),
.B(net7383),
.Y(net7419)
);

AND3x2_ASAP7_75t_R c7354(
.A(net7390),
.B(net7400),
.C(net7417),
.Y(net7420)
);

BUFx3_ASAP7_75t_R c7355(
.A(net7392),
.Y(net7421)
);

BUFx4_ASAP7_75t_R c7356(
.A(net7421),
.Y(net7422)
);

ICGx8DC_ASAP7_75t_R c7357(
.ENA(net7416),
.SE(net5574),
.CLK(clk),
.GCLK(net7423)
);

BUFx4f_ASAP7_75t_R c7358(
.A(net7409),
.Y(net7424)
);

BUFx5_ASAP7_75t_R c7359(
.A(net9325),
.Y(net7425)
);

BUFx6f_ASAP7_75t_R c7360(
.A(net7384),
.Y(net7426)
);

AND3x4_ASAP7_75t_R c7361(
.A(net7396),
.B(net7415),
.C(net7420),
.Y(net7427)
);

ICGx1_ASAP7_75t_R c7362(
.ENA(net7411),
.SE(net6522),
.CLK(clk),
.GCLK(net7428)
);

BUFx8_ASAP7_75t_R c7363(
.A(net9148),
.Y(net7429)
);

XOR2xp5_ASAP7_75t_R c7364(
.A(net7398),
.B(net7414),
.Y(net7430)
);

AND2x2_ASAP7_75t_R c7365(
.A(net7430),
.B(net6482),
.Y(net7431)
);

AO21x1_ASAP7_75t_R c7366(
.A1(net7430),
.A2(net7414),
.B(net7421),
.Y(net7432)
);

OA222x2_ASAP7_75t_R c7367(
.A1(net7432),
.A2(net7427),
.B1(net7419),
.B2(net6488),
.C1(net7374),
.C2(net7378),
.Y(net7433)
);

OR4x1_ASAP7_75t_R c7368(
.A(net5539),
.B(net5605),
.C(net7422),
.D(net7415),
.Y(net7434)
);

ICGx2_ASAP7_75t_R c7369(
.ENA(net7406),
.SE(net7415),
.CLK(clk),
.GCLK(net7435)
);

AO21x2_ASAP7_75t_R c7370(
.A1(net7435),
.A2(net7404),
.B(net10293),
.Y(net7436)
);

AOI21x1_ASAP7_75t_R c7371(
.A1(net7431),
.A2(net7410),
.B(net7392),
.Y(net7437)
);

ICGx2p67DC_ASAP7_75t_R c7372(
.ENA(net7413),
.SE(net7374),
.CLK(clk),
.GCLK(net7438)
);

SDFLx3_ASAP7_75t_R c7373(
.D(net7437),
.SE(net7431),
.SI(net10293),
.CLK(clk),
.QN(net7439)
);

OR5x2_ASAP7_75t_R c7374(
.A(net7418),
.B(net7404),
.C(net7393),
.D(net7399),
.E(net7415),
.Y(net7440)
);

AOI21xp33_ASAP7_75t_R c7375(
.A1(net7434),
.A2(net7435),
.B(net7415),
.Y(net7441)
);

SDFLx4_ASAP7_75t_R c7376(
.D(net7429),
.SE(net6533),
.SI(net7441),
.CLK(clk),
.QN(net7442)
);

ICGx3_ASAP7_75t_R c7377(
.ENA(net7438),
.SE(net7441),
.CLK(clk),
.GCLK(net7443)
);

AND2x4_ASAP7_75t_R c7378(
.A(net7416),
.B(net7442),
.Y(net7444)
);

ICGx4DC_ASAP7_75t_R c7379(
.ENA(net7419),
.SE(net7423),
.CLK(clk),
.GCLK(net7445)
);

AOI21xp5_ASAP7_75t_R c7380(
.A1(net7405),
.A2(net7442),
.B(net7429),
.Y(net7446)
);

OA33x2_ASAP7_75t_R c7381(
.A1(net7437),
.A2(net7444),
.A3(net7399),
.B1(net7415),
.B2(net907),
.B3(net10249),
.Y(net7447)
);

FAx1_ASAP7_75t_R c7382(
.A(net7442),
.B(net7406),
.CI(net10295),
.SN(net7448)
);

DFFASRHQNx1_ASAP7_75t_R c7383(
.D(net7385),
.RESETN(net9776),
.SETN(net10294),
.CLK(clk),
.QN(net7449)
);

MAJIxp5_ASAP7_75t_R c7384(
.A(net7445),
.B(net7428),
.C(net10295),
.Y(net7450)
);

MAJx2_ASAP7_75t_R c7385(
.A(net7403),
.B(net7450),
.C(net7439),
.Y(net7451)
);

MAJx3_ASAP7_75t_R c7386(
.A(net7443),
.B(net7445),
.C(net10294),
.Y(net7452)
);

CKINVDCx10_ASAP7_75t_R c7387(
.A(net4724),
.Y(net7453)
);

CKINVDCx11_ASAP7_75t_R c7388(
.A(net6591),
.Y(net7454)
);

CKINVDCx12_ASAP7_75t_R c7389(
.A(net6535),
.Y(net7455)
);

AND2x6_ASAP7_75t_R c7390(
.A(net3830),
.B(net6612),
.Y(net7456)
);

CKINVDCx14_ASAP7_75t_R c7391(
.A(net9211),
.Y(net7457)
);

CKINVDCx16_ASAP7_75t_R c7392(
.A(net6471),
.Y(net7458)
);

HAxp5_ASAP7_75t_R c7393(
.A(net6503),
.B(net7451),
.CON(net7459)
);

NAND3x1_ASAP7_75t_R c7394(
.A(net7443),
.B(net7404),
.C(net6595),
.Y(net7460)
);

CKINVDCx20_ASAP7_75t_R c7395(
.A(net6477),
.Y(net7461)
);

CKINVDCx5p33_ASAP7_75t_R c7396(
.A(net9091),
.Y(net7462)
);

CKINVDCx6p67_ASAP7_75t_R c7397(
.A(net5620),
.Y(net7463)
);

SDFHx1_ASAP7_75t_R c7398(
.D(net7461),
.SE(net7380),
.SI(net9951),
.CLK(clk),
.QN(net7464)
);

CKINVDCx8_ASAP7_75t_R c7399(
.A(net9091),
.Y(net7465)
);

NAND2x1_ASAP7_75t_R c7400(
.A(net7438),
.B(net5598),
.Y(net7466)
);

CKINVDCx9p33_ASAP7_75t_R c7401(
.A(net10267),
.Y(net7467)
);

NAND2x1p5_ASAP7_75t_R c7402(
.A(net7403),
.B(net10267),
.Y(net7468)
);

HB1xp67_ASAP7_75t_R c7403(
.A(net907),
.Y(net7469)
);

HB2xp67_ASAP7_75t_R c7404(
.A(net7455),
.Y(net7470)
);

NAND2x2_ASAP7_75t_R c7405(
.A(net7464),
.B(net7469),
.Y(net7471)
);

NAND2xp33_ASAP7_75t_R c7406(
.A(net5688),
.B(net6471),
.Y(net7472)
);

HB3xp67_ASAP7_75t_R c7407(
.A(net9253),
.Y(net7473)
);

HB4xp67_ASAP7_75t_R c7408(
.A(net3705),
.Y(net7474)
);

INVx11_ASAP7_75t_R c7409(
.A(net7474),
.Y(net7475)
);

NAND3x2_ASAP7_75t_R c7410(
.B(net4762),
.C(net7464),
.A(net10267),
.Y(net7476)
);

INVx13_ASAP7_75t_R c7411(
.A(net10550),
.Y(net7477)
);

INVx1_ASAP7_75t_R c7412(
.A(net6557),
.Y(net7478)
);

NAND2xp5_ASAP7_75t_R c7413(
.A(net7475),
.B(net5636),
.Y(net7479)
);

NAND2xp67_ASAP7_75t_R c7414(
.A(net6465),
.B(net10279),
.Y(net7480)
);

INVx2_ASAP7_75t_R c7415(
.A(net10437),
.Y(net7481)
);

INVx3_ASAP7_75t_R c7416(
.A(net10400),
.Y(net7482)
);

NAND3xp33_ASAP7_75t_R c7417(
.A(net7412),
.B(net7476),
.C(net5532),
.Y(net7483)
);

NOR3x1_ASAP7_75t_R c7418(
.A(net7467),
.B(net7469),
.C(net6461),
.Y(net7484)
);

NOR2x1_ASAP7_75t_R c7419(
.A(net7458),
.B(net7438),
.Y(net7485)
);

INVx4_ASAP7_75t_R c7420(
.A(net10559),
.Y(net7486)
);

INVx5_ASAP7_75t_R c7421(
.A(net7462),
.Y(net7487)
);

INVx6_ASAP7_75t_R c7422(
.A(net7478),
.Y(net7488)
);

NOR2x1p5_ASAP7_75t_R c7423(
.A(net7487),
.B(net7456),
.Y(net7489)
);

INVx8_ASAP7_75t_R c7424(
.A(net7372),
.Y(net7490)
);

NOR2x2_ASAP7_75t_R c7425(
.A(net7472),
.B(net5688),
.Y(net7491)
);

NOR3x2_ASAP7_75t_R c7426(
.B(net7460),
.C(net7372),
.A(net7412),
.Y(net7492)
);

INVxp33_ASAP7_75t_R c7427(
.A(net6461),
.Y(net7493)
);

INVxp67_ASAP7_75t_R c7428(
.A(net6535),
.Y(net7494)
);

BUFx10_ASAP7_75t_R c7429(
.A(net7480),
.Y(net7495)
);

NOR3xp33_ASAP7_75t_R c7430(
.A(net4696),
.B(net7453),
.C(net7475),
.Y(net7496)
);

BUFx12_ASAP7_75t_R c7431(
.A(net7468),
.Y(net7497)
);

NOR2xp33_ASAP7_75t_R c7432(
.A(net7465),
.B(net6550),
.Y(net7498)
);

NOR2xp67_ASAP7_75t_R c7433(
.A(net7490),
.B(net7496),
.Y(net7499)
);

BUFx12f_ASAP7_75t_R c7434(
.A(net7495),
.Y(net7500)
);

OR2x2_ASAP7_75t_R c7435(
.A(net7496),
.B(net7446),
.Y(net7501)
);

OR2x4_ASAP7_75t_R c7436(
.A(net7457),
.B(net6557),
.Y(net7502)
);

OA21x2_ASAP7_75t_R c7437(
.A1(net7451),
.A2(net7495),
.B(net6612),
.Y(net7503)
);

BUFx16f_ASAP7_75t_R c7438(
.A(net7446),
.Y(net7504)
);

OR2x6_ASAP7_75t_R c7439(
.A(net7501),
.B(net7492),
.Y(net7505)
);

XNOR2x1_ASAP7_75t_R c7440(
.B(net7471),
.A(net7500),
.Y(net7506)
);

XNOR2x2_ASAP7_75t_R c7441(
.A(net6550),
.B(net7496),
.Y(net7507)
);

BUFx24_ASAP7_75t_R c7442(
.A(net7500),
.Y(net7508)
);

XNOR2xp5_ASAP7_75t_R c7443(
.A(net7498),
.B(net7492),
.Y(net7509)
);

XOR2x1_ASAP7_75t_R c7444(
.A(net5649),
.B(net5628),
.Y(net7510)
);

ICGx4_ASAP7_75t_R c7445(
.ENA(net7484),
.SE(net7390),
.CLK(clk),
.GCLK(net7511)
);

XOR2x2_ASAP7_75t_R c7446(
.A(net7495),
.B(net7510),
.Y(net7512)
);

XOR2xp5_ASAP7_75t_R c7447(
.A(net7400),
.B(net7508),
.Y(net7513)
);

BUFx2_ASAP7_75t_R c7448(
.A(net7482),
.Y(net7514)
);

AND2x2_ASAP7_75t_R c7449(
.A(net7509),
.B(net7503),
.Y(net7515)
);

BUFx3_ASAP7_75t_R c7450(
.A(net7497),
.Y(net7516)
);

AND2x4_ASAP7_75t_R c7451(
.A(net7515),
.B(net7463),
.Y(net7517)
);

AND2x6_ASAP7_75t_R c7452(
.A(net7504),
.B(net7517),
.Y(net7518)
);

OAI21x1_ASAP7_75t_R c7453(
.A1(net7454),
.A2(net7516),
.B(net6615),
.Y(net7519)
);

BUFx4_ASAP7_75t_R c7454(
.A(net10487),
.Y(net7520)
);

OR4x2_ASAP7_75t_R c7455(
.A(net7503),
.B(net7511),
.C(net7508),
.D(net7378),
.Y(net7521)
);

HAxp5_ASAP7_75t_R c7456(
.A(net7517),
.B(net7508),
.CON(net7523),
.SN(net7522)
);

A2O1A1Ixp33_ASAP7_75t_R c7457(
.A1(net7511),
.A2(net7425),
.B(net6554),
.C(net7469),
.Y(net7524)
);

NAND2x1_ASAP7_75t_R c7458(
.A(net7375),
.B(net7503),
.Y(net7525)
);

SDFHx2_ASAP7_75t_R c7459(
.D(net7520),
.SE(net7523),
.SI(net7496),
.CLK(clk),
.QN(net7526)
);

OAI21xp33_ASAP7_75t_R c7460(
.A1(net7507),
.A2(net7517),
.B(net7510),
.Y(net7527)
);

OAI21xp5_ASAP7_75t_R c7461(
.A1(net7463),
.A2(net7509),
.B(net7510),
.Y(net7528)
);

NAND2x1p5_ASAP7_75t_R c7462(
.A(net7512),
.B(net7387),
.Y(net7529)
);

NAND2x2_ASAP7_75t_R c7463(
.A(net7489),
.B(net7526),
.Y(net7530)
);

OR3x1_ASAP7_75t_R c7464(
.A(net7476),
.B(net7516),
.C(net7529),
.Y(net7531)
);

OR3x2_ASAP7_75t_R c7465(
.A(net7519),
.B(net7511),
.C(net7492),
.Y(net7532)
);

NAND2xp33_ASAP7_75t_R c7466(
.A(net9908),
.B(net10296),
.Y(net7533)
);

OR3x4_ASAP7_75t_R c7467(
.A(net137),
.B(net7533),
.C(net7529),
.Y(net7534)
);

A2O1A1O1Ixp25_ASAP7_75t_R c7468(
.A1(net7529),
.A2(net7509),
.B(net7533),
.C(net7534),
.D(net6508),
.Y(net7535)
);

AND5x1_ASAP7_75t_R c7469(
.A(net7470),
.B(net7533),
.C(net7534),
.D(net6612),
.E(net10297),
.Y(net7536)
);

BUFx4f_ASAP7_75t_R c7470(
.A(net9235),
.Y(net7537)
);

BUFx5_ASAP7_75t_R c7471(
.A(net10123),
.Y(net7538)
);

BUFx6f_ASAP7_75t_R c7472(
.A(net10509),
.Y(net7539)
);

SDFHx3_ASAP7_75t_R c7473(
.D(net7493),
.SE(net7494),
.SI(net10267),
.CLK(clk),
.QN(net7540)
);

NAND2xp5_ASAP7_75t_R c7474(
.A(net6691),
.B(net7540),
.Y(net7541)
);

BUFx8_ASAP7_75t_R c7475(
.A(net6635),
.Y(net7542)
);

CKINVDCx10_ASAP7_75t_R c7476(
.A(net7435),
.Y(net7543)
);

NAND2xp67_ASAP7_75t_R c7477(
.A(net7449),
.B(net7543),
.Y(net7544)
);

CKINVDCx11_ASAP7_75t_R c7478(
.A(net5718),
.Y(net7545)
);

CKINVDCx12_ASAP7_75t_R c7479(
.A(net7491),
.Y(net7546)
);

CKINVDCx14_ASAP7_75t_R c7480(
.A(net9993),
.Y(net7547)
);

NOR2x1_ASAP7_75t_R c7481(
.A(net6532),
.B(net4827),
.Y(net7548)
);

NOR2x1p5_ASAP7_75t_R c7482(
.A(net6644),
.B(net7461),
.Y(net7549)
);

CKINVDCx16_ASAP7_75t_R c7483(
.A(net9177),
.Y(net7550)
);

CKINVDCx20_ASAP7_75t_R c7484(
.A(net7450),
.Y(net7551)
);

CKINVDCx5p33_ASAP7_75t_R c7485(
.A(net10486),
.Y(net7552)
);

NOR2x2_ASAP7_75t_R c7486(
.A(net7552),
.B(net6684),
.Y(net7553)
);

NOR2xp33_ASAP7_75t_R c7487(
.A(net5771),
.B(net7543),
.Y(net7554)
);

NOR2xp67_ASAP7_75t_R c7488(
.A(net6506),
.B(net7449),
.Y(net7555)
);

AND3x1_ASAP7_75t_R c7489(
.A(net7488),
.B(net5598),
.C(net7540),
.Y(net7556)
);

OR2x2_ASAP7_75t_R c7490(
.A(net5738),
.B(net7435),
.Y(net7557)
);

OR2x4_ASAP7_75t_R c7491(
.A(net6684),
.B(net4738),
.Y(net7558)
);

OR2x6_ASAP7_75t_R c7492(
.A(net7486),
.B(net5689),
.Y(net7559)
);

CKINVDCx6p67_ASAP7_75t_R c7493(
.A(net7545),
.Y(net7560)
);

XNOR2x1_ASAP7_75t_R c7494(
.B(net7528),
.A(net7544),
.Y(net7561)
);

AND3x2_ASAP7_75t_R c7495(
.A(net7557),
.B(net7548),
.C(net6643),
.Y(net7562)
);

CKINVDCx8_ASAP7_75t_R c7496(
.A(net9325),
.Y(net7563)
);

XNOR2x2_ASAP7_75t_R c7497(
.A(net3767),
.B(net7559),
.Y(net7564)
);

CKINVDCx9p33_ASAP7_75t_R c7498(
.A(net9216),
.Y(net7565)
);

HB1xp67_ASAP7_75t_R c7499(
.A(net7530),
.Y(net7566)
);

HB2xp67_ASAP7_75t_R c7500(
.A(net10513),
.Y(net7567)
);

XNOR2xp5_ASAP7_75t_R c7501(
.A(net7560),
.B(net7549),
.Y(net7568)
);

XOR2x1_ASAP7_75t_R c7502(
.A(net7516),
.B(net7540),
.Y(net7569)
);

HB3xp67_ASAP7_75t_R c7503(
.A(net10458),
.Y(net7570)
);

HB4xp67_ASAP7_75t_R c7504(
.A(net9667),
.Y(net7571)
);

XOR2x2_ASAP7_75t_R c7505(
.A(net7537),
.B(net6569),
.Y(net7572)
);

XOR2xp5_ASAP7_75t_R c7506(
.A(net7556),
.B(net6681),
.Y(net7573)
);

AND3x4_ASAP7_75t_R c7507(
.A(net6561),
.B(net7486),
.C(net6681),
.Y(net7574)
);

AO21x1_ASAP7_75t_R c7508(
.A1(net4834),
.A2(net7564),
.B(net9719),
.Y(net7575)
);

AND2x2_ASAP7_75t_R c7509(
.A(net6616),
.B(net7537),
.Y(net7576)
);

INVx11_ASAP7_75t_R c7510(
.A(net9667),
.Y(net7577)
);

AO21x2_ASAP7_75t_R c7511(
.A1(net7554),
.A2(net7576),
.B(net7534),
.Y(net7578)
);

INVx13_ASAP7_75t_R c7512(
.A(net7551),
.Y(net7579)
);

AOI21x1_ASAP7_75t_R c7513(
.A1(net7563),
.A2(net7564),
.B(net10116),
.Y(net7580)
);

INVx1_ASAP7_75t_R c7514(
.A(net10503),
.Y(net7581)
);

INVx2_ASAP7_75t_R c7515(
.A(net6676),
.Y(net7582)
);

INVx3_ASAP7_75t_R c7516(
.A(net10093),
.Y(net7583)
);

AND2x4_ASAP7_75t_R c7517(
.A(net6585),
.B(net6561),
.Y(net7584)
);

AND2x6_ASAP7_75t_R c7518(
.A(net6522),
.B(net7450),
.Y(net7585)
);

INVx4_ASAP7_75t_R c7519(
.A(net7565),
.Y(net7586)
);

AOI21xp33_ASAP7_75t_R c7520(
.A1(net6629),
.A2(net7578),
.B(net7399),
.Y(net7587)
);

HAxp5_ASAP7_75t_R c7521(
.A(net7469),
.B(net10171),
.CON(net7588)
);

INVx5_ASAP7_75t_R c7522(
.A(net9177),
.Y(net7589)
);

NAND2x1_ASAP7_75t_R c7523(
.A(net5730),
.B(net7426),
.Y(net7590)
);

AOI21xp5_ASAP7_75t_R c7524(
.A1(net7436),
.A2(net6666),
.B(net10050),
.Y(net7591)
);

NAND2x1p5_ASAP7_75t_R c7525(
.A(net6487),
.B(net7581),
.Y(net7592)
);

NAND2x2_ASAP7_75t_R c7526(
.A(net7410),
.B(net7583),
.Y(net7593)
);

INVx6_ASAP7_75t_R c7527(
.A(net7569),
.Y(net7594)
);

FAx1_ASAP7_75t_R c7528(
.A(net7583),
.B(net7573),
.CI(net9642),
.SN(net7595)
);

NAND2xp33_ASAP7_75t_R c7529(
.A(net7553),
.B(net7583),
.Y(net7596)
);

AND4x1_ASAP7_75t_R c7530(
.A(net7594),
.B(net7592),
.C(net7532),
.D(net7435),
.Y(net7597)
);

MAJIxp5_ASAP7_75t_R c7531(
.A(net7548),
.B(net7494),
.C(net6635),
.Y(net7598)
);

MAJx2_ASAP7_75t_R c7532(
.A(net7572),
.B(net7548),
.C(net6624),
.Y(net7599)
);

NAND2xp5_ASAP7_75t_R c7533(
.A(net7510),
.B(net7543),
.Y(net7600)
);

NAND2xp67_ASAP7_75t_R c7534(
.A(net7586),
.B(net10116),
.Y(net7601)
);

INVx8_ASAP7_75t_R c7535(
.A(net7595),
.Y(net7602)
);

NOR2x1_ASAP7_75t_R c7536(
.A(net7586),
.B(net9675),
.Y(net7603)
);

NOR2x1p5_ASAP7_75t_R c7537(
.A(net7589),
.B(net10050),
.Y(net7604)
);

SDFHx4_ASAP7_75t_R c7538(
.D(net7575),
.SE(net7576),
.SI(net7578),
.CLK(clk),
.QN(net7605)
);

NOR2x2_ASAP7_75t_R c7539(
.A(net7563),
.B(net7542),
.Y(net7606)
);

MAJx3_ASAP7_75t_R c7540(
.A(net5725),
.B(net7606),
.C(net7597),
.Y(net7607)
);

AND5x2_ASAP7_75t_R c7541(
.A(net7543),
.B(net7585),
.C(net4738),
.D(net7544),
.E(net7435),
.Y(net7608)
);

INVxp33_ASAP7_75t_R c7542(
.A(net10509),
.Y(net7609)
);

NAND3x1_ASAP7_75t_R c7543(
.A(net7556),
.B(net7542),
.C(net10123),
.Y(net7610)
);

NAND3x2_ASAP7_75t_R c7544(
.B(net7603),
.C(net7600),
.A(net7593),
.Y(net7611)
);

AND4x2_ASAP7_75t_R c7545(
.A(net7548),
.B(net7605),
.C(net6669),
.D(net9785),
.Y(net7612)
);

NAND3xp33_ASAP7_75t_R c7546(
.A(net7608),
.B(net7605),
.C(net4845),
.Y(net7613)
);

INVxp67_ASAP7_75t_R c7547(
.A(net10123),
.Y(net7614)
);

NOR2xp33_ASAP7_75t_R c7548(
.A(net7610),
.B(net7614),
.Y(net7615)
);

AO211x2_ASAP7_75t_R c7549(
.A1(net7555),
.A2(net7614),
.B(net7615),
.C(net4827),
.Y(net7616)
);

NOR3x1_ASAP7_75t_R c7550(
.A(net7425),
.B(net7435),
.C(net10028),
.Y(net7617)
);

AO221x1_ASAP7_75t_R c7551(
.A1(net7538),
.A2(net7616),
.B1(net7605),
.B2(net7617),
.C(net7399),
.Y(net7618)
);

AO221x2_ASAP7_75t_R c7552(
.A1(net7609),
.A2(net7596),
.B1(net7615),
.B2(net7618),
.C(net7544),
.Y(net7619)
);

NOR2xp67_ASAP7_75t_R c7553(
.A(net7532),
.B(net6782),
.Y(net7620)
);

OR2x2_ASAP7_75t_R c7554(
.A(net6658),
.B(net6649),
.Y(net7621)
);

OR2x4_ASAP7_75t_R c7555(
.A(net7492),
.B(net7550),
.Y(net7622)
);

OR2x6_ASAP7_75t_R c7556(
.A(net7622),
.B(net7581),
.Y(net7623)
);

XNOR2x1_ASAP7_75t_R c7557(
.B(net7436),
.A(net6658),
.Y(net7624)
);

XNOR2x2_ASAP7_75t_R c7558(
.A(net6482),
.B(net7473),
.Y(net7625)
);

XNOR2xp5_ASAP7_75t_R c7559(
.A(net3034),
.B(net5779),
.Y(net7626)
);

XOR2x1_ASAP7_75t_R c7560(
.A(net7623),
.B(net7542),
.Y(net7627)
);

XOR2x2_ASAP7_75t_R c7561(
.A(net7621),
.B(net7624),
.Y(net7628)
);

XOR2xp5_ASAP7_75t_R c7562(
.A(net4749),
.B(net6773),
.Y(net7629)
);

AND2x2_ASAP7_75t_R c7563(
.A(net7588),
.B(net6482),
.Y(net7630)
);

BUFx10_ASAP7_75t_R c7564(
.A(net10431),
.Y(net7631)
);

AND2x4_ASAP7_75t_R c7565(
.A(net7626),
.B(net7630),
.Y(net7632)
);

AND2x6_ASAP7_75t_R c7566(
.A(net7631),
.B(net10298),
.Y(net7633)
);

BUFx12_ASAP7_75t_R c7567(
.A(net6738),
.Y(net7634)
);

NOR3x2_ASAP7_75t_R c7568(
.B(net6569),
.C(net7620),
.A(net7466),
.Y(net7635)
);

HAxp5_ASAP7_75t_R c7569(
.A(net7625),
.B(net7633),
.CON(net7637),
.SN(net7636)
);

BUFx12f_ASAP7_75t_R c7570(
.A(net10053),
.Y(net7638)
);

NAND2x1_ASAP7_75t_R c7571(
.A(net6600),
.B(net7583),
.Y(net7639)
);

NAND2x1p5_ASAP7_75t_R c7572(
.A(net7505),
.B(net7573),
.Y(net7640)
);

NAND2x2_ASAP7_75t_R c7573(
.A(net7633),
.B(net7621),
.Y(net7641)
);

NAND2xp33_ASAP7_75t_R c7574(
.A(net7630),
.B(net7576),
.Y(net7642)
);

ICGx5_ASAP7_75t_R c7575(
.ENA(net6718),
.SE(net6738),
.CLK(clk),
.GCLK(net7643)
);

BUFx16f_ASAP7_75t_R c7576(
.A(net7635),
.Y(net7644)
);

BUFx24_ASAP7_75t_R c7577(
.A(net7539),
.Y(net7645)
);

AO22x1_ASAP7_75t_R c7578(
.A1(net7581),
.A2(net6777),
.B1(net7506),
.B2(net6764),
.Y(net7646)
);

NAND2xp5_ASAP7_75t_R c7579(
.A(net7627),
.B(net7559),
.Y(net7647)
);

NAND2xp67_ASAP7_75t_R c7580(
.A(net7643),
.B(net7645),
.Y(net7648)
);

NOR2x1_ASAP7_75t_R c7581(
.A(net6642),
.B(net7606),
.Y(net7649)
);

NOR2x1p5_ASAP7_75t_R c7582(
.A(net7628),
.B(net7559),
.Y(net7650)
);

NOR2x2_ASAP7_75t_R c7583(
.A(net7633),
.B(net10298),
.Y(net7651)
);

NOR2xp33_ASAP7_75t_R c7584(
.A(net7634),
.B(net7611),
.Y(net7652)
);

NOR2xp67_ASAP7_75t_R c7585(
.A(net7624),
.B(net6714),
.Y(net7653)
);

OR2x2_ASAP7_75t_R c7586(
.A(net7644),
.B(net6714),
.Y(net7654)
);

BUFx2_ASAP7_75t_R c7587(
.A(net7654),
.Y(net7655)
);

NOR3xp33_ASAP7_75t_R c7588(
.A(net6595),
.B(net7532),
.C(net7651),
.Y(net7656)
);

OR2x4_ASAP7_75t_R c7589(
.A(net7656),
.B(net6642),
.Y(net7657)
);

OA21x2_ASAP7_75t_R c7590(
.A1(net4738),
.A2(net7643),
.B(net7622),
.Y(net7658)
);

BUFx3_ASAP7_75t_R c7591(
.A(net10410),
.Y(net7659)
);

OR2x6_ASAP7_75t_R c7592(
.A(net7579),
.B(net7645),
.Y(net7660)
);

BUFx4_ASAP7_75t_R c7593(
.A(net10501),
.Y(net7661)
);

XNOR2x1_ASAP7_75t_R c7594(
.B(net7648),
.A(net7652),
.Y(net7662)
);

SDFLx1_ASAP7_75t_R c7595(
.D(net7484),
.SE(net6669),
.SI(net7622),
.CLK(clk),
.QN(net7663)
);

XNOR2x2_ASAP7_75t_R c7596(
.A(net6669),
.B(net7597),
.Y(net7664)
);

SDFLx2_ASAP7_75t_R c7597(
.D(net7662),
.SE(net6595),
.SI(net7574),
.CLK(clk),
.QN(net7665)
);

AO22x2_ASAP7_75t_R c7598(
.A1(net6777),
.A2(net7661),
.B1(net7621),
.B2(net7658),
.Y(net7666)
);

XNOR2xp5_ASAP7_75t_R c7599(
.A(net7596),
.B(net6738),
.Y(net7667)
);

XOR2x1_ASAP7_75t_R c7600(
.A(net7559),
.B(net5841),
.Y(net7668)
);

ICGx5p33DC_ASAP7_75t_R c7601(
.ENA(net6747),
.SE(net9642),
.CLK(clk),
.GCLK(net7669)
);

XOR2x2_ASAP7_75t_R c7602(
.A(net7629),
.B(net7667),
.Y(net7670)
);

XOR2xp5_ASAP7_75t_R c7603(
.A(net7506),
.B(net7573),
.Y(net7671)
);

BUFx4f_ASAP7_75t_R c7604(
.A(net10360),
.Y(net7672)
);

AO31x2_ASAP7_75t_R c7605(
.A1(net7672),
.A2(net4940),
.A3(net5689),
.B(net7669),
.Y(net7673)
);

AND2x2_ASAP7_75t_R c7606(
.A(net7665),
.B(net7652),
.Y(net7674)
);

AND2x4_ASAP7_75t_R c7607(
.A(net4940),
.B(net4845),
.Y(net7675)
);

AND2x6_ASAP7_75t_R c7608(
.A(net7649),
.B(net7667),
.Y(net7676)
);

HAxp5_ASAP7_75t_R c7609(
.A(net7646),
.B(net7665),
.CON(net7677)
);

BUFx5_ASAP7_75t_R c7610(
.A(net10463),
.Y(net7678)
);

NAND2x1_ASAP7_75t_R c7611(
.A(net7502),
.B(net4749),
.Y(net7679)
);

AOI211x1_ASAP7_75t_R c7612(
.A1(net7632),
.A2(net7677),
.B(net4870),
.C(net7618),
.Y(net7680)
);

OAI21x1_ASAP7_75t_R c7613(
.A1(net5726),
.A2(net7663),
.B(net10099),
.Y(net7681)
);

NAND2x1p5_ASAP7_75t_R c7614(
.A(net7681),
.B(net7673),
.Y(net7682)
);

NAND2x2_ASAP7_75t_R c7615(
.A(net7577),
.B(net7645),
.Y(net7683)
);

AO32x1_ASAP7_75t_R c7616(
.A1(net7439),
.A2(net6600),
.A3(net6747),
.B1(net7622),
.B2(net7651),
.Y(net7684)
);

BUFx6f_ASAP7_75t_R c7617(
.A(net10128),
.Y(net7685)
);

NAND2xp33_ASAP7_75t_R c7618(
.A(net7685),
.B(net10299),
.Y(net7686)
);

SDFLx3_ASAP7_75t_R c7619(
.D(net7661),
.SE(net6747),
.SI(net7673),
.CLK(clk),
.QN(net7687)
);

OAI21xp33_ASAP7_75t_R c7620(
.A1(net5598),
.A2(net7456),
.B(net7667),
.Y(net7688)
);

NAND2xp5_ASAP7_75t_R c7621(
.A(net7660),
.B(net7687),
.Y(net7689)
);

OAI21xp5_ASAP7_75t_R c7622(
.A1(net6773),
.A2(net7633),
.B(net7678),
.Y(net7690)
);

OR3x1_ASAP7_75t_R c7623(
.A(net7639),
.B(net7688),
.C(net7687),
.Y(net7691)
);

OAI222xp33_ASAP7_75t_R c7624(
.A1(net7679),
.A2(net7687),
.B1(net4940),
.B2(net7651),
.C1(net7469),
.C2(net10023),
.Y(net7692)
);

NAND2xp67_ASAP7_75t_R c7625(
.A(net7678),
.B(net7690),
.Y(net7693)
);

AOI211xp5_ASAP7_75t_R c7626(
.A1(net7663),
.A2(net7685),
.B(net7662),
.C(net10299),
.Y(net7694)
);

OR3x2_ASAP7_75t_R c7627(
.A(net7693),
.B(net7690),
.C(net10146),
.Y(net7695)
);

BUFx8_ASAP7_75t_R c7628(
.A(net10053),
.Y(net7696)
);

OR3x4_ASAP7_75t_R c7629(
.A(net6666),
.B(net7436),
.C(net10023),
.Y(net7697)
);

AND3x1_ASAP7_75t_R c7630(
.A(net7689),
.B(net7673),
.C(net9979),
.Y(net7698)
);

AOI22x1_ASAP7_75t_R c7631(
.A1(net7688),
.A2(net7686),
.B1(net6705),
.B2(net9979),
.Y(net7699)
);

NOR2x1_ASAP7_75t_R c7632(
.A(net7671),
.B(net7698),
.Y(net7700)
);

AND3x2_ASAP7_75t_R c7633(
.A(net7692),
.B(net7700),
.C(net7688),
.Y(net7701)
);

OAI321xp33_ASAP7_75t_R c7634(
.A1(net7669),
.A2(net7670),
.A3(net7667),
.B1(net7673),
.B2(net7651),
.C(net10134),
.Y(net7702)
);

AND3x4_ASAP7_75t_R c7635(
.A(net7700),
.B(net6760),
.C(net7670),
.Y(net7703)
);

NOR2x1p5_ASAP7_75t_R c7636(
.A(net7696),
.B(net6519),
.Y(net7704)
);

NOR2x2_ASAP7_75t_R c7637(
.A(net5858),
.B(net7564),
.Y(net7705)
);

AO21x1_ASAP7_75t_R c7638(
.A1(net7690),
.A2(net6825),
.B(net7481),
.Y(net7706)
);

NOR2xp33_ASAP7_75t_R c7639(
.A(net6719),
.B(net7673),
.Y(net7707)
);

AOI22xp33_ASAP7_75t_R c7640(
.A1(net6618),
.A2(net4870),
.B1(net5879),
.B2(net5910),
.Y(net7708)
);

CKINVDCx10_ASAP7_75t_R c7641(
.A(net7673),
.Y(net7709)
);

NOR2xp67_ASAP7_75t_R c7642(
.A(net7524),
.B(net7708),
.Y(net7710)
);

CKINVDCx11_ASAP7_75t_R c7643(
.A(net10157),
.Y(net7711)
);

OR2x2_ASAP7_75t_R c7644(
.A(net6838),
.B(net7696),
.Y(net7712)
);

CKINVDCx12_ASAP7_75t_R c7645(
.A(net10333),
.Y(net7713)
);

AO21x2_ASAP7_75t_R c7646(
.A1(net7699),
.A2(net10081),
.B(net10281),
.Y(net7714)
);

OR2x4_ASAP7_75t_R c7647(
.A(net7690),
.B(net9818),
.Y(net7715)
);

OR2x6_ASAP7_75t_R c7648(
.A(net7546),
.B(net7704),
.Y(net7716)
);

XNOR2x1_ASAP7_75t_R c7649(
.B(net5910),
.A(net9841),
.Y(net7717)
);

XNOR2x2_ASAP7_75t_R c7650(
.A(net7713),
.B(net5836),
.Y(net7718)
);

XNOR2xp5_ASAP7_75t_R c7651(
.A(net6798),
.B(net6795),
.Y(net7719)
);

XOR2x1_ASAP7_75t_R c7652(
.A(net2163),
.B(net7645),
.Y(net7720)
);

CKINVDCx14_ASAP7_75t_R c7653(
.A(net7719),
.Y(net7721)
);

XOR2x2_ASAP7_75t_R c7654(
.A(net7717),
.B(net10296),
.Y(net7722)
);

CKINVDCx16_ASAP7_75t_R c7655(
.A(net10471),
.Y(net7723)
);

XOR2xp5_ASAP7_75t_R c7656(
.A(net7711),
.B(net7481),
.Y(net7724)
);

AOI21x1_ASAP7_75t_R c7657(
.A1(net6788),
.A2(net7668),
.B(net7456),
.Y(net7725)
);

CKINVDCx20_ASAP7_75t_R c7658(
.A(net4870),
.Y(net7726)
);

CKINVDCx5p33_ASAP7_75t_R c7659(
.A(net10369),
.Y(net7727)
);

CKINVDCx6p67_ASAP7_75t_R c7660(
.A(net10117),
.Y(net7728)
);

AND2x2_ASAP7_75t_R c7661(
.A(net5879),
.B(net7606),
.Y(net7729)
);

AND2x4_ASAP7_75t_R c7662(
.A(net4099),
.B(net9774),
.Y(net7730)
);

CKINVDCx8_ASAP7_75t_R c7663(
.A(net10543),
.Y(net7731)
);

AND2x6_ASAP7_75t_R c7664(
.A(net6869),
.B(net9876),
.Y(net7732)
);

HAxp5_ASAP7_75t_R c7665(
.A(net7718),
.B(net7466),
.CON(net7734),
.SN(net7733)
);

ICGx6p67DC_ASAP7_75t_R c7666(
.ENA(net7604),
.SE(net6870),
.CLK(clk),
.GCLK(net7735)
);

NAND2x1_ASAP7_75t_R c7667(
.A(net6714),
.B(net7735),
.Y(net7736)
);

NAND2x1p5_ASAP7_75t_R c7668(
.A(net7652),
.B(net6825),
.Y(net7737)
);

AOI21xp33_ASAP7_75t_R c7669(
.A1(net7722),
.A2(net4962),
.B(net6796),
.Y(net7738)
);

NAND2x2_ASAP7_75t_R c7670(
.A(net7730),
.B(net2163),
.Y(net7739)
);

NAND2xp33_ASAP7_75t_R c7671(
.A(net7602),
.B(net6868),
.Y(net7740)
);

AOI21xp5_ASAP7_75t_R c7672(
.A1(net7725),
.A2(net5836),
.B(net7734),
.Y(net7741)
);

NAND2xp5_ASAP7_75t_R c7673(
.A(net7739),
.B(net6847),
.Y(net7742)
);

CKINVDCx9p33_ASAP7_75t_R c7674(
.A(net10533),
.Y(net7743)
);

HB1xp67_ASAP7_75t_R c7675(
.A(net10103),
.Y(net7744)
);

NAND2xp67_ASAP7_75t_R c7676(
.A(net6843),
.B(net7725),
.Y(net7745)
);

FAx1_ASAP7_75t_R c7677(
.A(net7734),
.B(net7686),
.CI(net10299),
.SN(net7746)
);

ICGx8DC_ASAP7_75t_R c7678(
.ENA(net7715),
.SE(net6832),
.CLK(clk),
.GCLK(net7747)
);

NOR2x1_ASAP7_75t_R c7679(
.A(net6868),
.B(net6852),
.Y(out13)
);

NOR2x1p5_ASAP7_75t_R c7680(
.A(net7736),
.B(net4652),
.Y(net7748)
);

NOR2x2_ASAP7_75t_R c7681(
.A(net5010),
.B(net2163),
.Y(net7749)
);

NOR2xp33_ASAP7_75t_R c7682(
.A(net7744),
.B(net7749),
.Y(net7750)
);

NOR2xp67_ASAP7_75t_R c7683(
.A(net7645),
.B(net7747),
.Y(net7751)
);

OR2x2_ASAP7_75t_R c7684(
.A(net7743),
.B(net6618),
.Y(net7752)
);

HB2xp67_ASAP7_75t_R c7685(
.A(net10401),
.Y(net7753)
);

ICGx1_ASAP7_75t_R c7686(
.ENA(net7737),
.SE(net7477),
.CLK(clk),
.GCLK(net7754)
);

HB3xp67_ASAP7_75t_R c7687(
.A(net10534),
.Y(net7755)
);

AO32x2_ASAP7_75t_R c7688(
.A1(net4065),
.A2(net7586),
.A3(net7753),
.B1(net7704),
.B2(net7721),
.Y(net7756)
);

SDFLx4_ASAP7_75t_R c7689(
.D(net7378),
.SE(net7750),
.SI(net7749),
.CLK(clk),
.QN(net7757)
);

MAJIxp5_ASAP7_75t_R c7690(
.A(net7731),
.B(net7726),
.C(net7704),
.Y(net7758)
);

AOI221x1_ASAP7_75t_R c7691(
.A1(net7753),
.A2(net6787),
.B1(net7733),
.B2(out13),
.C(net7651),
.Y(net7759)
);

HB4xp67_ASAP7_75t_R c7692(
.A(net10359),
.Y(net7760)
);

OR2x4_ASAP7_75t_R c7693(
.A(net7748),
.B(net7711),
.Y(net7761)
);

OR2x6_ASAP7_75t_R c7694(
.A(net7740),
.B(net6795),
.Y(net7762)
);

INVx11_ASAP7_75t_R c7695(
.A(net10439),
.Y(net7763)
);

XNOR2x1_ASAP7_75t_R c7696(
.B(net7757),
.A(net7712),
.Y(net7764)
);

MAJx2_ASAP7_75t_R c7697(
.A(net6825),
.B(net7762),
.C(net7757),
.Y(net7765)
);

XNOR2x2_ASAP7_75t_R c7698(
.A(net7752),
.B(net6868),
.Y(net7766)
);

XNOR2xp5_ASAP7_75t_R c7699(
.A(net7766),
.B(net7757),
.Y(net7767)
);

MAJx3_ASAP7_75t_R c7700(
.A(net7650),
.B(net7767),
.C(net6624),
.Y(net7768)
);

INVx13_ASAP7_75t_R c7701(
.A(net10360),
.Y(net7769)
);

INVx1_ASAP7_75t_R c7702(
.A(net10333),
.Y(net7770)
);

NAND3x1_ASAP7_75t_R c7703(
.A(net7756),
.B(net7752),
.C(net7764),
.Y(net7771)
);

NAND3x2_ASAP7_75t_R c7704(
.B(net7723),
.C(net7640),
.A(net7751),
.Y(net7772)
);

NAND3xp33_ASAP7_75t_R c7705(
.A(net4951),
.B(net7765),
.C(net7705),
.Y(net7773)
);

XOR2x1_ASAP7_75t_R c7706(
.A(net7763),
.B(net2163),
.Y(net7774)
);

NOR3x1_ASAP7_75t_R c7707(
.A(net7761),
.B(net7755),
.C(net7748),
.Y(net7775)
);

XOR2x2_ASAP7_75t_R c7708(
.A(net7770),
.B(net9640),
.Y(net7776)
);

NOR3x2_ASAP7_75t_R c7709(
.B(net7751),
.C(net6846),
.A(net7775),
.Y(net7777)
);

NOR3xp33_ASAP7_75t_R c7710(
.A(net6847),
.B(net7753),
.C(net7775),
.Y(net7778)
);

OAI33xp33_ASAP7_75t_R c7711(
.A1(net7749),
.A2(net7745),
.A3(net7778),
.B1(net7767),
.B2(net6832),
.B3(net6869),
.Y(net7779)
);

OA21x2_ASAP7_75t_R c7712(
.A1(net7525),
.A2(net7771),
.B(net10301),
.Y(net7780)
);

OAI21x1_ASAP7_75t_R c7713(
.A1(net7772),
.A2(net7776),
.B(net7775),
.Y(net7781)
);

OAI21xp33_ASAP7_75t_R c7714(
.A1(net7778),
.A2(net7770),
.B(net7780),
.Y(net7782)
);

OAI21xp5_ASAP7_75t_R c7715(
.A1(net7760),
.A2(net6847),
.B(net9640),
.Y(net7783)
);

DFFASRHQNx1_ASAP7_75t_R c7716(
.D(net7709),
.RESETN(net7753),
.SETN(net7742),
.CLK(clk),
.QN(net7784)
);

OR3x1_ASAP7_75t_R c7717(
.A(net7746),
.B(net7784),
.C(net7650),
.Y(net7785)
);

AO222x2_ASAP7_75t_R c7718(
.A1(net7770),
.A2(net7775),
.B1(net7752),
.B2(net7784),
.C1(net6869),
.C2(out13),
.Y(net7786)
);

INVx2_ASAP7_75t_R c7719(
.A(net4963),
.Y(net7787)
);

XOR2xp5_ASAP7_75t_R c7720(
.A(net7601),
.B(net6764),
.Y(net7788)
);

AND2x2_ASAP7_75t_R c7721(
.A(net5960),
.B(net9789),
.Y(net7789)
);

AND2x4_ASAP7_75t_R c7722(
.A(net6909),
.B(net6749),
.Y(net7790)
);

INVx3_ASAP7_75t_R c7723(
.A(net5957),
.Y(net7791)
);

INVx4_ASAP7_75t_R c7724(
.A(net9152),
.Y(net7792)
);

AND2x6_ASAP7_75t_R c7725(
.A(net5689),
.B(net5960),
.Y(net7793)
);

HAxp5_ASAP7_75t_R c7726(
.A(net7582),
.B(net5926),
.CON(net7794)
);

AOI22xp5_ASAP7_75t_R c7727(
.A1(net6764),
.A2(net5584),
.B1(net6899),
.B2(net7759),
.Y(net7795)
);

INVx5_ASAP7_75t_R c7728(
.A(net10417),
.Y(net7796)
);

NAND2x1_ASAP7_75t_R c7729(
.A(net6899),
.B(net6749),
.Y(net7797)
);

INVx6_ASAP7_75t_R c7730(
.A(net7777),
.Y(net7798)
);

ICGx2_ASAP7_75t_R c7731(
.ENA(net6954),
.SE(net5991),
.CLK(clk),
.GCLK(net7799)
);

AO33x2_ASAP7_75t_R c7732(
.A1(net7687),
.A2(net7477),
.A3(net6925),
.B1(net7469),
.B2(net7586),
.B3(net10281),
.Y(net7800)
);

INVx8_ASAP7_75t_R c7733(
.A(net7593),
.Y(net7801)
);

NAND2x1p5_ASAP7_75t_R c7734(
.A(net7735),
.B(net6925),
.Y(net7802)
);

OR3x2_ASAP7_75t_R c7735(
.A(net6945),
.B(net6869),
.C(net10110),
.Y(net7803)
);

NAND2x2_ASAP7_75t_R c7736(
.A(net7796),
.B(net7793),
.Y(net7804)
);

INVxp33_ASAP7_75t_R c7737(
.A(net10372),
.Y(net7805)
);

INVxp67_ASAP7_75t_R c7738(
.A(net6900),
.Y(net7806)
);

NAND2xp33_ASAP7_75t_R c7739(
.A(net5991),
.B(net6749),
.Y(net7807)
);

BUFx10_ASAP7_75t_R c7740(
.A(net10365),
.Y(net7808)
);

NAND2xp5_ASAP7_75t_R c7741(
.A(net7567),
.B(net6895),
.Y(net7809)
);

NAND2xp67_ASAP7_75t_R c7742(
.A(net7573),
.B(net7658),
.Y(net7810)
);

NOR2x1_ASAP7_75t_R c7743(
.A(net5960),
.B(net5609),
.Y(net7811)
);

NOR2x1p5_ASAP7_75t_R c7744(
.A(net7668),
.B(net5836),
.Y(net7812)
);

NOR2x2_ASAP7_75t_R c7745(
.A(net6952),
.B(net7619),
.Y(net7813)
);

NOR2xp33_ASAP7_75t_R c7746(
.A(net7808),
.B(net6764),
.Y(net7814)
);

BUFx12_ASAP7_75t_R c7747(
.A(net10491),
.Y(net7815)
);

BUFx12f_ASAP7_75t_R c7748(
.A(net10380),
.Y(net7816)
);

NOR2xp67_ASAP7_75t_R c7749(
.A(net7790),
.B(net7619),
.Y(net7817)
);

SDFHx1_ASAP7_75t_R c7750(
.D(net7803),
.SE(net6952),
.SI(net7814),
.CLK(clk),
.QN(net7818)
);

AOI31xp33_ASAP7_75t_R c7751(
.A1(net7813),
.A2(net7564),
.A3(net10281),
.B(net10299),
.Y(net7819)
);

BUFx16f_ASAP7_75t_R c7752(
.A(net10146),
.Y(net7820)
);

BUFx24_ASAP7_75t_R c7753(
.A(net10365),
.Y(net7821)
);

ICGx2p67DC_ASAP7_75t_R c7754(
.ENA(net7804),
.SE(net7712),
.CLK(clk),
.GCLK(net7822)
);

OR2x2_ASAP7_75t_R c7755(
.A(net1336),
.B(net7806),
.Y(net7823)
);

OR2x4_ASAP7_75t_R c7756(
.A(net7812),
.B(net7791),
.Y(net7824)
);

BUFx2_ASAP7_75t_R c7757(
.A(net10119),
.Y(net7825)
);

BUFx3_ASAP7_75t_R c7758(
.A(net6832),
.Y(net7826)
);

BUFx4_ASAP7_75t_R c7759(
.A(net10119),
.Y(net7827)
);

BUFx4f_ASAP7_75t_R c7760(
.A(net7728),
.Y(net7828)
);

OR2x6_ASAP7_75t_R c7761(
.A(net7818),
.B(net7826),
.Y(net7829)
);

XNOR2x1_ASAP7_75t_R c7762(
.B(net5599),
.A(net7806),
.Y(net7830)
);

XNOR2x2_ASAP7_75t_R c7763(
.A(net6749),
.B(net7601),
.Y(net7831)
);

XNOR2xp5_ASAP7_75t_R c7764(
.A(net6615),
.B(net10302),
.Y(net7832)
);

XOR2x1_ASAP7_75t_R c7765(
.A(net7798),
.B(net7822),
.Y(net7833)
);

BUFx5_ASAP7_75t_R c7766(
.A(net6937),
.Y(net7834)
);

XOR2x2_ASAP7_75t_R c7767(
.A(out13),
.B(net10281),
.Y(net7835)
);

AOI31xp67_ASAP7_75t_R c7768(
.A1(net6924),
.A2(net7793),
.A3(net7826),
.B(net7831),
.Y(net7836)
);

XOR2xp5_ASAP7_75t_R c7769(
.A(net6787),
.B(net7708),
.Y(net7837)
);

AND2x2_ASAP7_75t_R c7770(
.A(net7834),
.B(net10110),
.Y(net7838)
);

AND2x4_ASAP7_75t_R c7771(
.A(net7829),
.B(net6869),
.Y(net7839)
);

BUFx6f_ASAP7_75t_R c7772(
.A(net10450),
.Y(net7840)
);

AOI221xp5_ASAP7_75t_R c7773(
.A1(net6943),
.A2(net7791),
.B1(net7812),
.B2(net6906),
.C(net7826),
.Y(net7841)
);

AND2x6_ASAP7_75t_R c7774(
.A(net7840),
.B(net7818),
.Y(net7842)
);

OR3x4_ASAP7_75t_R c7775(
.A(net7686),
.B(net7842),
.C(net10302),
.Y(net7843)
);

AND3x1_ASAP7_75t_R c7776(
.A(net7793),
.B(net7840),
.C(net7754),
.Y(net7844)
);

NAND4xp25_ASAP7_75t_R c7777(
.A(net7836),
.B(net7831),
.C(net7841),
.D(net6804),
.Y(net7845)
);

BUFx8_ASAP7_75t_R c7778(
.A(net10354),
.Y(net7846)
);

CKINVDCx10_ASAP7_75t_R c7779(
.A(net10036),
.Y(net7847)
);

HAxp5_ASAP7_75t_R c7780(
.A(net7823),
.B(net5779),
.CON(net7849),
.SN(net7848)
);

AND3x2_ASAP7_75t_R c7781(
.A(net7827),
.B(net7834),
.C(net6764),
.Y(net7850)
);

NAND2x1_ASAP7_75t_R c7782(
.A(net7708),
.B(net10301),
.Y(net7851)
);

AND3x4_ASAP7_75t_R c7783(
.A(net6846),
.B(net7810),
.C(net7735),
.Y(net7852)
);

SDFHx2_ASAP7_75t_R c7784(
.D(net7816),
.SE(net7849),
.SI(net7836),
.CLK(clk),
.QN(net7853)
);

NAND2x1p5_ASAP7_75t_R c7785(
.A(net7838),
.B(net7852),
.Y(net7854)
);

CKINVDCx11_ASAP7_75t_R c7786(
.A(net10455),
.Y(net7855)
);

NAND2x2_ASAP7_75t_R c7787(
.A(net7812),
.B(net9689),
.Y(net7856)
);

AO21x1_ASAP7_75t_R c7788(
.A1(net7788),
.A2(net7846),
.B(net7853),
.Y(net7857)
);

CKINVDCx12_ASAP7_75t_R c7789(
.A(net9152),
.Y(net7858)
);

NAND2xp33_ASAP7_75t_R c7790(
.A(net7835),
.B(net6764),
.Y(net7859)
);

NAND4xp75_ASAP7_75t_R c7791(
.A(net7856),
.B(net7834),
.C(net7823),
.D(net6906),
.Y(net7860)
);

AO21x2_ASAP7_75t_R c7792(
.A1(net7847),
.A2(net7854),
.B(net7856),
.Y(net7861)
);

AOI21x1_ASAP7_75t_R c7793(
.A1(net7832),
.A2(net7846),
.B(net7850),
.Y(net7862)
);

NAND2xp5_ASAP7_75t_R c7794(
.A(net7862),
.B(net9939),
.Y(net7863)
);

NOR4xp25_ASAP7_75t_R c7795(
.A(net7859),
.B(net7851),
.C(net7862),
.D(out13),
.Y(net7864)
);

AOI21xp33_ASAP7_75t_R c7796(
.A1(net7821),
.A2(net7823),
.B(net10144),
.Y(net7865)
);

AOI21xp5_ASAP7_75t_R c7797(
.A1(net7861),
.A2(net7858),
.B(net10144),
.Y(net7866)
);

AOI222xp33_ASAP7_75t_R c7798(
.A1(net7824),
.A2(net7865),
.B1(net7862),
.B2(net7841),
.C1(net6832),
.C2(net7822),
.Y(net7867)
);

SDFHx3_ASAP7_75t_R c7799(
.D(net7805),
.SE(net7769),
.SI(net7867),
.CLK(clk),
.QN(net7868)
);

AOI311xp33_ASAP7_75t_R c7800(
.A1(net7791),
.A2(net7861),
.A3(net7868),
.B(net7862),
.C(net9689),
.Y(net7869)
);

NOR4xp75_ASAP7_75t_R c7801(
.A(net7855),
.B(net7865),
.C(net7861),
.D(net7868),
.Y(net7870)
);

NAND2xp67_ASAP7_75t_R c7802(
.A(net6964),
.B(net6928),
.Y(net7871)
);

NOR2x1_ASAP7_75t_R c7803(
.A(net6075),
.B(net6701),
.Y(net7872)
);

CKINVDCx14_ASAP7_75t_R c7804(
.A(net10337),
.Y(net7873)
);

NOR2x1p5_ASAP7_75t_R c7805(
.A(net6928),
.B(net7831),
.Y(net7874)
);

NOR2x2_ASAP7_75t_R c7806(
.A(net531),
.B(net7814),
.Y(net7875)
);

FAx1_ASAP7_75t_R c7807(
.A(net7850),
.B(net7841),
.CI(net6979),
.SN(net7877),
.CON(net7876)
);

MAJIxp5_ASAP7_75t_R c7808(
.A(net7810),
.B(net6914),
.C(net10299),
.Y(net7878)
);

NOR2xp33_ASAP7_75t_R c7809(
.A(net6114),
.B(net10059),
.Y(net7879)
);

CKINVDCx16_ASAP7_75t_R c7810(
.A(net10566),
.Y(net7880)
);

CKINVDCx20_ASAP7_75t_R c7811(
.A(net10537),
.Y(net7881)
);

NOR2xp67_ASAP7_75t_R c7812(
.A(net7881),
.B(net6917),
.Y(net7882)
);

OR2x2_ASAP7_75t_R c7813(
.A(net6945),
.B(net6751),
.Y(net7883)
);

MAJx2_ASAP7_75t_R c7814(
.A(net7638),
.B(net7019),
.C(net6114),
.Y(net7884)
);

OR2x4_ASAP7_75t_R c7815(
.A(net7841),
.B(net7586),
.Y(net7885)
);

MAJx3_ASAP7_75t_R c7816(
.A(net7771),
.B(net6979),
.C(net4962),
.Y(net7886)
);

OR2x6_ASAP7_75t_R c7817(
.A(net7008),
.B(net6958),
.Y(net7887)
);

NAND3x1_ASAP7_75t_R c7818(
.A(net7837),
.B(net7882),
.C(net6945),
.Y(net7888)
);

XNOR2x1_ASAP7_75t_R c7819(
.B(net7030),
.A(net7019),
.Y(net7889)
);

CKINVDCx5p33_ASAP7_75t_R c7820(
.A(net10477),
.Y(net7890)
);

CKINVDCx6p67_ASAP7_75t_R c7821(
.A(net10129),
.Y(net7891)
);

XNOR2x2_ASAP7_75t_R c7822(
.A(net7831),
.B(net9859),
.Y(net7892)
);

XNOR2xp5_ASAP7_75t_R c7823(
.A(net7023),
.B(net5152),
.Y(net7893)
);

NAND3x2_ASAP7_75t_R c7824(
.B(net5836),
.C(net7882),
.A(net7574),
.Y(net7894)
);

ICGx3_ASAP7_75t_R c7825(
.ENA(net7878),
.SE(net7877),
.CLK(clk),
.GCLK(net7895)
);

NAND3xp33_ASAP7_75t_R c7826(
.A(net7710),
.B(net6988),
.C(net7875),
.Y(net7896)
);

XOR2x1_ASAP7_75t_R c7827(
.A(net6050),
.B(net7886),
.Y(net7897)
);

XOR2x2_ASAP7_75t_R c7828(
.A(net7843),
.B(net6988),
.Y(net7898)
);

CKINVDCx8_ASAP7_75t_R c7829(
.A(net10118),
.Y(net7899)
);

CKINVDCx9p33_ASAP7_75t_R c7830(
.A(net10377),
.Y(net7900)
);

XOR2xp5_ASAP7_75t_R c7831(
.A(net7891),
.B(net7890),
.Y(net7901)
);

HB1xp67_ASAP7_75t_R c7832(
.A(net10356),
.Y(net7902)
);

NOR3x1_ASAP7_75t_R c7833(
.A(net7732),
.B(net7902),
.C(net7899),
.Y(net7903)
);

AND2x2_ASAP7_75t_R c7834(
.A(net5152),
.B(net7863),
.Y(net7904)
);

NOR3x2_ASAP7_75t_R c7835(
.B(net6994),
.C(net6928),
.A(net10143),
.Y(net7905)
);

AND2x4_ASAP7_75t_R c7836(
.A(net7564),
.B(net7892),
.Y(net7906)
);

HB2xp67_ASAP7_75t_R c7837(
.A(net10085),
.Y(net7907)
);

AND2x6_ASAP7_75t_R c7838(
.A(net7807),
.B(net7898),
.Y(net7908)
);

HAxp5_ASAP7_75t_R c7839(
.A(net6997),
.B(net7638),
.CON(net7909)
);

NAND2x1_ASAP7_75t_R c7840(
.A(net6914),
.B(net7901),
.Y(net7910)
);

NOR3xp33_ASAP7_75t_R c7841(
.A(net7712),
.B(net7875),
.C(net10011),
.Y(net7911)
);

OA21x2_ASAP7_75t_R c7842(
.A1(net7787),
.A2(net6751),
.B(net7771),
.Y(net7912)
);

OAI21x1_ASAP7_75t_R c7843(
.A1(net7909),
.A2(net6972),
.B(net7875),
.Y(net7913)
);

NAND2x1p5_ASAP7_75t_R c7844(
.A(net7800),
.B(net6025),
.Y(net7914)
);

NAND2x2_ASAP7_75t_R c7845(
.A(net7034),
.B(net4834),
.Y(net7915)
);

OAI21xp33_ASAP7_75t_R c7846(
.A1(net6101),
.A2(net6914),
.B(net3272),
.Y(net7916)
);

AOI32xp33_ASAP7_75t_R c7847(
.A1(net7809),
.A2(net7877),
.A3(net7822),
.B1(net6099),
.B2(net6508),
.Y(net7917)
);

NAND2xp33_ASAP7_75t_R c7848(
.A(net6114),
.B(net7884),
.Y(net7918)
);

ICGx4DC_ASAP7_75t_R c7849(
.ENA(net7914),
.SE(net7918),
.CLK(clk),
.GCLK(net7919)
);

AOI321xp33_ASAP7_75t_R c7850(
.A1(net7900),
.A2(net7889),
.A3(net6988),
.B1(net7841),
.B2(net7831),
.C(net7026),
.Y(net7920)
);

OAI21xp5_ASAP7_75t_R c7851(
.A1(net7916),
.A2(net5152),
.B(net6930),
.Y(net7921)
);

OR3x1_ASAP7_75t_R c7852(
.A(net5910),
.B(net7667),
.C(net7895),
.Y(net7922)
);

NAND2xp5_ASAP7_75t_R c7853(
.A(net3316),
.B(net9778),
.Y(net7923)
);

NAND2xp67_ASAP7_75t_R c7854(
.A(net7814),
.B(net7769),
.Y(net7924)
);

OR3x2_ASAP7_75t_R c7855(
.A(net5176),
.B(net7884),
.C(net6837),
.Y(net7925)
);

OR3x4_ASAP7_75t_R c7856(
.A(net7919),
.B(net7922),
.C(net10167),
.Y(net7926)
);

NOR2x1_ASAP7_75t_R c7857(
.A(net7849),
.B(net10018),
.Y(net7927)
);

NOR2x1p5_ASAP7_75t_R c7858(
.A(net7828),
.B(net10304),
.Y(net7928)
);

HB3xp67_ASAP7_75t_R c7859(
.A(net10384),
.Y(net7929)
);

NOR2x2_ASAP7_75t_R c7860(
.A(net3970),
.B(net7918),
.Y(net7930)
);

AOI33xp33_ASAP7_75t_R c7861(
.A1(net7895),
.A2(net7927),
.A3(net7898),
.B1(net7875),
.B2(net7841),
.B3(net7759),
.Y(net7931)
);

NOR2xp33_ASAP7_75t_R c7862(
.A(net7887),
.B(net7899),
.Y(net7932)
);

AND3x1_ASAP7_75t_R c7863(
.A(net7712),
.B(net6751),
.C(net10305),
.Y(net7933)
);

AND3x2_ASAP7_75t_R c7864(
.A(net7908),
.B(net7882),
.C(net7884),
.Y(net7934)
);

HB4xp67_ASAP7_75t_R c7865(
.A(net10448),
.Y(net7935)
);

NOR2xp67_ASAP7_75t_R c7866(
.A(net7932),
.B(net6930),
.Y(net7936)
);

OR2x2_ASAP7_75t_R c7867(
.A(net7928),
.B(net7907),
.Y(net7937)
);

AND3x4_ASAP7_75t_R c7868(
.A(net7911),
.B(net6945),
.C(net5910),
.Y(net7938)
);

SDFHx4_ASAP7_75t_R c7869(
.D(net7933),
.SE(net7012),
.SI(net7921),
.CLK(clk),
.QN(net7939)
);

AO21x1_ASAP7_75t_R c7870(
.A1(net7915),
.A2(net7911),
.B(net6917),
.Y(net7940)
);

AO21x2_ASAP7_75t_R c7871(
.A1(net6958),
.A2(net6945),
.B(net9759),
.Y(net7941)
);

AOI21x1_ASAP7_75t_R c7872(
.A1(net7937),
.A2(net7882),
.B(net7939),
.Y(net7942)
);

SDFLx1_ASAP7_75t_R c7873(
.D(net7930),
.SE(net7936),
.SI(net10304),
.CLK(clk),
.QN(net7943)
);

AOI21xp33_ASAP7_75t_R c7874(
.A1(net6988),
.A2(net7938),
.B(net7942),
.Y(net7944)
);

AOI21xp5_ASAP7_75t_R c7875(
.A1(net7792),
.A2(net7939),
.B(net7937),
.Y(net7945)
);

FAx1_ASAP7_75t_R c7876(
.A(net7686),
.B(net4835),
.CI(net7710),
.SN(net7946)
);

MAJIxp5_ASAP7_75t_R c7877(
.A(net6958),
.B(net7933),
.C(net10304),
.Y(net7947)
);

INVx11_ASAP7_75t_R c7878(
.A(net10337),
.Y(net7948)
);

NAND5xp2_ASAP7_75t_R c7879(
.A(net7944),
.B(net7945),
.C(net7947),
.D(net7921),
.E(net6869),
.Y(net7949)
);

OR2x4_ASAP7_75t_R c7880(
.A(net7948),
.B(net10143),
.Y(net7950)
);

OR2x6_ASAP7_75t_R c7881(
.A(net7938),
.B(net7942),
.Y(net7951)
);

MAJx2_ASAP7_75t_R c7882(
.A(net6643),
.B(net6087),
.C(net7939),
.Y(net7952)
);

MAJx3_ASAP7_75t_R c7883(
.A(net7951),
.B(net7952),
.C(net10143),
.Y(net7953)
);

SDFLx2_ASAP7_75t_R c7884(
.D(net7918),
.SE(net7952),
.SI(net7953),
.CLK(clk),
.QN(net7954)
);

INVx13_ASAP7_75t_R c7885(
.A(net10121),
.Y(net7955)
);

XNOR2x1_ASAP7_75t_R c7886(
.B(net5229),
.A(net6186),
.Y(net7956)
);

INVx1_ASAP7_75t_R c7887(
.A(net6869),
.Y(net7957)
);

INVx2_ASAP7_75t_R c7888(
.A(net10551),
.Y(net7958)
);

XNOR2x2_ASAP7_75t_R c7889(
.A(net4835),
.B(net10059),
.Y(net7959)
);

XNOR2xp5_ASAP7_75t_R c7890(
.A(net7902),
.B(net7853),
.Y(net7960)
);

INVx3_ASAP7_75t_R c7891(
.A(net9280),
.Y(net7961)
);

XOR2x1_ASAP7_75t_R c7892(
.A(net5193),
.B(net7929),
.Y(net7962)
);

INVx4_ASAP7_75t_R c7893(
.A(net9939),
.Y(net7963)
);

INVx5_ASAP7_75t_R c7894(
.A(net10094),
.Y(net7964)
);

INVx6_ASAP7_75t_R c7895(
.A(net6979),
.Y(net7965)
);

INVx8_ASAP7_75t_R c7896(
.A(net10285),
.Y(net7966)
);

INVxp33_ASAP7_75t_R c7897(
.A(net10355),
.Y(net7967)
);

XOR2x2_ASAP7_75t_R c7898(
.A(net6141),
.B(net7960),
.Y(net7968)
);

INVxp67_ASAP7_75t_R c7899(
.A(net10417),
.Y(net7969)
);

BUFx10_ASAP7_75t_R c7900(
.A(net10170),
.Y(net7970)
);

XOR2xp5_ASAP7_75t_R c7901(
.A(net7965),
.B(net7041),
.Y(net7971)
);

AND2x2_ASAP7_75t_R c7902(
.A(net7963),
.B(net5229),
.Y(net7972)
);

BUFx12_ASAP7_75t_R c7903(
.A(net10170),
.Y(net7973)
);

AND2x4_ASAP7_75t_R c7904(
.A(net7853),
.B(net7967),
.Y(net7974)
);

AND2x6_ASAP7_75t_R c7905(
.A(net7961),
.B(net6930),
.Y(net7975)
);

BUFx12f_ASAP7_75t_R c7906(
.A(net10571),
.Y(net7976)
);

HAxp5_ASAP7_75t_R c7907(
.A(net7067),
.B(net7898),
.CON(net7978),
.SN(net7977)
);

O2A1O1Ixp33_ASAP7_75t_R c7908(
.A1(net7955),
.A2(net7956),
.B(net7826),
.C(net7868),
.Y(net7979)
);

NAND2x1_ASAP7_75t_R c7909(
.A(net7883),
.B(net7879),
.Y(net7980)
);

NAND2x1p5_ASAP7_75t_R c7910(
.A(net7967),
.B(net9863),
.Y(net7981)
);

NAND2x2_ASAP7_75t_R c7911(
.A(net7060),
.B(net7966),
.Y(net7982)
);

NAND2xp33_ASAP7_75t_R c7912(
.A(net7950),
.B(net9928),
.Y(net7983)
);

NAND2xp5_ASAP7_75t_R c7913(
.A(net6044),
.B(net6979),
.Y(net7984)
);

NAND2xp67_ASAP7_75t_R c7914(
.A(net7041),
.B(net7075),
.Y(net7985)
);

NOR2x1_ASAP7_75t_R c7915(
.A(net5964),
.B(net6930),
.Y(net7986)
);

NOR2x1p5_ASAP7_75t_R c7916(
.A(net7973),
.B(net5211),
.Y(net7987)
);

BUFx16f_ASAP7_75t_R c7917(
.A(net10494),
.Y(net7988)
);

BUFx24_ASAP7_75t_R c7918(
.A(net10362),
.Y(net7989)
);

NOR2x2_ASAP7_75t_R c7919(
.A(net6837),
.B(net7982),
.Y(net7990)
);

NOR2xp33_ASAP7_75t_R c7920(
.A(net7051),
.B(net10299),
.Y(net7991)
);

NAND3x1_ASAP7_75t_R c7921(
.A(net7976),
.B(net7987),
.C(net7977),
.Y(net7992)
);

NOR2xp67_ASAP7_75t_R c7922(
.A(net7964),
.B(net7967),
.Y(net7993)
);

OR2x2_ASAP7_75t_R c7923(
.A(net6972),
.B(net7941),
.Y(net7994)
);

NAND3x2_ASAP7_75t_R c7924(
.B(net7967),
.C(net7966),
.A(net2475),
.Y(net7995)
);

OR2x4_ASAP7_75t_R c7925(
.A(net7987),
.B(net7586),
.Y(net7996)
);

OR2x6_ASAP7_75t_R c7926(
.A(net7985),
.B(net9686),
.Y(net7997)
);

XNOR2x1_ASAP7_75t_R c7927(
.B(net7958),
.A(net7986),
.Y(net7998)
);

O2A1O1Ixp5_ASAP7_75t_R c7928(
.A1(net7101),
.A2(net7986),
.B(net6136),
.C(net10285),
.Y(net7999)
);

XNOR2x2_ASAP7_75t_R c7929(
.A(net7053),
.B(net6930),
.Y(net8000)
);

BUFx2_ASAP7_75t_R c7930(
.A(net7992),
.Y(net8001)
);

XNOR2xp5_ASAP7_75t_R c7931(
.A(net7979),
.B(net7998),
.Y(net8002)
);

XOR2x1_ASAP7_75t_R c7932(
.A(net7984),
.B(net7956),
.Y(net8003)
);

XOR2x2_ASAP7_75t_R c7933(
.A(net6751),
.B(net10059),
.Y(net8004)
);

BUFx3_ASAP7_75t_R c7934(
.A(net8004),
.Y(net8005)
);

XOR2xp5_ASAP7_75t_R c7935(
.A(net7481),
.B(out13),
.Y(net8006)
);

BUFx4_ASAP7_75t_R c7936(
.A(net8003),
.Y(net8007)
);

AND2x2_ASAP7_75t_R c7937(
.A(net7586),
.B(net7987),
.Y(net8008)
);

OA211x2_ASAP7_75t_R c7938(
.A1(net7880),
.A2(net7985),
.B(net8008),
.C(net7053),
.Y(net8009)
);

NAND3xp33_ASAP7_75t_R c7939(
.A(net8007),
.B(net7990),
.C(net10272),
.Y(net8010)
);

AND2x4_ASAP7_75t_R c7940(
.A(net8000),
.B(net6930),
.Y(net8011)
);

BUFx4f_ASAP7_75t_R c7941(
.A(net10381),
.Y(net8012)
);

AND2x6_ASAP7_75t_R c7942(
.A(net7894),
.B(net7858),
.Y(net8013)
);

SDFLx3_ASAP7_75t_R c7943(
.D(net7980),
.SE(net7994),
.SI(net7922),
.CLK(clk),
.QN(net8014)
);

HAxp5_ASAP7_75t_R c7944(
.A(net5211),
.B(net8013),
.CON(net8015)
);

NAND2x1_ASAP7_75t_R c7945(
.A(net7970),
.B(net7996),
.Y(net8016)
);

NOR3x1_ASAP7_75t_R c7946(
.A(net5076),
.B(net7998),
.C(net7994),
.Y(net8017)
);

NAND2x1p5_ASAP7_75t_R c7947(
.A(net6069),
.B(net7083),
.Y(net8018)
);

NAND2x2_ASAP7_75t_R c7948(
.A(net7966),
.B(net8007),
.Y(net8019)
);

NOR3x2_ASAP7_75t_R c7949(
.B(net8008),
.C(net7990),
.A(net7983),
.Y(net8020)
);

NAND2xp33_ASAP7_75t_R c7950(
.A(net7991),
.B(net7833),
.Y(net8021)
);

NAND2xp5_ASAP7_75t_R c7951(
.A(net7996),
.B(net7053),
.Y(net8022)
);

OA22x2_ASAP7_75t_R c7952(
.A1(net8007),
.A2(net8019),
.B1(net8011),
.B2(net7060),
.Y(net8023)
);

NOR3xp33_ASAP7_75t_R c7953(
.A(net7993),
.B(net8006),
.C(net7969),
.Y(net8024)
);

OA21x2_ASAP7_75t_R c7954(
.A1(net8020),
.A2(net8024),
.B(net10306),
.Y(net8025)
);

BUFx5_ASAP7_75t_R c7955(
.A(net10142),
.Y(net8026)
);

OAI21x1_ASAP7_75t_R c7956(
.A1(net7988),
.A2(net8020),
.B(net10306),
.Y(net8027)
);

OA31x2_ASAP7_75t_R c7957(
.A1(net7912),
.A2(net8021),
.A3(net8025),
.B1(net7054),
.Y(net8028)
);

OAI21xp33_ASAP7_75t_R c7958(
.A1(net7074),
.A2(net8006),
.B(net10306),
.Y(net8029)
);

SDFLx4_ASAP7_75t_R c7959(
.D(net8001),
.SE(net6080),
.SI(net8024),
.CLK(clk),
.QN(net8030)
);

DFFASRHQNx1_ASAP7_75t_R c7960(
.D(net2475),
.RESETN(net8030),
.SETN(net7759),
.CLK(clk),
.QN(net8031)
);

OAI21xp5_ASAP7_75t_R c7961(
.A1(net8015),
.A2(net8031),
.B(net8030),
.Y(net8032)
);

OR3x1_ASAP7_75t_R c7962(
.A(net6973),
.B(net8026),
.C(net8031),
.Y(net8033)
);

OA222x2_ASAP7_75t_R c7963(
.A1(net8005),
.A2(net7892),
.B1(net5260),
.B2(net9959),
.C1(net10272),
.C2(net10306),
.Y(net8034)
);

NOR5xp2_ASAP7_75t_R c7964(
.A(net7960),
.B(net8027),
.C(net8019),
.D(net6972),
.E(net10307),
.Y(net8035)
);

OAI211xp5_ASAP7_75t_R c7965(
.A1(net7997),
.A2(net7991),
.B(net8030),
.C(net10307),
.Y(net8036)
);

OAI22x1_ASAP7_75t_R c7966(
.A1(net8025),
.A2(net7989),
.B1(net9759),
.B2(net10307),
.Y(net8037)
);

OR3x2_ASAP7_75t_R c7967(
.A(net8024),
.B(net9894),
.C(net10048),
.Y(net8038)
);

BUFx6f_ASAP7_75t_R c7968(
.A(net10114),
.Y(net8039)
);

OAI22xp33_ASAP7_75t_R c7969(
.A1(net6198),
.A2(net7892),
.B1(net7190),
.B2(net7161),
.Y(net8040)
);

OR3x4_ASAP7_75t_R c7970(
.A(net5996),
.B(net7138),
.C(net7956),
.Y(net8041)
);

BUFx8_ASAP7_75t_R c7971(
.A(net10141),
.Y(net8042)
);

NAND2xp67_ASAP7_75t_R c7972(
.A(net7898),
.B(net6085),
.Y(net8043)
);

NOR2x1_ASAP7_75t_R c7973(
.A(net7205),
.B(net7165),
.Y(net8044)
);

NOR2x1p5_ASAP7_75t_R c7974(
.A(net7910),
.B(net8043),
.Y(net8045)
);

NOR2x2_ASAP7_75t_R c7975(
.A(net7190),
.B(net10307),
.Y(net8046)
);

AND3x1_ASAP7_75t_R c7976(
.A(net8022),
.B(net8045),
.C(net7051),
.Y(net8047)
);

NOR2xp33_ASAP7_75t_R c7977(
.A(net8042),
.B(net7971),
.Y(net8048)
);

AND3x2_ASAP7_75t_R c7978(
.A(net5325),
.B(net6213),
.C(net7064),
.Y(net8049)
);

NOR2xp67_ASAP7_75t_R c7979(
.A(net7075),
.B(net7954),
.Y(net8050)
);

OR2x2_ASAP7_75t_R c7980(
.A(net7989),
.B(net8013),
.Y(net8051)
);

AND3x4_ASAP7_75t_R c7981(
.A(net7983),
.B(net7950),
.C(net7198),
.Y(net8052)
);

AO21x1_ASAP7_75t_R c7982(
.A1(net7200),
.A2(net8045),
.B(net7026),
.Y(net8053)
);

CKINVDCx10_ASAP7_75t_R c7983(
.A(net10397),
.Y(net8054)
);

CKINVDCx11_ASAP7_75t_R c7984(
.A(net10403),
.Y(net8055)
);

SDFHx1_ASAP7_75t_R c7985(
.D(net7191),
.SE(net8044),
.SI(net8043),
.CLK(clk),
.QN(net8056)
);

OR2x4_ASAP7_75t_R c7986(
.A(net7134),
.B(net8045),
.Y(net8057)
);

OR2x6_ASAP7_75t_R c7987(
.A(net8053),
.B(net9671),
.Y(net8058)
);

AO21x2_ASAP7_75t_R c7988(
.A1(net8050),
.A2(net8014),
.B(net7163),
.Y(net8059)
);

AOI21x1_ASAP7_75t_R c7989(
.A1(net1653),
.A2(net8057),
.B(net10304),
.Y(net8060)
);

AOI21xp33_ASAP7_75t_R c7990(
.A1(net8038),
.A2(net5332),
.B(net10305),
.Y(net8061)
);

CKINVDCx12_ASAP7_75t_R c7991(
.A(net9280),
.Y(net8062)
);

CKINVDCx14_ASAP7_75t_R c7992(
.A(net10355),
.Y(net8063)
);

XNOR2x1_ASAP7_75t_R c7993(
.B(net7981),
.A(net8043),
.Y(net8064)
);

AOI21xp5_ASAP7_75t_R c7994(
.A1(net6085),
.A2(net8047),
.B(net8056),
.Y(net8065)
);

CKINVDCx16_ASAP7_75t_R c7995(
.A(net10396),
.Y(net8066)
);

SDFHx2_ASAP7_75t_R c7996(
.D(net7172),
.SE(net8065),
.SI(net8058),
.CLK(clk),
.QN(net8067)
);

XNOR2x2_ASAP7_75t_R c7997(
.A(net6209),
.B(net7868),
.Y(net8068)
);

XNOR2xp5_ASAP7_75t_R c7998(
.A(net7064),
.B(net8064),
.Y(net8069)
);

SDFHx3_ASAP7_75t_R c7999(
.D(net8062),
.SE(net8059),
.SI(net8064),
.CLK(clk),
.QN(net8070)
);

CKINVDCx20_ASAP7_75t_R c8000(
.A(net10350),
.Y(net8071)
);

FAx1_ASAP7_75t_R c8001(
.A(net8068),
.B(net7122),
.CI(net10287),
.SN(net8072)
);

XOR2x1_ASAP7_75t_R c8002(
.A(net6058),
.B(net8055),
.Y(net8073)
);

XOR2x2_ASAP7_75t_R c8003(
.A(net7119),
.B(net8054),
.Y(net8074)
);

MAJIxp5_ASAP7_75t_R c8004(
.A(net8066),
.B(net6085),
.C(net7148),
.Y(net8075)
);

MAJx2_ASAP7_75t_R c8005(
.A(net7126),
.B(net6256),
.C(net7956),
.Y(net8076)
);

XOR2xp5_ASAP7_75t_R c8006(
.A(net6751),
.B(net7138),
.Y(net8077)
);

SDFHx4_ASAP7_75t_R c8007(
.D(net7122),
.SE(net8068),
.SI(net8019),
.CLK(clk),
.QN(net8078)
);

MAJx3_ASAP7_75t_R c8008(
.A(net4166),
.B(net8055),
.C(net7026),
.Y(net8079)
);

AND2x2_ASAP7_75t_R c8009(
.A(net8049),
.B(net10286),
.Y(net8080)
);

NAND3x1_ASAP7_75t_R c8010(
.A(net8075),
.B(net7956),
.C(net8076),
.Y(net8081)
);

OAI22xp5_ASAP7_75t_R c8011(
.A1(net8071),
.A2(net4369),
.B1(net8070),
.B2(net10304),
.Y(net8082)
);

CKINVDCx5p33_ASAP7_75t_R c8012(
.A(net10159),
.Y(net8083)
);

AND2x4_ASAP7_75t_R c8013(
.A(net8077),
.B(net8078),
.Y(net8084)
);

AND2x6_ASAP7_75t_R c8014(
.A(net8084),
.B(net7983),
.Y(net8085)
);

NAND3x2_ASAP7_75t_R c8015(
.B(net8073),
.C(net8064),
.A(net8076),
.Y(net8086)
);

OAI31xp33_ASAP7_75t_R c8016(
.A1(net8038),
.A2(net8085),
.A3(net8076),
.B(net8054),
.Y(net8087)
);

NAND3xp33_ASAP7_75t_R c8017(
.A(net4369),
.B(net8067),
.C(net2578),
.Y(net8088)
);

OA221x2_ASAP7_75t_R c8018(
.A1(net7969),
.A2(net7481),
.B1(net8086),
.B2(net8064),
.C(net7921),
.Y(net8089)
);

NOR3x1_ASAP7_75t_R c8019(
.A(net7919),
.B(net8088),
.C(net8078),
.Y(net8090)
);

OAI31xp67_ASAP7_75t_R c8020(
.A1(net8056),
.A2(net6085),
.A3(net5260),
.B(net9686),
.Y(net8091)
);

NOR3x2_ASAP7_75t_R c8021(
.B(net7924),
.C(net8083),
.A(net8086),
.Y(net8092)
);

NOR3xp33_ASAP7_75t_R c8022(
.A(net7833),
.B(net7058),
.C(net10309),
.Y(net8093)
);

SDFLx1_ASAP7_75t_R c8023(
.D(net8019),
.SE(net8085),
.SI(net7190),
.CLK(clk),
.QN(net8094)
);

OAI221xp5_ASAP7_75t_R c8024(
.A1(net8081),
.A2(net8019),
.B1(net8031),
.B2(net10021),
.C(net10288),
.Y(net8095)
);

OA21x2_ASAP7_75t_R c8025(
.A1(net6206),
.A2(net7051),
.B(net10004),
.Y(net8096)
);

SDFLx2_ASAP7_75t_R c8026(
.D(net8074),
.SE(net8088),
.SI(net7393),
.CLK(clk),
.QN(net8097)
);

OAI21x1_ASAP7_75t_R c8027(
.A1(net7052),
.A2(net6206),
.B(net8094),
.Y(net8098)
);

OAI21xp33_ASAP7_75t_R c8028(
.A1(net8097),
.A2(net8064),
.B(net8082),
.Y(net8099)
);

OAI311xp33_ASAP7_75t_R c8029(
.A1(net5330),
.A2(net7921),
.A3(net7574),
.B1(net7899),
.C1(net10309),
.Y(net8100)
);

OAI21xp5_ASAP7_75t_R c8030(
.A1(net7051),
.A2(net8094),
.B(net10055),
.Y(net8101)
);

HAxp5_ASAP7_75t_R c8031(
.A(net8083),
.B(net7910),
.CON(net8102)
);

OR3x1_ASAP7_75t_R c8032(
.A(net8094),
.B(net4363),
.C(net9761),
.Y(net8103)
);

OR3x2_ASAP7_75t_R c8033(
.A(net6256),
.B(net8058),
.C(net5105),
.Y(net8104)
);

OR3x4_ASAP7_75t_R c8034(
.A(net8101),
.B(net7921),
.C(net8099),
.Y(net8105)
);

SDFLx3_ASAP7_75t_R c8035(
.D(net7978),
.SE(net7181),
.SI(net7759),
.CLK(clk),
.QN(net8106)
);

AND3x1_ASAP7_75t_R c8036(
.A(net8092),
.B(net8051),
.C(net8064),
.Y(net8107)
);

OR4x1_ASAP7_75t_R c8037(
.A(net8067),
.B(net8079),
.C(net3432),
.D(net10309),
.Y(net8108)
);

CKINVDCx6p67_ASAP7_75t_R c8038(
.A(net10141),
.Y(net8109)
);

AND3x2_ASAP7_75t_R c8039(
.A(net8070),
.B(net7954),
.C(net9662),
.Y(net8110)
);

NAND2x1_ASAP7_75t_R c8040(
.A(net9972),
.B(net10021),
.Y(net8111)
);

SDFLx4_ASAP7_75t_R c8041(
.D(net8039),
.SE(net8108),
.SI(net8018),
.CLK(clk),
.QN(net8112)
);

NAND2x1p5_ASAP7_75t_R c8042(
.A(net8063),
.B(net9662),
.Y(net8113)
);

AND3x4_ASAP7_75t_R c8043(
.A(net8102),
.B(net8109),
.C(net8110),
.Y(net8114)
);

AO21x1_ASAP7_75t_R c8044(
.A1(net8114),
.A2(net8110),
.B(net8074),
.Y(net8115)
);

AO21x2_ASAP7_75t_R c8045(
.A1(net8111),
.A2(net8054),
.B(net9894),
.Y(net8116)
);

AOI21x1_ASAP7_75t_R c8046(
.A1(net8096),
.A2(net8111),
.B(net10029),
.Y(net8117)
);

AOI21xp33_ASAP7_75t_R c8047(
.A1(net7058),
.A2(net8116),
.B(net8115),
.Y(net8118)
);

AOI21xp5_ASAP7_75t_R c8048(
.A1(net8112),
.A2(net9790),
.B(net10001),
.Y(net8119)
);

DFFASRHQNx1_ASAP7_75t_R c8049(
.D(net7189),
.RESETN(net8113),
.SETN(net8097),
.CLK(clk),
.QN(net8120)
);

OA33x2_ASAP7_75t_R c8050(
.A1(net8112),
.A2(net8119),
.A3(net8120),
.B1(net7899),
.B2(net8056),
.B3(net10309),
.Y(net8121)
);

NAND2x2_ASAP7_75t_R c8051(
.A(net7941),
.B(net8086),
.Y(net8122)
);

NAND2xp33_ASAP7_75t_R c8052(
.A(net8033),
.B(net2617),
.Y(net8123)
);

NAND2xp5_ASAP7_75t_R c8053(
.A(net3443),
.B(out25),
.Y(net8124)
);

FAx1_ASAP7_75t_R c8054(
.A(net803),
.B(net8030),
.CI(net6975),
.SN(net8125)
);

SDFHx1_ASAP7_75t_R c8055(
.D(net7922),
.SE(net7875),
.SI(net5105),
.CLK(clk),
.QN(net8126)
);

NAND2xp67_ASAP7_75t_R c8056(
.A(net5394),
.B(net7226),
.Y(net8127)
);

MAJIxp5_ASAP7_75t_R c8057(
.A(net7892),
.B(net4513),
.C(net6342),
.Y(net8128)
);

SDFHx2_ASAP7_75t_R c8058(
.D(net8057),
.SE(net7269),
.SI(net5197),
.CLK(clk),
.QN(net8129)
);

MAJx2_ASAP7_75t_R c8059(
.A(net7226),
.B(net6335),
.C(net7268),
.Y(net8130)
);

MAJx3_ASAP7_75t_R c8060(
.A(net8130),
.B(net2475),
.C(net10309),
.Y(net8131)
);

OAI32xp33_ASAP7_75t_R c8061(
.A1(net7161),
.A2(net8129),
.A3(net7226),
.B1(net6166),
.B2(net7178),
.Y(net8132)
);

SDFHx3_ASAP7_75t_R c8062(
.D(net7858),
.SE(net6975),
.SI(net8031),
.CLK(clk),
.QN(net8133)
);

NOR2x1_ASAP7_75t_R c8063(
.A(net5168),
.B(net1652),
.Y(net8134)
);

NAND3x1_ASAP7_75t_R c8064(
.A(net7260),
.B(net7161),
.C(net7239),
.Y(net8135)
);

NAND3x2_ASAP7_75t_R c8065(
.B(net3557),
.C(out25),
.A(net3272),
.Y(net8136)
);

NOR2x1p5_ASAP7_75t_R c8066(
.A(net8014),
.B(net8082),
.Y(net8137)
);

NAND3xp33_ASAP7_75t_R c8067(
.A(net8132),
.B(net5411),
.C(net10307),
.Y(net8138)
);

CKINVDCx8_ASAP7_75t_R c8068(
.A(net10114),
.Y(net8139)
);

SDFHx4_ASAP7_75t_R c8069(
.D(net7282),
.SE(net8126),
.SI(net8134),
.CLK(clk),
.QN(net8140)
);

SDFLx1_ASAP7_75t_R c8070(
.D(net7162),
.SE(net7284),
.SI(net7287),
.CLK(clk),
.QN(net8141)
);

NOR3x1_ASAP7_75t_R c8071(
.A(net6342),
.B(net8118),
.C(net7268),
.Y(net8142)
);

OR5x1_ASAP7_75t_R c8072(
.A(net7289),
.B(net8057),
.C(net8103),
.D(net7875),
.E(net8133),
.Y(net8143)
);

SDFLx2_ASAP7_75t_R c8073(
.D(net8054),
.SE(net8051),
.SI(net10286),
.CLK(clk),
.QN(net8144)
);

OR4x2_ASAP7_75t_R c8074(
.A(net6332),
.B(net4307),
.C(net6975),
.D(net8133),
.Y(net8145)
);

NOR3x2_ASAP7_75t_R c8075(
.B(net3564),
.C(net8140),
.A(net8141),
.Y(net8146)
);

NOR3xp33_ASAP7_75t_R c8076(
.A(net8130),
.B(net5168),
.C(net10046),
.Y(net8147)
);

SDFLx3_ASAP7_75t_R c8077(
.D(net5197),
.SE(net5411),
.SI(net3557),
.CLK(clk),
.QN(net8148)
);

OA21x2_ASAP7_75t_R c8078(
.A1(net8012),
.A2(net8057),
.B(net3564),
.Y(net8149)
);

NOR2x2_ASAP7_75t_R c8079(
.A(net7286),
.B(net7826),
.Y(net8150)
);

OAI21x1_ASAP7_75t_R c8080(
.A1(net7057),
.A2(net8129),
.B(net8148),
.Y(net8151)
);

OAI21xp33_ASAP7_75t_R c8081(
.A1(net8024),
.A2(net6830),
.B(net9843),
.Y(net8152)
);

OAI21xp5_ASAP7_75t_R c8082(
.A1(net7239),
.A2(net8134),
.B(net8103),
.Y(net8153)
);

OR3x1_ASAP7_75t_R c8083(
.A(net7268),
.B(net8098),
.C(net8024),
.Y(net8154)
);

OR3x2_ASAP7_75t_R c8084(
.A(net8054),
.B(net8141),
.C(net8144),
.Y(net8155)
);

NOR2xp33_ASAP7_75t_R c8085(
.A(net7257),
.B(net10149),
.Y(net8156)
);

OR3x4_ASAP7_75t_R c8086(
.A(net6213),
.B(net8031),
.C(net6214),
.Y(net8157)
);

AND3x1_ASAP7_75t_R c8087(
.A(net6166),
.B(net8156),
.C(net8141),
.Y(net8158)
);

CKINVDCx9p33_ASAP7_75t_R c8088(
.A(net10342),
.Y(net8159)
);

AND3x2_ASAP7_75t_R c8089(
.A(net8158),
.B(net8156),
.C(net8099),
.Y(net8160)
);

AND3x4_ASAP7_75t_R c8090(
.A(net8123),
.B(net8155),
.C(net10286),
.Y(net8161)
);

HB1xp67_ASAP7_75t_R c8091(
.A(net10353),
.Y(net8162)
);

OAI222xp33_ASAP7_75t_R c8092(
.A1(net5394),
.A2(net7178),
.B1(net8134),
.B2(net8141),
.C1(net9968),
.C2(net10061),
.Y(net8163)
);

AO21x1_ASAP7_75t_R c8093(
.A1(net6367),
.A2(net8140),
.B(net2642),
.Y(net8164)
);

AO21x2_ASAP7_75t_R c8094(
.A1(net7879),
.A2(net8133),
.B(net8123),
.Y(net8165)
);

AOI21x1_ASAP7_75t_R c8095(
.A1(net8123),
.A2(net9757),
.B(net10308),
.Y(net8166)
);

AOI21xp33_ASAP7_75t_R c8096(
.A1(net4357),
.A2(net3564),
.B(net8133),
.Y(net8167)
);

SDFLx4_ASAP7_75t_R c8097(
.D(net8159),
.SE(net7287),
.SI(net9906),
.CLK(clk),
.QN(net8168)
);

AOI21xp5_ASAP7_75t_R c8098(
.A1(net8133),
.A2(net6332),
.B(net8141),
.Y(net8169)
);

FAx1_ASAP7_75t_R c8099(
.A(net4513),
.B(net8137),
.CI(net8155),
.SN(net8170)
);

MAJIxp5_ASAP7_75t_R c8100(
.A(net6323),
.B(net6366),
.C(net9814),
.Y(net8171)
);

MAJx2_ASAP7_75t_R c8101(
.A(net8088),
.B(net8152),
.C(net8167),
.Y(net8172)
);

MAJx3_ASAP7_75t_R c8102(
.A(net7227),
.B(net8162),
.C(net8144),
.Y(net8173)
);

OR5x2_ASAP7_75t_R c8103(
.A(net6335),
.B(net8162),
.C(net8123),
.D(net7269),
.E(net6204),
.Y(net8174)
);

NAND3x1_ASAP7_75t_R c8104(
.A(net6204),
.B(net8168),
.C(net8123),
.Y(net8175)
);

NAND3x2_ASAP7_75t_R c8105(
.B(net6214),
.C(net8150),
.A(net8167),
.Y(net8176)
);

A2O1A1Ixp33_ASAP7_75t_R c8106(
.A1(net8133),
.A2(net8148),
.B(net10030),
.C(net10033),
.Y(net8177)
);

NAND3xp33_ASAP7_75t_R c8107(
.A(net8177),
.B(net8170),
.C(net8167),
.Y(net8178)
);

NOR2xp67_ASAP7_75t_R c8108(
.A(net8171),
.B(net8178),
.Y(net8179)
);

NOR3x1_ASAP7_75t_R c8109(
.A(net7875),
.B(net8141),
.C(net6366),
.Y(net8180)
);

NOR3x2_ASAP7_75t_R c8110(
.B(net8167),
.C(net8155),
.A(net8136),
.Y(net8181)
);

NOR3xp33_ASAP7_75t_R c8111(
.A(net7269),
.B(net8174),
.C(net8180),
.Y(net8182)
);

AND4x1_ASAP7_75t_R c8112(
.A(net6335),
.B(net8133),
.C(net9814),
.D(net10149),
.Y(net8183)
);

OA21x2_ASAP7_75t_R c8113(
.A1(net8099),
.A2(net8182),
.B(net8133),
.Y(net8184)
);

OAI21x1_ASAP7_75t_R c8114(
.A1(net8086),
.A2(net8181),
.B(net8179),
.Y(net8185)
);

OR2x2_ASAP7_75t_R c8115(
.A(net8180),
.B(net9877),
.Y(net8186)
);

OAI21xp33_ASAP7_75t_R c8116(
.A1(net7950),
.A2(net8156),
.B(net8167),
.Y(net8187)
);

OR2x4_ASAP7_75t_R c8117(
.A(net8187),
.B(net8160),
.Y(net8188)
);

OAI21xp5_ASAP7_75t_R c8118(
.A1(net7893),
.A2(net8188),
.B(net8030),
.Y(net8189)
);

OR3x1_ASAP7_75t_R c8119(
.A(net8175),
.B(net8080),
.C(net8168),
.Y(net8190)
);

DFFASRHQNx1_ASAP7_75t_R c8120(
.D(net7083),
.RESETN(net8185),
.SETN(net10309),
.CLK(clk),
.QN(net8191)
);

OR3x2_ASAP7_75t_R c8121(
.A(net8169),
.B(net8106),
.C(net9895),
.Y(net8192)
);

OR3x4_ASAP7_75t_R c8122(
.A(net8179),
.B(net8123),
.C(net9757),
.Y(net8193)
);

AND3x1_ASAP7_75t_R c8123(
.A(net8051),
.B(net8165),
.C(net8164),
.Y(net8194)
);

SDFHx1_ASAP7_75t_R c8124(
.D(net7263),
.SE(net7287),
.SI(net10151),
.CLK(clk),
.QN(net8195)
);

AND3x2_ASAP7_75t_R c8125(
.A(net8173),
.B(net8192),
.C(net8169),
.Y(net8196)
);

AND3x4_ASAP7_75t_R c8126(
.A(net8196),
.B(net6366),
.C(net3557),
.Y(net8197)
);

HB2xp67_ASAP7_75t_R c8127(
.A(net10342),
.Y(net8198)
);

AO21x1_ASAP7_75t_R c8128(
.A1(net7268),
.A2(net9762),
.B(net9843),
.Y(net8199)
);

AO21x2_ASAP7_75t_R c8129(
.A1(net7118),
.A2(net8164),
.B(net8199),
.Y(net8200)
);

AOI21x1_ASAP7_75t_R c8130(
.A1(net8183),
.A2(net7287),
.B(net8190),
.Y(net8201)
);

AOI21xp33_ASAP7_75t_R c8131(
.A1(net8151),
.A2(net8197),
.B(net8167),
.Y(net8202)
);

AOI21xp5_ASAP7_75t_R c8132(
.A1(net8082),
.A2(net8148),
.B(net10058),
.Y(net8203)
);

FAx1_ASAP7_75t_R c8133(
.A(net8202),
.B(net8134),
.CI(net9997),
.SN(net8204)
);

AND4x2_ASAP7_75t_R c8160(
.A(net6419),
.B(net4549),
.C(out3),
.D(net5492),
.Y(net8205)
);

SDFHx2_ASAP7_75t_R c8161(
.D(net8134),
.SE(net7954),
.SI(net8240),
.CLK(clk),
.QN(net8206)
);

AO211x2_ASAP7_75t_R c8162(
.A1(net7362),
.A2(net8195),
.B(net6426),
.C(net8245),
.Y(net8207)
);

MAJIxp5_ASAP7_75t_R c8163(
.A(net7148),
.B(net8206),
.C(net8242),
.Y(net8208)
);

HB3xp67_ASAP7_75t_R c8164(
.A(net10341),
.Y(out6)
);

AO22x1_ASAP7_75t_R c8165(
.A1(net6263),
.A2(net6444),
.B1(net5495),
.B2(net8134),
.Y(net8209)
);

AO22x2_ASAP7_75t_R c8166(
.A1(net7311),
.A2(net7369),
.B1(net8234),
.B2(net10069),
.Y(net8210)
);

AO31x2_ASAP7_75t_R c8167(
.A1(net7340),
.A2(net7232),
.A3(net8242),
.B(net9638),
.Y(net8211)
);

MAJx2_ASAP7_75t_R c8168(
.A(net8206),
.B(net8234),
.C(net10075),
.Y(net8212)
);

MAJx3_ASAP7_75t_R c8169(
.A(net8210),
.B(net8212),
.C(net8161),
.Y(net8213)
);

NAND3x1_ASAP7_75t_R c8170(
.A(net5495),
.B(net7354),
.C(net8234),
.Y(net8214)
);

NAND3x2_ASAP7_75t_R c8171(
.B(net8098),
.C(net8212),
.A(net8245),
.Y(net8215)
);

AOI211x1_ASAP7_75t_R c8172(
.A1(net8241),
.A2(net8239),
.B(net6444),
.C(net8247),
.Y(net8216)
);

NAND3xp33_ASAP7_75t_R c8173(
.A(net8106),
.B(net8195),
.C(net7369),
.Y(net8217)
);

NOR3x1_ASAP7_75t_R c8174(
.A(net5446),
.B(net7184),
.C(net8247),
.Y(net8218)
);

NOR3x2_ASAP7_75t_R c8175(
.B(net5290),
.C(net7184),
.A(net8236),
.Y(out20)
);

A2O1A1O1Ixp25_ASAP7_75t_R c8176(
.A1(net8214),
.A2(net8245),
.B(net8206),
.C(net8234),
.D(net8134),
.Y(net8219)
);

NOR3xp33_ASAP7_75t_R c8177(
.A(net6300),
.B(net8247),
.C(net5511),
.Y(net8220)
);

OA21x2_ASAP7_75t_R c8178(
.A1(net8103),
.A2(net8251),
.B(net8205),
.Y(net8221)
);

OAI21x1_ASAP7_75t_R c8179(
.A1(net8233),
.A2(net10069),
.B(net10310),
.Y(out21)
);

OAI21xp33_ASAP7_75t_R c8180(
.A1(net8248),
.A2(net8249),
.B(net10290),
.Y(net8222)
);

OAI21xp5_ASAP7_75t_R c8181(
.A1(net8234),
.A2(net8208),
.B(net8206),
.Y(net8223)
);

OR3x1_ASAP7_75t_R c8182(
.A(net8205),
.B(net7148),
.C(net10310),
.Y(out11)
);

OR3x2_ASAP7_75t_R c8183(
.A(net2747),
.B(net7350),
.C(net9924),
.Y(net8224)
);

SDFHx3_ASAP7_75t_R c8184(
.D(net8118),
.SE(net8221),
.SI(net10075),
.CLK(clk),
.QN(out17)
);

AND5x1_ASAP7_75t_R c8185(
.A(net8238),
.B(net7328),
.C(net8106),
.D(net6446),
.Y(net8225)
);

OAI321xp33_ASAP7_75t_R c8186(
.A1(net8240),
.A2(net8207),
.A3(net8206),
.B1(out17),
.B2(out25),
.C(net7232),
.Y(net8226)
);

AOI211xp5_ASAP7_75t_R c8187(
.A1(net8217),
.A2(out17),
.B(out1),
.C(out23),
.Y(net8227)
);

AND5x2_ASAP7_75t_R c8188(
.A(net4549),
.B(out17),
.C(net8247),
.D(net9968),
.E(net10005),
.Y(net8228)
);

OAI33xp33_ASAP7_75t_R c8189(
.A1(net6426),
.A2(net8222),
.A3(net8247),
.B1(out17),
.B2(net5411),
.B3(net8191),
.Y(net8229)
);

AO222x2_ASAP7_75t_R c8190(
.A1(net8211),
.A2(net8245),
.B1(net7354),
.B2(net8234),
.C1(out10),
.C2(net10289),
.Y(net8230)
);

OR3x4_ASAP7_75t_R c8191(
.A(net8242),
.B(net5492),
.C(net9638),
.Y(out18)
);

AND3x1_ASAP7_75t_R c8192(
.A(out18),
.B(net10008),
.C(net10121),
.Y(net8231)
);

AND3x2_ASAP7_75t_R c8193(
.A(net6381),
.B(net7365),
.C(net5411),
.Y(net8232)
);

SDFHx4_ASAP7_75t_R c8194(
.D(net7321),
.SE(net7369),
.SI(net5462),
.CLK(clk),
.QN(net8233)
);

AND3x4_ASAP7_75t_R c8195(
.A(net4549),
.B(net7340),
.C(net8115),
.Y(out24)
);

AO21x1_ASAP7_75t_R c8196(
.A1(net7271),
.A2(net7304),
.B(net8233),
.Y(net8234)
);

AO21x2_ASAP7_75t_R c8197(
.A1(net7232),
.A2(net8161),
.B(net5492),
.Y(net8235)
);

SDFLx1_ASAP7_75t_R c8198(
.D(net7293),
.SE(net5411),
.SI(net2747),
.CLK(clk),
.QN(net8236)
);

AOI21x1_ASAP7_75t_R c8199(
.A1(net6378),
.A2(out9),
.B(net6300),
.Y(net8237)
);

AOI21xp33_ASAP7_75t_R c8200(
.A1(net8237),
.A2(net4600),
.B(net8106),
.Y(net8238)
);

AOI22x1_ASAP7_75t_R c8201(
.A1(net7341),
.A2(net8236),
.B1(net8161),
.B2(out9),
.Y(net8239)
);

AOI21xp5_ASAP7_75t_R c8202(
.A1(net8235),
.A2(net8234),
.B(net10290),
.Y(net8240)
);

FAx1_ASAP7_75t_R c8203(
.A(net7265),
.B(net7311),
.CI(net5411),
.SN(net8241)
);

MAJIxp5_ASAP7_75t_R c8204(
.A(net5511),
.B(net6419),
.C(net7232),
.Y(net8242)
);

AOI22xp33_ASAP7_75t_R c8205(
.A1(net6413),
.A2(net6300),
.B1(net8242),
.B2(net9925),
.Y(out22)
);

MAJx2_ASAP7_75t_R c8206(
.A(net2745),
.B(net6446),
.C(net7369),
.Y(net8243)
);

AOI22xp5_ASAP7_75t_R c8207(
.A1(net8124),
.A2(net7350),
.B1(net7354),
.B2(net6300),
.Y(net8244)
);

SDFLx2_ASAP7_75t_R c8208(
.D(net7240),
.SE(net7365),
.SI(net10292),
.CLK(clk),
.QN(net8245)
);

MAJx3_ASAP7_75t_R c8209(
.A(net6383),
.B(net6263),
.C(net8195),
.Y(out14)
);

NAND3x1_ASAP7_75t_R c8210(
.A(net8115),
.B(net8134),
.C(net4549),
.Y(net8246)
);

NAND3x2_ASAP7_75t_R c8211(
.B(net7363),
.C(net8242),
.A(net7311),
.Y(net8247)
);

NAND3xp33_ASAP7_75t_R c8212(
.A(net5492),
.B(net4600),
.C(net9892),
.Y(net8248)
);

SDFLx3_ASAP7_75t_R c8213(
.D(net8244),
.SE(net8245),
.SI(net7184),
.CLK(clk),
.QN(net8249)
);

NOR3x1_ASAP7_75t_R c8214(
.A(net7328),
.B(net8249),
.C(net8247),
.Y(net8250)
);

NOR3x2_ASAP7_75t_R c8215(
.B(net7954),
.C(net7271),
.A(net10043),
.Y(out12)
);

HB4xp67_ASAP7_75t_R c8216(
.A(net10341),
.Y(net8251)
);

INVx11_ASAP7_75t_R c8217(
.A(net7444),
.Y(net8252)
);

INVx13_ASAP7_75t_R c8218(
.A(net9173),
.Y(net8253)
);

OR2x6_ASAP7_75t_R c8219(
.A(net4609),
.B(net7415),
.Y(net8254)
);

INVx1_ASAP7_75t_R c8220(
.A(net8252),
.Y(net8255)
);

INVx2_ASAP7_75t_R c8221(
.A(net7427),
.Y(net8256)
);

INVx3_ASAP7_75t_R c8222(
.A(net8253),
.Y(net8257)
);

INVx4_ASAP7_75t_R c8223(
.A(net6533),
.Y(net8258)
);

INVx5_ASAP7_75t_R c8224(
.A(net7444),
.Y(net8259)
);

XNOR2x1_ASAP7_75t_R c8225(
.B(net5584),
.A(net6510),
.Y(net8260)
);

INVx6_ASAP7_75t_R c8226(
.A(net6480),
.Y(net8261)
);

INVx8_ASAP7_75t_R c8227(
.A(net7423),
.Y(net8262)
);

INVxp33_ASAP7_75t_R c8228(
.A(net8253),
.Y(net8263)
);

NOR3xp33_ASAP7_75t_R c8229(
.A(net8259),
.B(net7382),
.C(net10249),
.Y(net8264)
);

XNOR2x2_ASAP7_75t_R c8230(
.A(net6519),
.B(net7444),
.Y(net8265)
);

INVxp67_ASAP7_75t_R c8231(
.A(net5599),
.Y(net8266)
);

BUFx10_ASAP7_75t_R c8232(
.A(net8266),
.Y(net8267)
);

BUFx12_ASAP7_75t_R c8233(
.A(net8259),
.Y(net8268)
);

BUFx12f_ASAP7_75t_R c8234(
.A(net9173),
.Y(net8269)
);

BUFx16f_ASAP7_75t_R c8235(
.A(net7408),
.Y(net8270)
);

BUFx24_ASAP7_75t_R c8236(
.A(net8259),
.Y(net8271)
);

BUFx2_ASAP7_75t_R c8237(
.A(net8257),
.Y(net8272)
);

BUFx3_ASAP7_75t_R c8238(
.A(net7415),
.Y(net8273)
);

BUFx4_ASAP7_75t_R c8239(
.A(net7452),
.Y(net8274)
);

XNOR2xp5_ASAP7_75t_R c8240(
.A(net8261),
.B(net7399),
.Y(net8275)
);

XOR2x1_ASAP7_75t_R c8241(
.A(net8266),
.B(net8275),
.Y(net8276)
);

BUFx4f_ASAP7_75t_R c8242(
.A(net8276),
.Y(net8277)
);

BUFx5_ASAP7_75t_R c8243(
.A(net8275),
.Y(net8278)
);

BUFx6f_ASAP7_75t_R c8244(
.A(net8256),
.Y(net8279)
);

BUFx8_ASAP7_75t_R c8245(
.A(net7428),
.Y(net8280)
);

ICGx4_ASAP7_75t_R c8246(
.ENA(net5574),
.SE(net8264),
.CLK(clk),
.GCLK(net8281)
);

CKINVDCx10_ASAP7_75t_R c8247(
.A(net5532),
.Y(net8282)
);

CKINVDCx11_ASAP7_75t_R c8248(
.A(net8268),
.Y(net8283)
);

CKINVDCx12_ASAP7_75t_R c8249(
.A(net6528),
.Y(net8284)
);

CKINVDCx14_ASAP7_75t_R c8250(
.A(net8255),
.Y(net8285)
);

CKINVDCx16_ASAP7_75t_R c8251(
.A(net7407),
.Y(net8286)
);

CKINVDCx20_ASAP7_75t_R c8252(
.A(net9217),
.Y(net8287)
);

CKINVDCx5p33_ASAP7_75t_R c8253(
.A(net8281),
.Y(net8288)
);

CKINVDCx6p67_ASAP7_75t_R c8254(
.A(net8278),
.Y(net8289)
);

CKINVDCx8_ASAP7_75t_R c8255(
.A(net8287),
.Y(net8290)
);

XOR2x2_ASAP7_75t_R c8256(
.A(net8286),
.B(net8274),
.Y(net8291)
);

XOR2xp5_ASAP7_75t_R c8257(
.A(net8285),
.B(net8275),
.Y(net8292)
);

AND2x2_ASAP7_75t_R c8258(
.A(net8280),
.B(net8260),
.Y(net8293)
);

AND2x4_ASAP7_75t_R c8259(
.A(net8268),
.B(net8290),
.Y(net8294)
);

AND2x6_ASAP7_75t_R c8260(
.A(net8292),
.B(net8262),
.Y(net8295)
);

CKINVDCx9p33_ASAP7_75t_R c8261(
.A(net8291),
.Y(net8296)
);

HAxp5_ASAP7_75t_R c8262(
.A(net7422),
.B(net8280),
.CON(net8298),
.SN(net8297)
);

HB1xp67_ASAP7_75t_R c8263(
.A(net7445),
.Y(net8299)
);

NAND2x1_ASAP7_75t_R c8264(
.A(net8283),
.B(net7444),
.Y(net8300)
);

HB2xp67_ASAP7_75t_R c8265(
.A(net8290),
.Y(net8301)
);

NAND2x1p5_ASAP7_75t_R c8266(
.A(net8269),
.B(net8297),
.Y(net8302)
);

HB3xp67_ASAP7_75t_R c8267(
.A(net8301),
.Y(net8303)
);

NAND2x2_ASAP7_75t_R c8268(
.A(net8283),
.B(net8263),
.Y(net8304)
);

NAND2xp33_ASAP7_75t_R c8269(
.A(net8304),
.B(net8290),
.Y(net8305)
);

HB4xp67_ASAP7_75t_R c8270(
.A(net8272),
.Y(net8306)
);

NAND2xp5_ASAP7_75t_R c8271(
.A(net8295),
.B(net8291),
.Y(net8307)
);

NAND2xp67_ASAP7_75t_R c8272(
.A(net8277),
.B(net8307),
.Y(net8308)
);

NOR2x1_ASAP7_75t_R c8273(
.A(net6510),
.B(net8296),
.Y(net8309)
);

OA21x2_ASAP7_75t_R c8274(
.A1(net8270),
.A2(net8287),
.B(net8296),
.Y(net8310)
);

NOR2x1p5_ASAP7_75t_R c8275(
.A(net8254),
.B(net8307),
.Y(net8311)
);

NOR2x2_ASAP7_75t_R c8276(
.A(net8274),
.B(net8260),
.Y(net8312)
);

NOR2xp33_ASAP7_75t_R c8277(
.A(net8298),
.B(net8287),
.Y(net8313)
);

NOR2xp67_ASAP7_75t_R c8278(
.A(net8313),
.B(net8302),
.Y(net8314)
);

OR2x2_ASAP7_75t_R c8279(
.A(net8288),
.B(net6510),
.Y(net8315)
);

OR2x4_ASAP7_75t_R c8280(
.A(net8292),
.B(net8301),
.Y(net8316)
);

OR2x6_ASAP7_75t_R c8281(
.A(net8314),
.B(net8315),
.Y(net8317)
);

AOI31xp33_ASAP7_75t_R c8282(
.A1(net8305),
.A2(net8313),
.A3(net8315),
.B(net8279),
.Y(net8318)
);

XNOR2x1_ASAP7_75t_R c8283(
.B(net8265),
.A(net8317),
.Y(net8319)
);

AOI31xp67_ASAP7_75t_R c8284(
.A1(net8319),
.A2(net8317),
.A3(net7445),
.B(net8315),
.Y(net8320)
);

NAND4xp25_ASAP7_75t_R c8285(
.A(net8308),
.B(net7428),
.C(net7397),
.D(net8296),
.Y(net8321)
);

OAI21x1_ASAP7_75t_R c8286(
.A1(net8284),
.A2(net5588),
.B(net10311),
.Y(net8322)
);

OAI21xp33_ASAP7_75t_R c8287(
.A1(net8316),
.A2(net8310),
.B(net8302),
.Y(net8323)
);

SDFLx4_ASAP7_75t_R c8288(
.D(net8281),
.SE(net8317),
.SI(net8318),
.CLK(clk),
.QN(net8324)
);

DFFASRHQNx1_ASAP7_75t_R c8289(
.D(net8309),
.RESETN(net8308),
.SETN(net8317),
.CLK(clk),
.QN(net8325)
);

XNOR2x2_ASAP7_75t_R c8290(
.A(net7423),
.B(net8319),
.Y(net8326)
);

XNOR2xp5_ASAP7_75t_R c8291(
.A(net7408),
.B(net8313),
.Y(net8327)
);

NAND4xp75_ASAP7_75t_R c8292(
.A(net8306),
.B(net8324),
.C(net8311),
.D(net8323),
.Y(net8328)
);

NOR4xp25_ASAP7_75t_R c8293(
.A(net8300),
.B(net8288),
.C(net8254),
.D(net8296),
.Y(net8329)
);

XOR2x1_ASAP7_75t_R c8294(
.A(net8329),
.B(net8327),
.Y(net8330)
);

OAI21xp5_ASAP7_75t_R c8295(
.A1(net8271),
.A2(net8263),
.B(net8323),
.Y(net8331)
);

NOR4xp75_ASAP7_75t_R c8296(
.A(net8331),
.B(net8287),
.C(net8317),
.Y(net8332)
);

SDFHx1_ASAP7_75t_R c8297(
.D(net8310),
.SE(net8309),
.SI(net8331),
.CLK(clk),
.QN(net8333)
);

O2A1O1Ixp33_ASAP7_75t_R c8298(
.A1(net8331),
.A2(net8316),
.B(net8275),
.C(net9659),
.Y(net8334)
);

AO33x2_ASAP7_75t_R c8299(
.A1(net8331),
.A2(net8333),
.A3(net8279),
.B1(net8275),
.B2(net7399),
.B3(net9817),
.Y(net8335)
);

XOR2x2_ASAP7_75t_R c8300(
.A(net7485),
.B(net8299),
.Y(net8336)
);

XOR2xp5_ASAP7_75t_R c8301(
.A(net7404),
.B(net10278),
.Y(net8337)
);

AND2x2_ASAP7_75t_R c8302(
.A(net8323),
.B(net8273),
.Y(net8338)
);

INVx11_ASAP7_75t_R c8303(
.A(net9187),
.Y(net8339)
);

AND2x4_ASAP7_75t_R c8304(
.A(net8326),
.B(net7513),
.Y(net8340)
);

AND2x6_ASAP7_75t_R c8305(
.A(net8302),
.B(net8323),
.Y(net8341)
);

HAxp5_ASAP7_75t_R c8306(
.A(net6560),
.B(net10311),
.CON(net8342)
);

INVx13_ASAP7_75t_R c8307(
.A(net3767),
.Y(net8343)
);

NAND2x1_ASAP7_75t_R c8308(
.A(net7397),
.B(net5628),
.Y(net8344)
);

NAND2x1p5_ASAP7_75t_R c8309(
.A(net8317),
.B(net8280),
.Y(net8345)
);

NAND2x2_ASAP7_75t_R c8310(
.A(net5576),
.B(net8256),
.Y(net8346)
);

INVx1_ASAP7_75t_R c8311(
.A(net8261),
.Y(net8347)
);

NAND2xp33_ASAP7_75t_R c8312(
.A(net8342),
.B(net6612),
.Y(net8348)
);

INVx2_ASAP7_75t_R c8313(
.A(net10294),
.Y(net8349)
);

NAND2xp5_ASAP7_75t_R c8314(
.A(net8322),
.B(net6542),
.Y(net8350)
);

INVx3_ASAP7_75t_R c8315(
.A(net8273),
.Y(net8351)
);

NAND2xp67_ASAP7_75t_R c8316(
.A(net6480),
.B(net3767),
.Y(net8352)
);

NOR2x1_ASAP7_75t_R c8317(
.A(net8320),
.B(net10312),
.Y(net8353)
);

INVx4_ASAP7_75t_R c8318(
.A(net10297),
.Y(net8354)
);

NOR2x1p5_ASAP7_75t_R c8319(
.A(net7382),
.B(net8279),
.Y(net8355)
);

NOR2x2_ASAP7_75t_R c8320(
.A(net8330),
.B(net6519),
.Y(net8356)
);

NOR2xp33_ASAP7_75t_R c8321(
.A(net8333),
.B(net10312),
.Y(net8357)
);

NOR2xp67_ASAP7_75t_R c8322(
.A(net8324),
.B(net8337),
.Y(net8358)
);

INVx5_ASAP7_75t_R c8323(
.A(net8353),
.Y(net8359)
);

OR2x2_ASAP7_75t_R c8324(
.A(net8349),
.B(net10294),
.Y(net8360)
);

INVx6_ASAP7_75t_R c8325(
.A(net8348),
.Y(net8361)
);

OR3x1_ASAP7_75t_R c8326(
.A(net8359),
.B(net5588),
.C(net8358),
.Y(net8362)
);

OR2x4_ASAP7_75t_R c8327(
.A(net7513),
.B(net7404),
.Y(net8363)
);

INVx8_ASAP7_75t_R c8328(
.A(net8289),
.Y(net8364)
);

OR2x6_ASAP7_75t_R c8329(
.A(net7461),
.B(net10278),
.Y(net8365)
);

INVxp33_ASAP7_75t_R c8330(
.A(net8299),
.Y(net8366)
);

INVxp67_ASAP7_75t_R c8331(
.A(net9187),
.Y(net8367)
);

XNOR2x1_ASAP7_75t_R c8332(
.B(net8263),
.A(net8344),
.Y(net8368)
);

XNOR2x2_ASAP7_75t_R c8333(
.A(net8356),
.B(net8282),
.Y(net8369)
);

SDFHx2_ASAP7_75t_R c8334(
.D(net8311),
.SE(net8366),
.SI(net8323),
.CLK(clk),
.QN(net8370)
);

OR3x2_ASAP7_75t_R c8335(
.A(net8354),
.B(net6615),
.C(net7513),
.Y(net8371)
);

XNOR2xp5_ASAP7_75t_R c8336(
.A(net8361),
.B(net8366),
.Y(net8372)
);

XOR2x1_ASAP7_75t_R c8337(
.A(net7526),
.B(net9737),
.Y(net8373)
);

XOR2x2_ASAP7_75t_R c8338(
.A(net8256),
.B(net8293),
.Y(net8374)
);

OR3x4_ASAP7_75t_R c8339(
.A(net7420),
.B(net8365),
.C(net8347),
.Y(net8375)
);

BUFx10_ASAP7_75t_R c8340(
.A(net10405),
.Y(net8376)
);

XOR2xp5_ASAP7_75t_R c8341(
.A(net8340),
.B(net8367),
.Y(net8377)
);

BUFx12_ASAP7_75t_R c8342(
.A(net8363),
.Y(net8378)
);

ICGx5_ASAP7_75t_R c8343(
.ENA(net8377),
.SE(net8363),
.CLK(clk),
.GCLK(net8379)
);

AND2x2_ASAP7_75t_R c8344(
.A(net8365),
.B(net8357),
.Y(net8380)
);

BUFx12f_ASAP7_75t_R c8345(
.A(net8351),
.Y(net8381)
);

AND3x1_ASAP7_75t_R c8346(
.A(net8307),
.B(net8352),
.C(net8273),
.Y(net8382)
);

AND2x4_ASAP7_75t_R c8347(
.A(net8280),
.B(net8273),
.Y(net8383)
);

AND2x6_ASAP7_75t_R c8348(
.A(net8380),
.B(net8365),
.Y(net8384)
);

BUFx16f_ASAP7_75t_R c8349(
.A(net10559),
.Y(net8385)
);

ICGx5p33DC_ASAP7_75t_R c8350(
.ENA(net8282),
.SE(net8311),
.CLK(clk),
.GCLK(net8386)
);

HAxp5_ASAP7_75t_R c8351(
.A(net8371),
.B(net8381),
.CON(net8388),
.SN(net8387)
);

NAND2x1_ASAP7_75t_R c8352(
.A(net7387),
.B(net8361),
.Y(net8389)
);

AND3x2_ASAP7_75t_R c8353(
.A(net8301),
.B(net8363),
.C(net8352),
.Y(net8390)
);

NAND2x1p5_ASAP7_75t_R c8354(
.A(net8379),
.B(net8375),
.Y(net8391)
);

AND3x4_ASAP7_75t_R c8355(
.A(net8262),
.B(net8388),
.C(net6560),
.Y(net8392)
);

AO221x1_ASAP7_75t_R c8356(
.A1(net8345),
.A2(net8367),
.B1(net8386),
.B2(net8366),
.C(net8376),
.Y(net8393)
);

AO21x1_ASAP7_75t_R c8357(
.A1(net8303),
.A2(net8378),
.B(net7466),
.Y(net8394)
);

AO21x2_ASAP7_75t_R c8358(
.A1(net8372),
.A2(net8386),
.B(net8387),
.Y(net8395)
);

SDFHx3_ASAP7_75t_R c8359(
.D(net8390),
.SE(net8320),
.SI(net7382),
.CLK(clk),
.QN(net8396)
);

AOI21x1_ASAP7_75t_R c8360(
.A1(net8333),
.A2(net8379),
.B(net8386),
.Y(net8397)
);

NAND2x2_ASAP7_75t_R c8361(
.A(net7514),
.B(net8296),
.Y(net8398)
);

AOI21xp33_ASAP7_75t_R c8362(
.A1(net8375),
.A2(net8396),
.B(net8367),
.Y(net8399)
);

AOI21xp5_ASAP7_75t_R c8363(
.A1(net8398),
.A2(net8397),
.B(net8396),
.Y(net8400)
);

FAx1_ASAP7_75t_R c8364(
.A(net6521),
.B(net8399),
.CI(net10297),
.SN(net8401)
);

MAJIxp5_ASAP7_75t_R c8365(
.A(net6554),
.B(net5689),
.C(net8357),
.Y(net8402)
);

NAND2xp33_ASAP7_75t_R c8366(
.A(net8401),
.B(net8396),
.Y(net8403)
);

MAJx2_ASAP7_75t_R c8367(
.A(net8312),
.B(net8388),
.C(net8323),
.Y(net8404)
);

MAJx3_ASAP7_75t_R c8368(
.A(net8403),
.B(net8387),
.C(net9951),
.Y(net8405)
);

NAND2xp5_ASAP7_75t_R c8369(
.A(net8386),
.B(net8400),
.Y(net8406)
);

NAND3x1_ASAP7_75t_R c8370(
.A(net5532),
.B(net8318),
.C(net8403),
.Y(net8407)
);

NAND2xp67_ASAP7_75t_R c8371(
.A(net8369),
.B(net8336),
.Y(net8408)
);

NAND3x2_ASAP7_75t_R c8372(
.B(net8406),
.C(net8389),
.A(net8307),
.Y(net8409)
);

SDFHx4_ASAP7_75t_R c8373(
.D(net8378),
.SE(net8408),
.SI(net9975),
.CLK(clk),
.QN(net8410)
);

NAND3xp33_ASAP7_75t_R c8374(
.A(net8409),
.B(net8408),
.C(net8383),
.Y(net8411)
);

NOR3x1_ASAP7_75t_R c8375(
.A(net8384),
.B(net8404),
.C(net7420),
.Y(net8412)
);

AO221x2_ASAP7_75t_R c8376(
.A1(net8402),
.A2(net7526),
.B1(net8400),
.B2(net7456),
.C(net8258),
.Y(net8413)
);

NOR2x1_ASAP7_75t_R c8377(
.A(net8389),
.B(net8379),
.Y(net8414)
);

AOI222xp33_ASAP7_75t_R c8378(
.A1(net8358),
.A2(net8414),
.B1(net8397),
.B2(net8376),
.C1(net7469),
.C2(net10313),
.Y(net8415)
);

NOR3x2_ASAP7_75t_R c8379(
.B(net8382),
.C(net4652),
.A(net9830),
.Y(net8416)
);

NOR3xp33_ASAP7_75t_R c8380(
.A(net8403),
.B(net7500),
.C(net8410),
.Y(net8417)
);

O2A1O1Ixp5_ASAP7_75t_R c8381(
.A1(net8341),
.A2(net8409),
.B(net7456),
.C(net9817),
.Y(net8418)
);

OA211x2_ASAP7_75t_R c8382(
.A1(net9737),
.A2(net9800),
.B(net10313),
.C(net10314),
.Y(net8419)
);

NOR2x1p5_ASAP7_75t_R c8383(
.A(net6681),
.B(net6615),
.Y(net8420)
);

NOR2x2_ASAP7_75t_R c8384(
.A(net7461),
.B(net8293),
.Y(net8421)
);

NOR2xp33_ASAP7_75t_R c8385(
.A(net8400),
.B(net10279),
.Y(net8422)
);

NOR2xp67_ASAP7_75t_R c8386(
.A(net8376),
.B(net9789),
.Y(net8423)
);

OA21x2_ASAP7_75t_R c8387(
.A1(net7499),
.A2(net8410),
.B(net8279),
.Y(net8424)
);

OR2x2_ASAP7_75t_R c8388(
.A(net8421),
.B(net7585),
.Y(net8425)
);

BUFx24_ASAP7_75t_R c8389(
.A(net10115),
.Y(net8426)
);

BUFx2_ASAP7_75t_R c8390(
.A(net8325),
.Y(net8427)
);

BUFx3_ASAP7_75t_R c8391(
.A(net10433),
.Y(net8428)
);

OR2x4_ASAP7_75t_R c8392(
.A(net8341),
.B(net7570),
.Y(net8429)
);

OR2x6_ASAP7_75t_R c8393(
.A(net8426),
.B(net6690),
.Y(net8430)
);

XNOR2x1_ASAP7_75t_R c8394(
.B(net7414),
.A(net4835),
.Y(net8431)
);

AO32x1_ASAP7_75t_R c8395(
.A1(net8352),
.A2(net8408),
.A3(net7615),
.B1(net7574),
.B2(net8376),
.Y(net8432)
);

XNOR2x2_ASAP7_75t_R c8396(
.A(net8343),
.B(net5772),
.Y(net8433)
);

XNOR2xp5_ASAP7_75t_R c8397(
.A(net8346),
.B(net10313),
.Y(net8434)
);

XOR2x1_ASAP7_75t_R c8398(
.A(net7570),
.B(net8427),
.Y(net8435)
);

XOR2x2_ASAP7_75t_R c8399(
.A(net8383),
.B(net8424),
.Y(net8436)
);

XOR2xp5_ASAP7_75t_R c8400(
.A(net8431),
.B(net10314),
.Y(net8437)
);

AND2x2_ASAP7_75t_R c8401(
.A(net6682),
.B(net8293),
.Y(net8438)
);

AND2x4_ASAP7_75t_R c8402(
.A(net8367),
.B(net8279),
.Y(net8439)
);

BUFx4_ASAP7_75t_R c8403(
.A(net10513),
.Y(net8440)
);

AND2x6_ASAP7_75t_R c8404(
.A(net7374),
.B(net8391),
.Y(net8441)
);

SDFLx1_ASAP7_75t_R c8405(
.D(net8439),
.SE(net7477),
.SI(net8352),
.CLK(clk),
.QN(net8442)
);

HAxp5_ASAP7_75t_R c8406(
.A(net6527),
.B(net8440),
.CON(net8443)
);

OAI21x1_ASAP7_75t_R c8407(
.A1(net7526),
.A2(net8431),
.B(net8435),
.Y(net8444)
);

NAND2x1_ASAP7_75t_R c8408(
.A(net8400),
.B(net9706),
.Y(net8445)
);

BUFx4f_ASAP7_75t_R c8409(
.A(net10486),
.Y(net8446)
);

BUFx5_ASAP7_75t_R c8410(
.A(net10492),
.Y(net8447)
);

NAND2x1p5_ASAP7_75t_R c8411(
.A(net4852),
.B(net8445),
.Y(net8448)
);

NAND2x2_ASAP7_75t_R c8412(
.A(net6690),
.B(net8367),
.Y(net8449)
);

NAND2xp33_ASAP7_75t_R c8413(
.A(net8264),
.B(net8385),
.Y(net8450)
);

OAI21xp33_ASAP7_75t_R c8414(
.A1(net8339),
.A2(net7617),
.B(net6542),
.Y(net8451)
);

NAND2xp5_ASAP7_75t_R c8415(
.A(net8385),
.B(net8442),
.Y(net8452)
);

OAI21xp5_ASAP7_75t_R c8416(
.A1(net8449),
.A2(net8325),
.B(net7374),
.Y(net8453)
);

OR3x1_ASAP7_75t_R c8417(
.A(net7494),
.B(net7542),
.C(net8452),
.Y(net8454)
);

NAND2xp67_ASAP7_75t_R c8418(
.A(net8296),
.B(net8450),
.Y(net8455)
);

NOR2x1_ASAP7_75t_R c8419(
.A(net8410),
.B(net10050),
.Y(net8456)
);

BUFx6f_ASAP7_75t_R c8420(
.A(net10433),
.Y(net8457)
);

NOR2x1p5_ASAP7_75t_R c8421(
.A(net8293),
.B(net8393),
.Y(net8458)
);

BUFx8_ASAP7_75t_R c8422(
.A(net10338),
.Y(net8459)
);

NOR2x2_ASAP7_75t_R c8423(
.A(net6630),
.B(net6649),
.Y(net8460)
);

AO32x2_ASAP7_75t_R c8424(
.A1(net8360),
.A2(net3767),
.A3(net8420),
.B1(net10050),
.B2(net10313),
.Y(net8461)
);

OA22x2_ASAP7_75t_R c8425(
.A1(net7508),
.A2(net8433),
.B1(net8435),
.B2(net8431),
.Y(net8462)
);

SDFLx2_ASAP7_75t_R c8426(
.D(net8456),
.SE(net8425),
.SI(net8460),
.CLK(clk),
.QN(net8463)
);

OA31x2_ASAP7_75t_R c8427(
.A1(net8395),
.A2(net8460),
.A3(net8397),
.B1(net10313),
.Y(net8464)
);

NOR2xp33_ASAP7_75t_R c8428(
.A(net8435),
.B(net7617),
.Y(net8465)
);

AOI221x1_ASAP7_75t_R c8429(
.A1(net8394),
.A2(net8454),
.B1(net8419),
.B2(net7469),
.C(net8366),
.Y(net8466)
);

NOR2xp67_ASAP7_75t_R c8430(
.A(net8433),
.B(net10083),
.Y(net8467)
);

OR2x2_ASAP7_75t_R c8431(
.A(net8397),
.B(net10316),
.Y(net8468)
);

OR3x2_ASAP7_75t_R c8432(
.A(net6542),
.B(net8258),
.C(net8337),
.Y(net8469)
);

OAI211xp5_ASAP7_75t_R c8433(
.A1(net8318),
.A2(net7544),
.B(net8425),
.C(net8294),
.Y(net8470)
);

AOI221xp5_ASAP7_75t_R c8434(
.A1(net8446),
.A2(net8444),
.B1(net5772),
.B2(net8260),
.C(net10315),
.Y(net8471)
);

OR3x4_ASAP7_75t_R c8435(
.A(net8431),
.B(net8433),
.C(net10315),
.Y(net8472)
);

ICGx6p67DC_ASAP7_75t_R c8436(
.ENA(net8279),
.SE(net7566),
.CLK(clk),
.GCLK(net8473)
);

OR2x4_ASAP7_75t_R c8437(
.A(net8315),
.B(net10009),
.Y(net8474)
);

OR2x6_ASAP7_75t_R c8438(
.A(net8430),
.B(net8445),
.Y(net8475)
);

CKINVDCx10_ASAP7_75t_R c8439(
.A(net10115),
.Y(net8476)
);

XNOR2x1_ASAP7_75t_R c8440(
.B(net8373),
.A(net7615),
.Y(net8477)
);

XNOR2x2_ASAP7_75t_R c8441(
.A(net8443),
.B(net7544),
.Y(net8478)
);

CKINVDCx11_ASAP7_75t_R c8442(
.A(net10553),
.Y(net8479)
);

XNOR2xp5_ASAP7_75t_R c8443(
.A(net8457),
.B(net8463),
.Y(net8480)
);

XOR2x1_ASAP7_75t_R c8444(
.A(net8480),
.B(net5726),
.Y(net8481)
);

XOR2x2_ASAP7_75t_R c8445(
.A(net7544),
.B(net8444),
.Y(net8482)
);

XOR2xp5_ASAP7_75t_R c8446(
.A(net8450),
.B(net8400),
.Y(net8483)
);

AND2x2_ASAP7_75t_R c8447(
.A(net8483),
.B(net9965),
.Y(net8484)
);

AND2x4_ASAP7_75t_R c8448(
.A(net8447),
.B(net8410),
.Y(net8485)
);

AND3x1_ASAP7_75t_R c8449(
.A(net8455),
.B(net8483),
.C(net10315),
.Y(net8486)
);

AND2x6_ASAP7_75t_R c8450(
.A(net8483),
.B(net10314),
.Y(net8487)
);

HAxp5_ASAP7_75t_R c8451(
.A(net7615),
.B(net10083),
.CON(net8489),
.SN(net8488)
);

CKINVDCx12_ASAP7_75t_R c8452(
.A(net10338),
.Y(net8490)
);

AND3x2_ASAP7_75t_R c8453(
.A(net8350),
.B(net8433),
.C(net10316),
.Y(net8491)
);

AND3x4_ASAP7_75t_R c8454(
.A(net8490),
.B(net8451),
.C(net8480),
.Y(net8492)
);

CKINVDCx14_ASAP7_75t_R c8455(
.A(net10459),
.Y(net8493)
);

NAND2x1_ASAP7_75t_R c8456(
.A(net8461),
.B(net8480),
.Y(net8494)
);

AO21x1_ASAP7_75t_R c8457(
.A1(net6649),
.A2(net7494),
.B(net10123),
.Y(net8495)
);

NAND2x1p5_ASAP7_75t_R c8458(
.A(net8474),
.B(net8476),
.Y(net8496)
);

AO21x2_ASAP7_75t_R c8459(
.A1(net6694),
.A2(net9706),
.B(net10315),
.Y(net8497)
);

NAND2x2_ASAP7_75t_R c8460(
.A(net8497),
.B(net8487),
.Y(net8498)
);

NAND2xp33_ASAP7_75t_R c8461(
.A(net8374),
.B(net6643),
.Y(net8499)
);

AOI21x1_ASAP7_75t_R c8462(
.A1(net8482),
.A2(net8494),
.B(net8463),
.Y(net8500)
);

OAI22x1_ASAP7_75t_R c8463(
.A1(net7617),
.A2(net8488),
.B1(net8374),
.B2(net8478),
.Y(net8501)
);

AOI311xp33_ASAP7_75t_R c8464(
.A1(net8498),
.A2(net8496),
.A3(net8499),
.B(net8480),
.C(net7393),
.Y(net8502)
);

NAND2xp5_ASAP7_75t_R c8465(
.A(net8465),
.B(net10318),
.Y(net8503)
);

CKINVDCx16_ASAP7_75t_R c8466(
.A(net10093),
.Y(net8504)
);

NAND2xp67_ASAP7_75t_R c8467(
.A(net6612),
.B(net8493),
.Y(net8505)
);

CKINVDCx20_ASAP7_75t_R c8468(
.A(net10053),
.Y(net8506)
);

NOR2x1_ASAP7_75t_R c8469(
.A(net6705),
.B(net7658),
.Y(net8507)
);

AOI21xp33_ASAP7_75t_R c8470(
.A1(net7550),
.A2(net8267),
.B(net7399),
.Y(net8508)
);

AOI21xp5_ASAP7_75t_R c8471(
.A1(net7675),
.A2(net8460),
.B(net10052),
.Y(net8509)
);

CKINVDCx5p33_ASAP7_75t_R c8472(
.A(net10121),
.Y(net8510)
);

NOR2x1p5_ASAP7_75t_R c8473(
.A(net8509),
.B(net10166),
.Y(net8511)
);

CKINVDCx6p67_ASAP7_75t_R c8474(
.A(net10521),
.Y(net8512)
);

FAx1_ASAP7_75t_R c8475(
.A(net8391),
.B(net8479),
.CI(net8442),
.SN(net8514),
.CON(net8513)
);

NOR2x2_ASAP7_75t_R c8476(
.A(net7500),
.B(net7647),
.Y(net8515)
);

MAJIxp5_ASAP7_75t_R c8477(
.A(net7698),
.B(net8493),
.C(net8431),
.Y(net8516)
);

NOR2xp33_ASAP7_75t_R c8478(
.A(net7541),
.B(net6705),
.Y(net8517)
);

NOR2xp67_ASAP7_75t_R c8479(
.A(net7653),
.B(net7636),
.Y(net8518)
);

MAJx2_ASAP7_75t_R c8480(
.A(net3922),
.B(net8518),
.C(net8444),
.Y(net8519)
);

OR2x2_ASAP7_75t_R c8481(
.A(net5628),
.B(net8357),
.Y(net8520)
);

OR2x4_ASAP7_75t_R c8482(
.A(net5841),
.B(net8514),
.Y(net8521)
);

MAJx3_ASAP7_75t_R c8483(
.A(net6782),
.B(net6560),
.C(net8260),
.Y(net8522)
);

OR2x6_ASAP7_75t_R c8484(
.A(net7473),
.B(net10171),
.Y(net8523)
);

XNOR2x1_ASAP7_75t_R c8485(
.B(net6781),
.A(net7606),
.Y(net8524)
);

NAND3x1_ASAP7_75t_R c8486(
.A(net7547),
.B(net8258),
.C(net9938),
.Y(net8525)
);

SDFLx3_ASAP7_75t_R c8487(
.D(net6747),
.SE(net8444),
.SI(net8357),
.CLK(clk),
.QN(net8526)
);

ICGx8DC_ASAP7_75t_R c8488(
.ENA(net5772),
.SE(net8495),
.CLK(clk),
.GCLK(net8527)
);

NAND3x2_ASAP7_75t_R c8489(
.B(net8364),
.C(net8344),
.A(net7453),
.Y(net8528)
);

NAND3xp33_ASAP7_75t_R c8490(
.A(net7641),
.B(net8445),
.C(net8315),
.Y(net8529)
);

XNOR2x2_ASAP7_75t_R c8491(
.A(net6666),
.B(net10014),
.Y(net8530)
);

SDFLx4_ASAP7_75t_R c8492(
.D(net8508),
.SE(net7670),
.SI(net8419),
.CLK(clk),
.QN(net8531)
);

NOR3x1_ASAP7_75t_R c8493(
.A(net8522),
.B(net7574),
.C(net7500),
.Y(net8532)
);

NOR3x2_ASAP7_75t_R c8494(
.B(net8423),
.C(net8523),
.A(net8376),
.Y(net8533)
);

XNOR2xp5_ASAP7_75t_R c8495(
.A(net8473),
.B(net10317),
.Y(net8534)
);

ICGx1_ASAP7_75t_R c8496(
.ENA(net7670),
.SE(net8506),
.CLK(clk),
.GCLK(net8535)
);

DFFASRHQNx1_ASAP7_75t_R c8497(
.D(net8392),
.RESETN(net7658),
.SETN(net8522),
.CLK(clk),
.QN(net8536)
);

XOR2x1_ASAP7_75t_R c8498(
.A(net6761),
.B(net5628),
.Y(net8537)
);

NOR3xp33_ASAP7_75t_R c8499(
.A(net7611),
.B(net8473),
.C(net8438),
.Y(net8538)
);

XOR2x2_ASAP7_75t_R c8500(
.A(net7637),
.B(net8267),
.Y(net8539)
);

XOR2xp5_ASAP7_75t_R c8501(
.A(net8532),
.B(net7542),
.Y(net8540)
);

CKINVDCx8_ASAP7_75t_R c8502(
.A(net10521),
.Y(net8541)
);

AND2x2_ASAP7_75t_R c8503(
.A(net8473),
.B(net9947),
.Y(net8542)
);

AND2x4_ASAP7_75t_R c8504(
.A(net8542),
.B(net10318),
.Y(net8543)
);

AND2x6_ASAP7_75t_R c8505(
.A(net8499),
.B(net10316),
.Y(net8544)
);

HAxp5_ASAP7_75t_R c8506(
.A(net8260),
.B(net8463),
.CON(net8546),
.SN(net8545)
);

NAND2x1_ASAP7_75t_R c8507(
.A(net6666),
.B(net8540),
.Y(net8547)
);

NAND2x1p5_ASAP7_75t_R c8508(
.A(net8503),
.B(net8509),
.Y(net8548)
);

SDFHx1_ASAP7_75t_R c8509(
.D(net7399),
.SE(net8536),
.SI(net8521),
.CLK(clk),
.QN(net8549)
);

OA21x2_ASAP7_75t_R c8510(
.A1(net8517),
.A2(net6705),
.B(net8370),
.Y(net8550)
);

NAND2x2_ASAP7_75t_R c8511(
.A(net7669),
.B(net9991),
.Y(net8551)
);

CKINVDCx9p33_ASAP7_75t_R c8512(
.A(net10539),
.Y(net8552)
);

ICGx2_ASAP7_75t_R c8513(
.ENA(net8538),
.SE(net8267),
.CLK(clk),
.GCLK(net8553)
);

NAND2xp33_ASAP7_75t_R c8514(
.A(net8549),
.B(net8459),
.Y(net8554)
);

OAI21x1_ASAP7_75t_R c8515(
.A1(net8515),
.A2(net8336),
.B(net6761),
.Y(net8555)
);

OAI21xp33_ASAP7_75t_R c8516(
.A1(net8535),
.A2(net8493),
.B(net8440),
.Y(net8556)
);

NAND2xp5_ASAP7_75t_R c8517(
.A(net6649),
.B(net8553),
.Y(net8557)
);

NAND2xp67_ASAP7_75t_R c8518(
.A(net8557),
.B(net8440),
.Y(net8558)
);

NOR2x1_ASAP7_75t_R c8519(
.A(net8485),
.B(net8364),
.Y(net8559)
);

NOR2x1p5_ASAP7_75t_R c8520(
.A(net8555),
.B(net8558),
.Y(net8560)
);

NOR2x2_ASAP7_75t_R c8521(
.A(net8556),
.B(net8294),
.Y(net8561)
);

OAI21xp5_ASAP7_75t_R c8522(
.A1(net7547),
.A2(net7675),
.B(net8392),
.Y(net8562)
);

OR3x1_ASAP7_75t_R c8523(
.A(net8511),
.B(net8370),
.C(net8509),
.Y(net8563)
);

HB1xp67_ASAP7_75t_R c8524(
.A(net10053),
.Y(net8564)
);

NOR2xp33_ASAP7_75t_R c8525(
.A(net8431),
.B(net9938),
.Y(net8565)
);

OAI22xp33_ASAP7_75t_R c8526(
.A1(net8557),
.A2(net8535),
.B1(net7688),
.B2(net10145),
.Y(net8566)
);

NOR2xp67_ASAP7_75t_R c8527(
.A(net8554),
.B(net6711),
.Y(net8567)
);

OR2x2_ASAP7_75t_R c8528(
.A(net8552),
.B(net9929),
.Y(net8568)
);

SDFHx2_ASAP7_75t_R c8529(
.D(net8568),
.SE(net8521),
.SI(net8564),
.CLK(clk),
.QN(net8569)
);

OR3x2_ASAP7_75t_R c8530(
.A(net8260),
.B(net8508),
.C(net9867),
.Y(net8570)
);

OR3x4_ASAP7_75t_R c8531(
.A(net7541),
.B(net8554),
.C(net10134),
.Y(net8571)
);

AND3x1_ASAP7_75t_R c8532(
.A(net8540),
.B(net8551),
.C(net8566),
.Y(net8572)
);

OR2x4_ASAP7_75t_R c8533(
.A(net8536),
.B(net8565),
.Y(net8573)
);

SDFHx3_ASAP7_75t_R c8534(
.D(net8344),
.SE(net8549),
.SI(net8478),
.CLK(clk),
.QN(net8574)
);

SDFHx4_ASAP7_75t_R c8535(
.D(net8336),
.SE(net8559),
.SI(net8574),
.CLK(clk),
.QN(net8575)
);

AND3x2_ASAP7_75t_R c8536(
.A(net8564),
.B(net8549),
.C(net8574),
.Y(net8576)
);

AND3x4_ASAP7_75t_R c8537(
.A(net8520),
.B(net8573),
.C(net8574),
.Y(net8577)
);

AO21x1_ASAP7_75t_R c8538(
.A1(net6734),
.A2(net8574),
.B(net7640),
.Y(net8578)
);

AO21x2_ASAP7_75t_R c8539(
.A1(net8565),
.A2(net9863),
.B(net9886),
.Y(net8579)
);

AOI21x1_ASAP7_75t_R c8540(
.A1(net8571),
.A2(net8557),
.B(net8513),
.Y(net8580)
);

AOI21xp33_ASAP7_75t_R c8541(
.A1(net8444),
.A2(net8534),
.B(net10052),
.Y(net8581)
);

AOI21xp5_ASAP7_75t_R c8542(
.A1(net8567),
.A2(net8575),
.B(net9912),
.Y(net8582)
);

SDFLx1_ASAP7_75t_R c8543(
.D(net8581),
.SE(net9975),
.SI(net10171),
.CLK(clk),
.QN(net8583)
);

FAx1_ASAP7_75t_R c8544(
.A(net8528),
.B(net8580),
.CI(net8583),
.SN(net8584)
);

OAI22xp5_ASAP7_75t_R c8545(
.A1(net8550),
.A2(net8561),
.B1(net8515),
.B2(net10313),
.Y(net8585)
);

OR2x6_ASAP7_75t_R c8546(
.A(net7664),
.B(net9785),
.Y(net8586)
);

AOI32xp33_ASAP7_75t_R c8547(
.A1(net8586),
.A2(net8582),
.A3(net8576),
.B1(net8574),
.B2(net7651),
.Y(net8587)
);

MAJIxp5_ASAP7_75t_R c8548(
.A(net8574),
.B(net9705),
.C(net9774),
.Y(net8588)
);

MAJx2_ASAP7_75t_R c8549(
.A(net7606),
.B(net8569),
.C(net8531),
.Y(net8589)
);

MAJx3_ASAP7_75t_R c8550(
.A(net7783),
.B(net8521),
.C(net8566),
.Y(net8590)
);

HB2xp67_ASAP7_75t_R c8551(
.A(net10092),
.Y(net8591)
);

XNOR2x1_ASAP7_75t_R c8552(
.B(net6560),
.A(net10318),
.Y(net8592)
);

XNOR2x2_ASAP7_75t_R c8553(
.A(net7704),
.B(net8489),
.Y(net8593)
);

XNOR2xp5_ASAP7_75t_R c8554(
.A(net7721),
.B(net8553),
.Y(net8594)
);

NAND3x1_ASAP7_75t_R c8555(
.A(net8428),
.B(net8593),
.C(net8575),
.Y(net8595)
);

XOR2x1_ASAP7_75t_R c8556(
.A(net8527),
.B(net8458),
.Y(net8596)
);

NAND3x2_ASAP7_75t_R c8557(
.B(net8533),
.C(net8575),
.A(net8486),
.Y(net8597)
);

NAND3xp33_ASAP7_75t_R c8558(
.A(net7473),
.B(net8484),
.C(net8593),
.Y(net8598)
);

AOI321xp33_ASAP7_75t_R c8559(
.A1(net8438),
.A2(net4962),
.A3(net8592),
.B1(net8521),
.B2(net8541),
.C(net8569),
.Y(net8599)
);

NOR3x1_ASAP7_75t_R c8560(
.A(net7597),
.B(net8506),
.C(net7683),
.Y(net8600)
);

NOR3x2_ASAP7_75t_R c8561(
.B(net8489),
.C(net8595),
.A(net8545),
.Y(net8601)
);

XOR2x2_ASAP7_75t_R c8562(
.A(net8294),
.B(net8601),
.Y(net8602)
);

ICGx2p67DC_ASAP7_75t_R c8563(
.ENA(net8388),
.SE(net8521),
.CLK(clk),
.GCLK(net8603)
);

NOR3xp33_ASAP7_75t_R c8564(
.A(net7453),
.B(net8603),
.C(net8463),
.Y(net8604)
);

HB3xp67_ASAP7_75t_R c8565(
.A(net10552),
.Y(net8605)
);

OA21x2_ASAP7_75t_R c8566(
.A1(net8524),
.A2(net7597),
.B(net7774),
.Y(net8606)
);

XOR2xp5_ASAP7_75t_R c8567(
.A(net8541),
.B(net8505),
.Y(net8607)
);

OAI21x1_ASAP7_75t_R c8568(
.A1(net8486),
.A2(net8294),
.B(net7784),
.Y(net8608)
);

HB4xp67_ASAP7_75t_R c8569(
.A(net10574),
.Y(net8609)
);

AND2x2_ASAP7_75t_R c8570(
.A(net7618),
.B(net8445),
.Y(net8610)
);

OAI21xp33_ASAP7_75t_R c8571(
.A1(net8543),
.A2(net8583),
.B(net9965),
.Y(net8611)
);

AND2x4_ASAP7_75t_R c8572(
.A(net8546),
.B(net8419),
.Y(net8612)
);

AND2x6_ASAP7_75t_R c8573(
.A(net8477),
.B(net8570),
.Y(net8613)
);

OAI21xp5_ASAP7_75t_R c8574(
.A1(net8610),
.A2(net7784),
.B(net7688),
.Y(net8614)
);

OR3x1_ASAP7_75t_R c8575(
.A(net7781),
.B(net8387),
.C(net10300),
.Y(net8615)
);

OR3x2_ASAP7_75t_R c8576(
.A(net7784),
.B(net8315),
.C(net5689),
.Y(net8616)
);

OR3x4_ASAP7_75t_R c8577(
.A(net5846),
.B(net8580),
.C(net6804),
.Y(net8617)
);

HAxp5_ASAP7_75t_R c8578(
.A(net7647),
.B(net7669),
.CON(net8619),
.SN(net8618)
);

AND3x1_ASAP7_75t_R c8579(
.A(net8587),
.B(net9942),
.C(net10317),
.Y(net8620)
);

SDFLx2_ASAP7_75t_R c8580(
.D(net8463),
.SE(net8588),
.SI(net6796),
.CLK(clk),
.QN(net8621)
);

NAND2x1_ASAP7_75t_R c8581(
.A(net9947),
.B(net10300),
.Y(net8622)
);

AND3x2_ASAP7_75t_R c8582(
.A(net7707),
.B(net8591),
.C(net8516),
.Y(net8623)
);

AOI33xp33_ASAP7_75t_R c8583(
.A1(net7640),
.A2(net8516),
.A3(net8592),
.B1(net8622),
.B2(net8606),
.B3(net7765),
.Y(net8624)
);

AND3x4_ASAP7_75t_R c8584(
.A(net7724),
.B(net8258),
.C(net8516),
.Y(net8625)
);

NAND2x1p5_ASAP7_75t_R c8585(
.A(net7620),
.B(net8526),
.Y(net8626)
);

AO21x1_ASAP7_75t_R c8586(
.A1(net8499),
.A2(net8616),
.B(net8347),
.Y(net8627)
);

AO21x2_ASAP7_75t_R c8587(
.A1(net7729),
.A2(net7456),
.B(net7747),
.Y(net8628)
);

AOI21x1_ASAP7_75t_R c8588(
.A1(net8612),
.A2(net8591),
.B(net7774),
.Y(net8629)
);

SDFLx3_ASAP7_75t_R c8589(
.D(net8603),
.SE(net8601),
.SI(net7774),
.CLK(clk),
.QN(net8630)
);

SDFLx4_ASAP7_75t_R c8590(
.D(net7469),
.SE(net8613),
.SI(net6796),
.CLK(clk),
.QN(net8631)
);

DFFASRHQNx1_ASAP7_75t_R c8591(
.D(net8559),
.RESETN(net8631),
.SETN(net9912),
.CLK(clk),
.QN(net8632)
);

AOI21xp33_ASAP7_75t_R c8592(
.A1(net8628),
.A2(net8613),
.B(net7618),
.Y(net8633)
);

AOI21xp5_ASAP7_75t_R c8593(
.A1(net6796),
.A2(net8614),
.B(net8294),
.Y(net8634)
);

FAx1_ASAP7_75t_R c8594(
.A(net8510),
.B(net8616),
.CI(net7667),
.SN(net8636),
.CON(net8635)
);

MAJIxp5_ASAP7_75t_R c8595(
.A(net8452),
.B(net8618),
.C(net5846),
.Y(net8637)
);

MAJx2_ASAP7_75t_R c8596(
.A(net8258),
.B(net8337),
.C(net8608),
.Y(net8638)
);

MAJx3_ASAP7_75t_R c8597(
.A(net8437),
.B(net7786),
.C(net8507),
.Y(net8639)
);

SDFHx1_ASAP7_75t_R c8598(
.D(net8608),
.SE(net10283),
.SI(net10317),
.CLK(clk),
.QN(net8640)
);

NAND3x1_ASAP7_75t_R c8599(
.A(net8637),
.B(net8451),
.C(net8621),
.Y(net8641)
);

NAND3x2_ASAP7_75t_R c8600(
.B(net7774),
.C(net8635),
.A(net8621),
.Y(net8642)
);

NAND3xp33_ASAP7_75t_R c8601(
.A(net7683),
.B(net8451),
.C(net8632),
.Y(net8643)
);

SDFHx2_ASAP7_75t_R c8602(
.D(net8445),
.SE(net8597),
.SI(net8531),
.CLK(clk),
.QN(net8644)
);

NOR3x1_ASAP7_75t_R c8603(
.A(net8600),
.B(net8595),
.C(net10014),
.Y(net8645)
);

SDFHx3_ASAP7_75t_R c8604(
.D(net8608),
.SE(net8619),
.SI(net8527),
.CLK(clk),
.QN(net8646)
);

INVx11_ASAP7_75t_R c8605(
.A(net10092),
.Y(net8647)
);

INVx13_ASAP7_75t_R c8606(
.A(net10439),
.Y(net8648)
);

NOR3x2_ASAP7_75t_R c8607(
.B(net8419),
.C(net8605),
.A(net10283),
.Y(net8649)
);

NAND5xp2_ASAP7_75t_R c8608(
.A(net7765),
.B(net7721),
.C(net8622),
.D(net8630),
.E(net8526),
.Y(net8650)
);

OA222x2_ASAP7_75t_R c8609(
.A1(net7669),
.A2(net8644),
.B1(net8643),
.B2(net8566),
.C1(net8576),
.C2(net8606),
.Y(net8651)
);

SDFHx4_ASAP7_75t_R c8610(
.D(net8548),
.SE(net7542),
.SI(net8643),
.CLK(clk),
.QN(net8652)
);

INVx1_ASAP7_75t_R c8611(
.A(net10354),
.Y(net8653)
);

NOR3xp33_ASAP7_75t_R c8612(
.A(net8267),
.B(net8581),
.C(net10115),
.Y(net8654)
);

OA21x2_ASAP7_75t_R c8613(
.A1(net8642),
.A2(net8645),
.B(net8644),
.Y(net8655)
);

SDFLx1_ASAP7_75t_R c8614(
.D(net8559),
.SE(net8652),
.SI(net7754),
.CLK(clk),
.QN(net8656)
);

OA33x2_ASAP7_75t_R c8615(
.A1(net8589),
.A2(net8656),
.A3(net8646),
.B1(net8575),
.B2(net8606),
.B3(net7759),
.Y(net8657)
);

INVx2_ASAP7_75t_R c8616(
.A(net10383),
.Y(net8658)
);

OAI21x1_ASAP7_75t_R c8617(
.A1(net8504),
.A2(net8294),
.B(net9875),
.Y(net8659)
);

OAI21xp33_ASAP7_75t_R c8618(
.A1(net8643),
.A2(net8658),
.B(net8647),
.Y(net8660)
);

OAI21xp5_ASAP7_75t_R c8619(
.A1(net8648),
.A2(net8575),
.B(net9886),
.Y(net8661)
);

OR3x1_ASAP7_75t_R c8620(
.A(net8608),
.B(net8653),
.C(net9661),
.Y(net8662)
);

OR3x2_ASAP7_75t_R c8621(
.A(net8644),
.B(net8419),
.C(net10092),
.Y(net8663)
);

OR3x4_ASAP7_75t_R c8622(
.A(net8659),
.B(net8510),
.C(net10144),
.Y(net8664)
);

AND3x1_ASAP7_75t_R c8623(
.A(net8653),
.B(net8658),
.C(net10009),
.Y(net8665)
);

SDFLx2_ASAP7_75t_R c8624(
.D(net8615),
.SE(net8611),
.SI(net8652),
.CLK(clk),
.QN(net8666)
);

AND3x2_ASAP7_75t_R c8625(
.A(net8588),
.B(net8666),
.C(net10092),
.Y(net8667)
);

SDFLx3_ASAP7_75t_R c8626(
.D(net8664),
.SE(net8636),
.SI(net8615),
.CLK(clk),
.QN(net8668)
);

AND3x4_ASAP7_75t_R c8627(
.A(net8667),
.B(net8656),
.C(net8649),
.Y(net8669)
);

AO21x1_ASAP7_75t_R c8628(
.A1(net8629),
.A2(net8579),
.B(net9942),
.Y(net8670)
);

AO21x2_ASAP7_75t_R c8629(
.A1(net8665),
.A2(net8606),
.B(net10059),
.Y(net8671)
);

ICGx3_ASAP7_75t_R c8630(
.ENA(net8581),
.SE(net8669),
.CLK(clk),
.GCLK(net8672)
);

SDFLx4_ASAP7_75t_R c8631(
.D(net8598),
.SE(net8649),
.SI(net9661),
.CLK(clk),
.QN(net8673)
);

AOI21x1_ASAP7_75t_R c8632(
.A1(net8620),
.A2(net8478),
.B(net8529),
.Y(net8674)
);

NAND2x2_ASAP7_75t_R c8633(
.A(net7708),
.B(net8583),
.Y(net8675)
);

AOI21xp33_ASAP7_75t_R c8634(
.A1(net8663),
.A2(net8620),
.B(net7839),
.Y(net8676)
);

INVx3_ASAP7_75t_R c8635(
.A(net10154),
.Y(net8677)
);

INVx4_ASAP7_75t_R c8636(
.A(net10154),
.Y(net8678)
);

NAND2xp33_ASAP7_75t_R c8637(
.A(net8595),
.B(net8420),
.Y(net8679)
);

AOI21xp5_ASAP7_75t_R c8638(
.A1(net8594),
.A2(net8460),
.B(net7846),
.Y(net8680)
);

FAx1_ASAP7_75t_R c8639(
.A(net8668),
.B(net8646),
.CI(net10132),
.SN(net8681)
);

MAJIxp5_ASAP7_75t_R c8640(
.A(net7747),
.B(net8506),
.C(net10154),
.Y(net8682)
);

NAND2xp5_ASAP7_75t_R c8641(
.A(net8569),
.B(net6925),
.Y(net8683)
);

DFFASRHQNx1_ASAP7_75t_R c8642(
.D(net7754),
.RESETN(net8632),
.SETN(net8675),
.CLK(clk),
.QN(net8684)
);

NAND2xp67_ASAP7_75t_R c8643(
.A(net8673),
.B(net6493),
.Y(net8685)
);

INVx5_ASAP7_75t_R c8644(
.A(net10518),
.Y(net8686)
);

NOR2x1_ASAP7_75t_R c8645(
.A(net8507),
.B(net8632),
.Y(net8687)
);

NOR2x1p5_ASAP7_75t_R c8646(
.A(net8593),
.B(net8587),
.Y(net8688)
);

NOR2x2_ASAP7_75t_R c8647(
.A(net6905),
.B(net8677),
.Y(net8689)
);

SDFHx1_ASAP7_75t_R c8648(
.D(net6804),
.SE(net7754),
.SI(net8688),
.CLK(clk),
.QN(net8690)
);

NOR2xp33_ASAP7_75t_R c8649(
.A(net8460),
.B(net8681),
.Y(net8691)
);

MAJx2_ASAP7_75t_R c8650(
.A(net8631),
.B(net7651),
.C(net10313),
.Y(net8692)
);

NOR2xp67_ASAP7_75t_R c8651(
.A(net7846),
.B(net6830),
.Y(net8693)
);

OR2x2_ASAP7_75t_R c8652(
.A(net7825),
.B(net8680),
.Y(net8694)
);

OR2x4_ASAP7_75t_R c8653(
.A(net7747),
.B(net6804),
.Y(net8695)
);

OR2x6_ASAP7_75t_R c8654(
.A(net7842),
.B(net8666),
.Y(net8696)
);

XNOR2x1_ASAP7_75t_R c8655(
.B(net7799),
.A(net7857),
.Y(net8697)
);

OAI31xp33_ASAP7_75t_R c8656(
.A1(net7839),
.A2(net8646),
.A3(net8684),
.B(net8506),
.Y(net8698)
);

XNOR2x2_ASAP7_75t_R c8657(
.A(net7806),
.B(net10320),
.Y(net8699)
);

MAJx3_ASAP7_75t_R c8658(
.A(net8570),
.B(net8605),
.C(net8699),
.Y(net8700)
);

XNOR2xp5_ASAP7_75t_R c8659(
.A(net8604),
.B(net10320),
.Y(net8701)
);

NAND3x1_ASAP7_75t_R c8660(
.A(net8647),
.B(net8690),
.C(net8673),
.Y(net8702)
);

NAND3x2_ASAP7_75t_R c8661(
.B(net8585),
.C(net7651),
.A(net9705),
.Y(net8703)
);

NAND3xp33_ASAP7_75t_R c8662(
.A(net8695),
.B(net7619),
.C(net10146),
.Y(net8704)
);

XOR2x1_ASAP7_75t_R c8663(
.A(net8592),
.B(net10026),
.Y(net8705)
);

NOR3x1_ASAP7_75t_R c8664(
.A(net8347),
.B(net7619),
.C(net8649),
.Y(net8706)
);

NOR3x2_ASAP7_75t_R c8665(
.B(net8693),
.C(net7830),
.A(net7799),
.Y(net8707)
);

NOR3xp33_ASAP7_75t_R c8666(
.A(net8692),
.B(net8668),
.C(net8622),
.Y(net8708)
);

OA21x2_ASAP7_75t_R c8667(
.A1(net8679),
.A2(net8706),
.B(net8675),
.Y(net8709)
);

OAI21x1_ASAP7_75t_R c8668(
.A1(net8702),
.A2(net8705),
.B(net7747),
.Y(net8710)
);

XOR2x2_ASAP7_75t_R c8669(
.A(net7658),
.B(net7764),
.Y(net8711)
);

OAI21xp33_ASAP7_75t_R c8670(
.A1(net8357),
.A2(net8507),
.B(net8512),
.Y(net8712)
);

OAI21xp5_ASAP7_75t_R c8671(
.A1(net8699),
.A2(net8621),
.B(net5105),
.Y(net8713)
);

SDFHx2_ASAP7_75t_R c8672(
.D(net8640),
.SE(net8706),
.SI(net7619),
.CLK(clk),
.QN(net8714)
);

OR3x1_ASAP7_75t_R c8673(
.A(net8531),
.B(net8695),
.C(net7799),
.Y(net8715)
);

OR3x2_ASAP7_75t_R c8674(
.A(net7651),
.B(net8366),
.C(net8690),
.Y(net8716)
);

OR3x4_ASAP7_75t_R c8675(
.A(net8604),
.B(net8682),
.C(net8695),
.Y(net8717)
);

AND3x1_ASAP7_75t_R c8676(
.A(net8711),
.B(net7754),
.C(net6016),
.Y(net8718)
);

AND3x2_ASAP7_75t_R c8677(
.A(net8696),
.B(net8347),
.C(net10313),
.Y(net8719)
);

OAI222xp33_ASAP7_75t_R c8678(
.A1(net8683),
.A2(net7619),
.B1(net7842),
.B2(net8695),
.C1(net8675),
.C2(net8666),
.Y(net8720)
);

AND3x4_ASAP7_75t_R c8679(
.A(net8704),
.B(net8715),
.C(net7839),
.Y(net8721)
);

XOR2xp5_ASAP7_75t_R c8680(
.A(net7688),
.B(net7825),
.Y(net8722)
);

AO21x1_ASAP7_75t_R c8681(
.A1(net6925),
.A2(net8717),
.B(net8640),
.Y(net8723)
);

AO21x2_ASAP7_75t_R c8682(
.A1(net8630),
.A2(net8719),
.B(net8675),
.Y(net8724)
);

SDFHx3_ASAP7_75t_R c8683(
.D(net8626),
.SE(net5105),
.SI(net8714),
.CLK(clk),
.QN(net8725)
);

AND2x2_ASAP7_75t_R c8684(
.A(net8506),
.B(net8479),
.Y(net8726)
);

AOI21x1_ASAP7_75t_R c8685(
.A1(net7764),
.A2(net8725),
.B(net10154),
.Y(net8727)
);

AOI21xp33_ASAP7_75t_R c8686(
.A1(net8605),
.A2(net8594),
.B(net9851),
.Y(net8728)
);

AOI21xp5_ASAP7_75t_R c8687(
.A1(net8727),
.A2(net8719),
.B(net8711),
.Y(net8729)
);

AND2x4_ASAP7_75t_R c8688(
.A(net9991),
.B(net10026),
.Y(net8730)
);

AND2x6_ASAP7_75t_R c8689(
.A(net7456),
.B(net8716),
.Y(net8731)
);

FAx1_ASAP7_75t_R c8690(
.A(net7830),
.B(net6947),
.CI(net7822),
.SN(net8733),
.CON(net8732)
);

MAJIxp5_ASAP7_75t_R c8691(
.A(net8731),
.B(net8729),
.C(net8715),
.Y(net8734)
);

MAJx2_ASAP7_75t_R c8692(
.A(net6599),
.B(net8494),
.C(net8658),
.Y(net8735)
);

MAJx3_ASAP7_75t_R c8693(
.A(net7862),
.B(net8678),
.C(net8606),
.Y(net8736)
);

HAxp5_ASAP7_75t_R c8694(
.A(net8734),
.B(net8512),
.CON(net8737)
);

OAI31xp67_ASAP7_75t_R c8695(
.A1(net8728),
.A2(net8686),
.A3(out13),
.B(net10132),
.Y(net8738)
);

NAND3x1_ASAP7_75t_R c8696(
.A(net8685),
.B(net8730),
.C(net8714),
.Y(net8739)
);

NAND3x2_ASAP7_75t_R c8697(
.B(net8479),
.C(net8723),
.A(net8731),
.Y(net8740)
);

NAND3xp33_ASAP7_75t_R c8698(
.A(net8712),
.B(net8739),
.C(net7830),
.Y(net8741)
);

NOR3x1_ASAP7_75t_R c8699(
.A(net8739),
.B(net8459),
.C(net7862),
.Y(net8742)
);

NOR3x2_ASAP7_75t_R c8700(
.B(net8494),
.C(net8742),
.A(net8630),
.Y(net8743)
);

NOR3xp33_ASAP7_75t_R c8701(
.A(net8741),
.B(net8699),
.C(net9974),
.Y(net8744)
);

NAND2x1_ASAP7_75t_R c8702(
.A(net8728),
.B(net8716),
.Y(net8745)
);

OR4x1_ASAP7_75t_R c8703(
.A(net6947),
.B(net8745),
.C(net8739),
.D(net8606),
.Y(net8746)
);

OA21x2_ASAP7_75t_R c8704(
.A1(net8579),
.A2(net8729),
.B(net8688),
.Y(net8747)
);

OAI21x1_ASAP7_75t_R c8705(
.A1(net8719),
.A2(net8739),
.B(net9851),
.Y(net8748)
);

OAI21xp33_ASAP7_75t_R c8706(
.A1(net8632),
.A2(net8459),
.B(net7764),
.Y(net8749)
);

NOR5xp2_ASAP7_75t_R c8707(
.A(net8701),
.B(net8740),
.C(net8732),
.D(net8585),
.E(net7826),
.Y(net8750)
);

OAI21xp5_ASAP7_75t_R c8708(
.A1(net7801),
.A2(net8730),
.B(net8725),
.Y(net8751)
);

OR4x2_ASAP7_75t_R c8709(
.A(net8726),
.B(net8742),
.C(net10025),
.D(net10321),
.Y(net8752)
);

OR3x1_ASAP7_75t_R c8710(
.A(net8609),
.B(net8715),
.C(net8745),
.Y(net8753)
);

OR3x2_ASAP7_75t_R c8711(
.A(net8752),
.B(net8749),
.C(net9915),
.Y(net8754)
);

A2O1A1Ixp33_ASAP7_75t_R c8712(
.A1(net8754),
.A2(net8745),
.B(net8587),
.C(net9974),
.Y(net8755)
);

OR3x4_ASAP7_75t_R c8713(
.A(net8723),
.B(net8725),
.C(net7651),
.Y(net8756)
);

OAI321xp33_ASAP7_75t_R c8714(
.A1(net8738),
.A2(net8756),
.A3(net8755),
.B1(net8688),
.B2(net8666),
.C(net8675),
.Y(net8757)
);

NAND2x1p5_ASAP7_75t_R c8715(
.A(net8697),
.B(net9882),
.Y(net8758)
);

AND4x1_ASAP7_75t_R c8716(
.A(net7884),
.B(net8622),
.C(net8478),
.D(net8695),
.Y(net8759)
);

NAND2x2_ASAP7_75t_R c8717(
.A(net7822),
.B(net8758),
.Y(net8760)
);

SDFHx4_ASAP7_75t_R c8718(
.D(net8575),
.SE(net8606),
.SI(net8337),
.CLK(clk),
.QN(net8761)
);

INVx6_ASAP7_75t_R c8719(
.A(net10104),
.Y(net8762)
);

AND3x1_ASAP7_75t_R c8720(
.A(net8537),
.B(net7393),
.C(net8606),
.Y(net8763)
);

SDFLx1_ASAP7_75t_R c8721(
.D(net7947),
.SE(net8755),
.SI(net8585),
.CLK(clk),
.QN(net8764)
);

NAND2xp33_ASAP7_75t_R c8722(
.A(net7935),
.B(net8420),
.Y(net8765)
);

AND3x2_ASAP7_75t_R c8723(
.A(net8587),
.B(net8672),
.C(net10001),
.Y(net8766)
);

INVx8_ASAP7_75t_R c8724(
.A(net10492),
.Y(net8767)
);

SDFLx2_ASAP7_75t_R c8725(
.D(net7885),
.SE(net6905),
.SI(net8753),
.CLK(clk),
.QN(net8768)
);

NAND2xp5_ASAP7_75t_R c8726(
.A(net8689),
.B(net8686),
.Y(net8769)
);

AND3x4_ASAP7_75t_R c8727(
.A(net8686),
.B(net7481),
.C(net9654),
.Y(net8770)
);

NAND2xp67_ASAP7_75t_R c8728(
.A(net7904),
.B(net7953),
.Y(net8771)
);

INVxp33_ASAP7_75t_R c8729(
.A(net10356),
.Y(net8772)
);

AO21x1_ASAP7_75t_R c8730(
.A1(net7873),
.A2(net7831),
.B(net8772),
.Y(net8773)
);

INVxp67_ASAP7_75t_R c8731(
.A(net10370),
.Y(net8774)
);

NOR2x1_ASAP7_75t_R c8732(
.A(net8758),
.B(net8529),
.Y(net8775)
);

NOR2x1p5_ASAP7_75t_R c8733(
.A(net8708),
.B(net7904),
.Y(net8776)
);

AO21x2_ASAP7_75t_R c8734(
.A1(net6025),
.A2(net8672),
.B(net8376),
.Y(net8777)
);

BUFx10_ASAP7_75t_R c8735(
.A(net10347),
.Y(net8778)
);

NOR2x2_ASAP7_75t_R c8736(
.A(net6016),
.B(net8691),
.Y(net8779)
);

OAI33xp33_ASAP7_75t_R c8737(
.A1(net7019),
.A2(net7820),
.A3(net8745),
.B1(net8315),
.B2(net8695),
.B3(net8675),
.Y(net8780)
);

AOI21x1_ASAP7_75t_R c8738(
.A1(net8762),
.A2(net3272),
.B(net8758),
.Y(net8781)
);

AOI21xp33_ASAP7_75t_R c8739(
.A1(net8742),
.A2(net7884),
.B(net10319),
.Y(net8782)
);

AOI21xp5_ASAP7_75t_R c8740(
.A1(net8621),
.A2(net8767),
.B(net8781),
.Y(net8783)
);

NOR2xp33_ASAP7_75t_R c8741(
.A(net8760),
.B(net8774),
.Y(net8784)
);

FAx1_ASAP7_75t_R c8742(
.A(net6917),
.B(net8697),
.CI(net8772),
.SN(net8786),
.CON(net8785)
);

MAJIxp5_ASAP7_75t_R c8743(
.A(net8770),
.B(net8622),
.C(net7822),
.Y(net8787)
);

MAJx2_ASAP7_75t_R c8744(
.A(net7769),
.B(net6917),
.C(net8733),
.Y(net8788)
);

MAJx3_ASAP7_75t_R c8745(
.A(net6099),
.B(net8772),
.C(net8427),
.Y(net8789)
);

SDFLx3_ASAP7_75t_R c8746(
.D(net8337),
.SE(net7759),
.SI(net7769),
.CLK(clk),
.QN(net8790)
);

NOR2xp67_ASAP7_75t_R c8747(
.A(net8753),
.B(net10303),
.Y(net8791)
);

SDFLx4_ASAP7_75t_R c8748(
.D(net8737),
.SE(net8786),
.SI(net6099),
.CLK(clk),
.QN(net8792)
);

NAND3x1_ASAP7_75t_R c8749(
.A(net8733),
.B(net8585),
.C(net7953),
.Y(net8793)
);

DFFASRHQNx1_ASAP7_75t_R c8750(
.D(net3272),
.RESETN(net8778),
.SETN(net8585),
.CLK(clk),
.QN(net8794)
);

NAND3x2_ASAP7_75t_R c8751(
.B(net6795),
.C(net8666),
.A(net8774),
.Y(net8795)
);

NAND3xp33_ASAP7_75t_R c8752(
.A(net8785),
.B(net8765),
.C(net9903),
.Y(net8796)
);

NOR3x1_ASAP7_75t_R c8753(
.A(net8605),
.B(net8768),
.C(net8675),
.Y(net8797)
);

BUFx12_ASAP7_75t_R c8754(
.A(net10377),
.Y(net8798)
);

OR2x2_ASAP7_75t_R c8755(
.A(net8687),
.B(net8776),
.Y(net8799)
);

NOR3x2_ASAP7_75t_R c8756(
.B(net8790),
.C(net8742),
.A(net8767),
.Y(net8800)
);

NOR3xp33_ASAP7_75t_R c8757(
.A(net7820),
.B(net8761),
.C(net8785),
.Y(net8801)
);

AND4x2_ASAP7_75t_R c8758(
.A(net8798),
.B(net8799),
.C(net6905),
.D(net10322),
.Y(net8802)
);

OA21x2_ASAP7_75t_R c8759(
.A1(net8791),
.A2(net8665),
.B(net9959),
.Y(net8803)
);

BUFx12f_ASAP7_75t_R c8760(
.A(net10347),
.Y(net8804)
);

OAI21x1_ASAP7_75t_R c8761(
.A1(net8778),
.A2(net8795),
.B(net8784),
.Y(net8805)
);

AO211x2_ASAP7_75t_R c8762(
.A1(net8716),
.A2(net8804),
.B(net8790),
.C(net7014),
.Y(net8806)
);

SDFHx1_ASAP7_75t_R c8763(
.D(net7831),
.SE(net8537),
.SI(net8801),
.CLK(clk),
.QN(net8807)
);

SDFHx2_ASAP7_75t_R c8764(
.D(net8505),
.SE(net8691),
.SI(net8606),
.CLK(clk),
.QN(net8808)
);

OR2x4_ASAP7_75t_R c8765(
.A(net8784),
.B(net8575),
.Y(net8809)
);

OAI21xp33_ASAP7_75t_R c8766(
.A1(net8799),
.A2(net8805),
.B(net6795),
.Y(net8810)
);

OAI21xp5_ASAP7_75t_R c8767(
.A1(net8583),
.A2(net8805),
.B(net9915),
.Y(net8811)
);

OA221x2_ASAP7_75t_R c8768(
.A1(net8675),
.A2(net8783),
.B1(net8478),
.B2(net7831),
.C(net10323),
.Y(net8812)
);

OR3x1_ASAP7_75t_R c8769(
.A(net8587),
.B(net8801),
.C(net10323),
.Y(net8813)
);

OR2x6_ASAP7_75t_R c8770(
.A(net8807),
.B(net10140),
.Y(net8814)
);

OR3x2_ASAP7_75t_R c8771(
.A(net8801),
.B(net8794),
.C(net7574),
.Y(net8815)
);

XNOR2x1_ASAP7_75t_R c8772(
.B(net8781),
.A(net9989),
.Y(net8816)
);

AO22x1_ASAP7_75t_R c8773(
.A1(net7466),
.A2(net8794),
.B1(net7822),
.B2(net10323),
.Y(net8817)
);

AO22x2_ASAP7_75t_R c8774(
.A1(net8714),
.A2(net8817),
.B1(net9875),
.B2(net10323),
.Y(net8818)
);

XNOR2x2_ASAP7_75t_R c8775(
.A(net8741),
.B(net8553),
.Y(net8819)
);

SDFHx3_ASAP7_75t_R c8776(
.D(net8813),
.SE(net8818),
.SI(net8801),
.CLK(clk),
.QN(net8820)
);

XNOR2xp5_ASAP7_75t_R c8777(
.A(net8815),
.B(net8816),
.Y(net8821)
);

AO31x2_ASAP7_75t_R c8778(
.A1(net8814),
.A2(net8807),
.A3(net3969),
.B(net8816),
.Y(net8822)
);

OAI221xp5_ASAP7_75t_R c8779(
.A1(net8748),
.A2(net8684),
.B1(net8751),
.B2(net7667),
.C(net8816),
.Y(net8823)
);

XOR2x1_ASAP7_75t_R c8780(
.A(net8665),
.B(net8505),
.Y(net8824)
);

OAI311xp33_ASAP7_75t_R c8781(
.A1(net8800),
.A2(net8818),
.A3(net8774),
.B1(net8675),
.C1(net10323),
.Y(net8825)
);

OR3x4_ASAP7_75t_R c8782(
.A(net8811),
.B(net8585),
.C(net8622),
.Y(net8826)
);

AND3x1_ASAP7_75t_R c8783(
.A(net8807),
.B(net8821),
.C(net6643),
.Y(net8827)
);

AND3x2_ASAP7_75t_R c8784(
.A(net8748),
.B(net9990),
.C(net10323),
.Y(net8828)
);

AND3x4_ASAP7_75t_R c8785(
.A(net7936),
.B(net8822),
.C(net6099),
.Y(net8829)
);

AOI211x1_ASAP7_75t_R c8786(
.A1(net8796),
.A2(net8828),
.B(net8794),
.C(net10323),
.Y(net8830)
);

AO21x1_ASAP7_75t_R c8787(
.A1(net8794),
.A2(net8741),
.B(net9988),
.Y(net8831)
);

SDFHx4_ASAP7_75t_R c8788(
.D(net8700),
.SE(net8427),
.SI(net8830),
.CLK(clk),
.QN(net8832)
);

XOR2x2_ASAP7_75t_R c8789(
.A(net8782),
.B(net8823),
.Y(net8833)
);

OAI32xp33_ASAP7_75t_R c8790(
.A1(net8833),
.A2(net8684),
.A3(net8804),
.B1(net8587),
.B2(net8675),
.Y(net8834)
);

SDFLx1_ASAP7_75t_R c8791(
.D(net8831),
.SE(net8818),
.SI(net9997),
.CLK(clk),
.QN(net8835)
);

AO21x2_ASAP7_75t_R c8792(
.A1(net8830),
.A2(net8828),
.B(net10032),
.Y(net8836)
);

AOI21x1_ASAP7_75t_R c8793(
.A1(net8529),
.A2(net8827),
.B(net8828),
.Y(net8837)
);

AOI21xp33_ASAP7_75t_R c8794(
.A1(net8821),
.A2(net8832),
.B(net8816),
.Y(net8838)
);

AOI21xp5_ASAP7_75t_R c8795(
.A1(net8838),
.A2(net8832),
.B(net9819),
.Y(net8839)
);

SDFLx2_ASAP7_75t_R c8796(
.D(net8688),
.SE(net8835),
.SI(net9787),
.CLK(clk),
.QN(net8840)
);

SDFLx3_ASAP7_75t_R c8797(
.D(net8835),
.SE(net8831),
.SI(net9928),
.CLK(clk),
.QN(net8841)
);

XOR2xp5_ASAP7_75t_R c8798(
.A(net7975),
.B(net8016),
.Y(net8842)
);

FAx1_ASAP7_75t_R c8799(
.A(net8820),
.B(net6519),
.CI(net10321),
.SN(net8844),
.CON(net8843)
);

AND2x2_ASAP7_75t_R c8800(
.A(net8583),
.B(net10322),
.Y(net8845)
);

AND2x4_ASAP7_75t_R c8801(
.A(net4307),
.B(net8661),
.Y(net8846)
);

MAJIxp5_ASAP7_75t_R c8802(
.A(net8773),
.B(net9654),
.C(net10323),
.Y(net8847)
);

BUFx16f_ASAP7_75t_R c8803(
.A(net10424),
.Y(net8848)
);

AND2x6_ASAP7_75t_R c8804(
.A(net8769),
.B(net8806),
.Y(net8849)
);

HAxp5_ASAP7_75t_R c8805(
.A(net10151),
.B(net10323),
.CON(net8850)
);

BUFx24_ASAP7_75t_R c8806(
.A(net10334),
.Y(net8851)
);

OR5x1_ASAP7_75t_R c8807(
.A(net8846),
.B(net7956),
.C(net8016),
.D(net8806),
.E(net8666),
.Y(net8852)
);

NAND2x1_ASAP7_75t_R c8808(
.A(net7826),
.B(net8576),
.Y(net8853)
);

MAJx2_ASAP7_75t_R c8809(
.A(net7789),
.B(net8376),
.C(net8820),
.Y(net8854)
);

MAJx3_ASAP7_75t_R c8810(
.A(net8842),
.B(net8661),
.C(net8764),
.Y(net8855)
);

NAND3x1_ASAP7_75t_R c8811(
.A(net8847),
.B(net8576),
.C(net7921),
.Y(net8856)
);

NAND2x1p5_ASAP7_75t_R c8812(
.A(net4962),
.B(net8844),
.Y(net8857)
);

ICGx4DC_ASAP7_75t_R c8813(
.ENA(net8566),
.SE(net8011),
.CLK(clk),
.GCLK(net8858)
);

BUFx2_ASAP7_75t_R c8814(
.A(net10094),
.Y(net8859)
);

AOI211xp5_ASAP7_75t_R c8815(
.A1(net7046),
.A2(net7116),
.B(net7953),
.C(net8855),
.Y(net8860)
);

AOI22x1_ASAP7_75t_R c8816(
.A1(net5971),
.A2(net7943),
.B1(net8792),
.B2(net8427),
.Y(net8861)
);

SDFLx4_ASAP7_75t_R c8817(
.D(net7759),
.SE(net6643),
.SI(net8855),
.CLK(clk),
.QN(net8862)
);

NAND3x2_ASAP7_75t_R c8818(
.B(net7477),
.C(net8855),
.A(net10321),
.Y(net8863)
);

NAND3xp33_ASAP7_75t_R c8819(
.A(net7988),
.B(out13),
.C(net8816),
.Y(net8864)
);

NOR3x1_ASAP7_75t_R c8820(
.A(net8749),
.B(net8672),
.C(net8847),
.Y(net8865)
);

NOR3x2_ASAP7_75t_R c8821(
.B(net8864),
.C(net8714),
.A(net8788),
.Y(net8866)
);

NOR3xp33_ASAP7_75t_R c8822(
.A(net8777),
.B(net10140),
.C(net10324),
.Y(net8867)
);

OA21x2_ASAP7_75t_R c8823(
.A1(net8011),
.A2(net8847),
.B(net8783),
.Y(net8868)
);

NAND2x2_ASAP7_75t_R c8824(
.A(net8861),
.B(net8859),
.Y(net8869)
);

OAI21x1_ASAP7_75t_R c8825(
.A1(net8765),
.A2(net6852),
.B(net10307),
.Y(net8870)
);

OAI21xp33_ASAP7_75t_R c8826(
.A1(net8859),
.A2(net8646),
.B(net8817),
.Y(net8871)
);

OAI21xp5_ASAP7_75t_R c8827(
.A1(net8787),
.A2(net8848),
.B(net7116),
.Y(net8872)
);

NAND2xp33_ASAP7_75t_R c8828(
.A(net8661),
.B(net8871),
.Y(net8873)
);

NAND2xp5_ASAP7_75t_R c8829(
.A(net8869),
.B(net8866),
.Y(net8874)
);

NAND2xp67_ASAP7_75t_R c8830(
.A(net8868),
.B(net8749),
.Y(net8875)
);

OR5x2_ASAP7_75t_R c8831(
.A(net8516),
.B(net8862),
.C(net8576),
.D(net7759),
.E(net7054),
.Y(net8876)
);

ICGx4_ASAP7_75t_R c8832(
.ENA(net8819),
.SE(net8853),
.CLK(clk),
.GCLK(net8877)
);

OR3x1_ASAP7_75t_R c8833(
.A(net8816),
.B(net7069),
.C(net8646),
.Y(net8878)
);

NOR2x1_ASAP7_75t_R c8834(
.A(net8745),
.B(net8868),
.Y(net8879)
);

OR3x2_ASAP7_75t_R c8835(
.A(net7116),
.B(net9787),
.C(net9913),
.Y(net8880)
);

BUFx3_ASAP7_75t_R c8836(
.A(net10424),
.Y(net8881)
);

DFFASRHQNx1_ASAP7_75t_R c8837(
.D(net7090),
.RESETN(net8787),
.SETN(net8516),
.CLK(clk),
.QN(net8882)
);

OR3x4_ASAP7_75t_R c8838(
.A(net8877),
.B(net8847),
.C(net8010),
.Y(net8883)
);

ICGx5_ASAP7_75t_R c8839(
.ENA(net7116),
.SE(net8875),
.CLK(clk),
.GCLK(net8884)
);

NOR2x1p5_ASAP7_75t_R c8840(
.A(net8376),
.B(net8873),
.Y(net8885)
);

AND3x1_ASAP7_75t_R c8841(
.A(net8010),
.B(net8478),
.C(net7943),
.Y(net8886)
);

AND3x2_ASAP7_75t_R c8842(
.A(net8878),
.B(net7014),
.C(net10307),
.Y(net8887)
);

NOR2x2_ASAP7_75t_R c8843(
.A(net7972),
.B(net8881),
.Y(net8888)
);

BUFx4_ASAP7_75t_R c8844(
.A(net10451),
.Y(net8889)
);

AND3x4_ASAP7_75t_R c8845(
.A(net7014),
.B(out13),
.C(net10029),
.Y(net8890)
);

AO21x1_ASAP7_75t_R c8846(
.A1(net8845),
.A2(net8882),
.B(net10057),
.Y(net8891)
);

BUFx4f_ASAP7_75t_R c8847(
.A(net10351),
.Y(net8892)
);

AO21x2_ASAP7_75t_R c8848(
.A1(net8768),
.A2(net8865),
.B(net10325),
.Y(net8893)
);

AOI21x1_ASAP7_75t_R c8849(
.A1(net8006),
.A2(net8890),
.B(net8806),
.Y(net8894)
);

AOI21xp33_ASAP7_75t_R c8850(
.A1(net8849),
.A2(net7090),
.B(net9761),
.Y(net8895)
);

AOI21xp5_ASAP7_75t_R c8851(
.A1(net8016),
.A2(net8862),
.B(net8776),
.Y(net8896)
);

FAx1_ASAP7_75t_R c8852(
.A(net8788),
.B(net8749),
.CI(net10325),
.SN(net8898),
.CON(net8897)
);

NOR2xp33_ASAP7_75t_R c8853(
.A(net8863),
.B(net8576),
.Y(net8899)
);

MAJIxp5_ASAP7_75t_R c8854(
.A(net8887),
.B(net7061),
.C(net8376),
.Y(net8900)
);

MAJx2_ASAP7_75t_R c8855(
.A(net8710),
.B(net8783),
.C(net8777),
.Y(net8901)
);

MAJx3_ASAP7_75t_R c8856(
.A(net8868),
.B(net7789),
.C(net9639),
.Y(net8902)
);

NAND3x1_ASAP7_75t_R c8857(
.A(net8866),
.B(net8882),
.C(net9903),
.Y(net8903)
);

NOR2xp67_ASAP7_75t_R c8858(
.A(net7953),
.B(net8786),
.Y(net8904)
);

NAND3x2_ASAP7_75t_R c8859(
.B(net7667),
.C(net8898),
.A(net8843),
.Y(net8905)
);

SDFHx1_ASAP7_75t_R c8860(
.D(net8892),
.SE(net8879),
.SI(net8865),
.CLK(clk),
.QN(net8906)
);

OR2x2_ASAP7_75t_R c8861(
.A(net8885),
.B(net8906),
.Y(net8907)
);

NAND3xp33_ASAP7_75t_R c8862(
.A(net8899),
.B(net8898),
.C(net10322),
.Y(net8908)
);

BUFx5_ASAP7_75t_R c8863(
.A(net10334),
.Y(net8909)
);

NOR3x1_ASAP7_75t_R c8864(
.A(net8891),
.B(net8907),
.C(net8858),
.Y(net8910)
);

NOR3x2_ASAP7_75t_R c8865(
.B(net8910),
.C(net8907),
.A(net8877),
.Y(net8911)
);

NOR3xp33_ASAP7_75t_R c8866(
.A(net8882),
.B(net9760),
.C(net10018),
.Y(net8912)
);

AO222x2_ASAP7_75t_R c8867(
.A1(net8870),
.A2(net8866),
.B1(net8666),
.B2(net8893),
.C1(net7956),
.C2(net8906),
.Y(net8913)
);

OA21x2_ASAP7_75t_R c8868(
.A1(net7962),
.A2(net8911),
.B(net8909),
.Y(net8914)
);

OAI21x1_ASAP7_75t_R c8869(
.A1(net8914),
.A2(net8909),
.B(net9960),
.Y(net8915)
);

OAI21xp33_ASAP7_75t_R c8870(
.A1(net8896),
.A2(net8890),
.B(net8010),
.Y(net8916)
);

OAI21xp5_ASAP7_75t_R c8871(
.A1(net8881),
.A2(net8914),
.B(net10303),
.Y(net8917)
);

OR2x4_ASAP7_75t_R c8872(
.A(net8909),
.B(net10049),
.Y(net8918)
);

OR3x1_ASAP7_75t_R c8873(
.A(net7026),
.B(net8850),
.C(net8772),
.Y(net8919)
);

OR2x6_ASAP7_75t_R c8874(
.A(net8772),
.B(net10324),
.Y(net8920)
);

AO33x2_ASAP7_75t_R c8875(
.A1(net8919),
.A2(net8920),
.A3(net8658),
.B1(net8893),
.B2(net8914),
.B3(net10322),
.Y(net8921)
);

OR3x2_ASAP7_75t_R c8876(
.A(net8884),
.B(net9902),
.C(net10004),
.Y(net8922)
);

OR3x4_ASAP7_75t_R c8877(
.A(net8922),
.B(net10057),
.C(net10321),
.Y(net8923)
);

AND3x1_ASAP7_75t_R c8878(
.A(net8918),
.B(net10025),
.C(net10326),
.Y(net8924)
);

AND3x2_ASAP7_75t_R c8879(
.A(net8923),
.B(net8924),
.C(net8695),
.Y(net8925)
);

A2O1A1O1Ixp25_ASAP7_75t_R c8880(
.A1(net8894),
.A2(net8887),
.B(net8925),
.C(net6132),
.D(net10326),
.Y(net8926)
);

XNOR2x1_ASAP7_75t_R c8881(
.B(net8315),
.A(net8884),
.Y(net8927)
);

AND3x4_ASAP7_75t_R c8882(
.A(net8909),
.B(net8755),
.C(net8889),
.Y(net8928)
);

AOI22xp33_ASAP7_75t_R c8883(
.A1(net7874),
.A2(net8121),
.B1(net8607),
.B2(net10308),
.Y(net8929)
);

AO21x1_ASAP7_75t_R c8884(
.A1(net8902),
.A2(net8777),
.B(net8607),
.Y(net8930)
);

AND5x1_ASAP7_75t_R c8885(
.A(net8764),
.B(net8879),
.C(net6132),
.D(net8855),
.E(net8909),
.Y(net8931)
);

AO21x2_ASAP7_75t_R c8886(
.A1(net7069),
.A2(net7026),
.B(net7124),
.Y(net8932)
);

XNOR2x2_ASAP7_75t_R c8887(
.A(net8880),
.B(net10125),
.Y(net8933)
);

XNOR2xp5_ASAP7_75t_R c8888(
.A(net8895),
.B(net7163),
.Y(net8934)
);

SDFHx2_ASAP7_75t_R c8889(
.D(net8718),
.SE(net9819),
.SI(net10055),
.CLK(clk),
.QN(net8935)
);

XOR2x1_ASAP7_75t_R c8890(
.A(net6830),
.B(net8933),
.Y(net8936)
);

AOI21x1_ASAP7_75t_R c8891(
.A1(net6852),
.A2(net8855),
.B(net8775),
.Y(net8937)
);

BUFx6f_ASAP7_75t_R c8892(
.A(net10335),
.Y(net8938)
);

SDFHx3_ASAP7_75t_R c8893(
.D(net8809),
.SE(net8914),
.SI(net9995),
.CLK(clk),
.QN(net8939)
);

SDFHx4_ASAP7_75t_R c8894(
.D(net8478),
.SE(net8806),
.SI(net10125),
.CLK(clk),
.QN(net8940)
);

AOI21xp33_ASAP7_75t_R c8895(
.A1(net8792),
.A2(net8940),
.B(net10140),
.Y(net8941)
);

XOR2x2_ASAP7_75t_R c8896(
.A(net6129),
.B(net8909),
.Y(net8942)
);

AOI21xp5_ASAP7_75t_R c8897(
.A1(net7054),
.A2(net8841),
.B(net10321),
.Y(net8943)
);

XOR2xp5_ASAP7_75t_R c8898(
.A(net8933),
.B(net10151),
.Y(net8944)
);

FAx1_ASAP7_75t_R c8899(
.A(net5311),
.B(net8933),
.CI(net8806),
.SN(net8945)
);

BUFx8_ASAP7_75t_R c8900(
.A(net10374),
.Y(net8946)
);

AND2x2_ASAP7_75t_R c8901(
.A(net8929),
.B(net8933),
.Y(net8947)
);

MAJIxp5_ASAP7_75t_R c8902(
.A(net8777),
.B(net7899),
.C(net8946),
.Y(net8948)
);

AND2x4_ASAP7_75t_R c8903(
.A(net8607),
.B(net7959),
.Y(net8949)
);

AND2x6_ASAP7_75t_R c8904(
.A(net7061),
.B(net7069),
.Y(net8950)
);

MAJx2_ASAP7_75t_R c8905(
.A(net7146),
.B(net8938),
.C(net8909),
.Y(net8951)
);

CKINVDCx10_ASAP7_75t_R c8906(
.A(net10335),
.Y(net8952)
);

AOI22xp5_ASAP7_75t_R c8907(
.A1(net8951),
.A2(net8666),
.B1(net8048),
.B2(net8939),
.Y(net8953)
);

MAJx3_ASAP7_75t_R c8908(
.A(net8895),
.B(net8764),
.C(net10325),
.Y(net8954)
);

AOI31xp33_ASAP7_75t_R c8909(
.A1(net8828),
.A2(net8935),
.A3(net8120),
.B(net8427),
.Y(net8955)
);

NAND3x1_ASAP7_75t_R c8910(
.A(net4363),
.B(net7786),
.C(net8048),
.Y(net8956)
);

NAND3x2_ASAP7_75t_R c8911(
.B(net8889),
.C(net8933),
.A(net8935),
.Y(net8957)
);

NAND3xp33_ASAP7_75t_R c8912(
.A(net8048),
.B(net8955),
.C(net8951),
.Y(net8958)
);

NOR3x1_ASAP7_75t_R c8913(
.A(net8952),
.B(net1652),
.C(net9877),
.Y(net8959)
);

AOI31xp67_ASAP7_75t_R c8914(
.A1(net5294),
.A2(net8858),
.A3(net8315),
.B(net9998),
.Y(net8960)
);

NOR3x2_ASAP7_75t_R c8915(
.B(net8882),
.C(net8946),
.A(net8607),
.Y(net8961)
);

NOR3xp33_ASAP7_75t_R c8916(
.A(net8952),
.B(net8658),
.C(net8934),
.Y(net8962)
);

OA21x2_ASAP7_75t_R c8917(
.A1(net8764),
.A2(net7054),
.B(net10125),
.Y(net8963)
);

HAxp5_ASAP7_75t_R c8918(
.A(net8961),
.B(net9687),
.CON(net8964)
);

OAI21x1_ASAP7_75t_R c8919(
.A1(net8946),
.A2(net7054),
.B(net10159),
.Y(net8965)
);

OAI21xp33_ASAP7_75t_R c8920(
.A1(net8852),
.A2(net8949),
.B(net8420),
.Y(net8966)
);

OAI21xp5_ASAP7_75t_R c8921(
.A1(net7206),
.A2(net8806),
.B(net3432),
.Y(net8967)
);

OR3x1_ASAP7_75t_R c8922(
.A(net8962),
.B(net8963),
.C(net8882),
.Y(net8968)
);

OR3x2_ASAP7_75t_R c8923(
.A(net8967),
.B(net8646),
.C(net8817),
.Y(net8969)
);

OR3x4_ASAP7_75t_R c8924(
.A(net8884),
.B(net8117),
.C(net8939),
.Y(net8970)
);

AND3x1_ASAP7_75t_R c8925(
.A(net8934),
.B(net8056),
.C(net10319),
.Y(net8971)
);

AND3x2_ASAP7_75t_R c8926(
.A(net8658),
.B(net8968),
.C(net8808),
.Y(net8972)
);

AND3x4_ASAP7_75t_R c8927(
.A(net7899),
.B(net8048),
.C(net9919),
.Y(net8973)
);

AO21x1_ASAP7_75t_R c8928(
.A1(net8072),
.A2(net7574),
.B(net8960),
.Y(net8974)
);

AO21x2_ASAP7_75t_R c8929(
.A1(net7160),
.A2(net8925),
.B(net8852),
.Y(net8975)
);

NAND4xp25_ASAP7_75t_R c8930(
.A(net8947),
.B(net8944),
.C(net8975),
.D(net10321),
.Y(net8976)
);

SDFLx1_ASAP7_75t_R c8931(
.D(net8954),
.SE(net8953),
.SI(net8960),
.CLK(clk),
.QN(net8977)
);

AOI21x1_ASAP7_75t_R c8932(
.A1(net8957),
.A2(net8973),
.B(net8828),
.Y(net8978)
);

AOI21xp33_ASAP7_75t_R c8933(
.A1(net8974),
.A2(net8945),
.B(net8893),
.Y(net8979)
);

AOI21xp5_ASAP7_75t_R c8934(
.A1(net8912),
.A2(net10159),
.B(net10327),
.Y(net8980)
);

FAx1_ASAP7_75t_R c8935(
.A(net7959),
.B(net8882),
.CI(net10098),
.SN(net8981)
);

MAJIxp5_ASAP7_75t_R c8936(
.A(net8880),
.B(net8946),
.C(net8828),
.Y(net8982)
);

MAJx2_ASAP7_75t_R c8937(
.A(net7164),
.B(net8977),
.C(net10327),
.Y(net8983)
);

NAND2x1_ASAP7_75t_R c8938(
.A(net7990),
.B(net8965),
.Y(net8984)
);

MAJx3_ASAP7_75t_R c8939(
.A(net8973),
.B(net8942),
.C(net8975),
.Y(net8985)
);

NAND2x1p5_ASAP7_75t_R c8940(
.A(net8950),
.B(net10321),
.Y(net8986)
);

NAND3x1_ASAP7_75t_R c8941(
.A(net8966),
.B(net8964),
.C(net8895),
.Y(net8987)
);

NAND3x2_ASAP7_75t_R c8942(
.B(net8984),
.C(net8975),
.A(net10327),
.Y(net8988)
);

NAND3xp33_ASAP7_75t_R c8943(
.A(net6132),
.B(net7145),
.C(net8884),
.Y(net8989)
);

NOR3x1_ASAP7_75t_R c8944(
.A(net3432),
.B(net5294),
.C(net8968),
.Y(net8990)
);

NOR3x2_ASAP7_75t_R c8945(
.B(net8986),
.C(net8970),
.A(net8046),
.Y(net8991)
);

NOR3xp33_ASAP7_75t_R c8946(
.A(net8969),
.B(net7165),
.C(net3442),
.Y(net8992)
);

CKINVDCx11_ASAP7_75t_R c8947(
.A(net10351),
.Y(net8993)
);

OA21x2_ASAP7_75t_R c8948(
.A1(net8983),
.A2(net8914),
.B(net10125),
.Y(net8994)
);

OAI21x1_ASAP7_75t_R c8949(
.A1(net8714),
.A2(net8809),
.B(net8056),
.Y(net8995)
);

OAI21xp33_ASAP7_75t_R c8950(
.A1(net8989),
.A2(net8959),
.B(net8960),
.Y(net8996)
);

OAI21xp5_ASAP7_75t_R c8951(
.A1(net8968),
.A2(net8940),
.B(net10141),
.Y(net8997)
);

OR3x1_ASAP7_75t_R c8952(
.A(net8997),
.B(net8934),
.C(net10033),
.Y(net8998)
);

AOI222xp33_ASAP7_75t_R c8953(
.A1(net8943),
.A2(net8990),
.B1(net8968),
.B2(net8056),
.C1(net7054),
.C2(net8851),
.Y(net8999)
);

OR3x2_ASAP7_75t_R c8954(
.A(net8858),
.B(net8972),
.C(net8968),
.Y(net9000)
);

AND5x2_ASAP7_75t_R c8955(
.A(net8971),
.B(net8056),
.C(net8975),
.D(net7054),
.E(net10328),
.Y(net9001)
);

OR3x4_ASAP7_75t_R c8956(
.A(net8992),
.B(net7054),
.C(net10043),
.Y(net9002)
);

AND3x1_ASAP7_75t_R c8957(
.A(net8980),
.B(net8996),
.C(net10325),
.Y(net9003)
);

AND3x2_ASAP7_75t_R c8958(
.A(net7956),
.B(net8995),
.C(net10328),
.Y(net9004)
);

AND3x4_ASAP7_75t_R c8959(
.A(net8969),
.B(net10058),
.C(net10319),
.Y(net9005)
);

AOI321xp33_ASAP7_75t_R c8960(
.A1(net8992),
.A2(net8984),
.A3(net9005),
.B1(net8960),
.B2(net8952),
.C(net10046),
.Y(net9006)
);

AO21x1_ASAP7_75t_R c8961(
.A1(net8069),
.A2(net9003),
.B(net8977),
.Y(net9007)
);

AO21x2_ASAP7_75t_R c8962(
.A1(net8982),
.A2(net9005),
.B(net9906),
.Y(net9008)
);

AO221x1_ASAP7_75t_R c8963(
.A1(net8934),
.A2(net9005),
.B1(net8975),
.B2(net10037),
.C(net10141),
.Y(net9009)
);

AOI21x1_ASAP7_75t_R c8964(
.A1(net8914),
.A2(net6830),
.B(net8940),
.Y(net9010)
);

AOI21xp33_ASAP7_75t_R c8965(
.A1(net7874),
.A2(net8154),
.B(net8427),
.Y(net9011)
);

NAND2x2_ASAP7_75t_R c8966(
.A(net7178),
.B(net7868),
.Y(net9012)
);

AOI21xp5_ASAP7_75t_R c8967(
.A1(net6975),
.A2(net8940),
.B(net8975),
.Y(net9013)
);

NAND2xp33_ASAP7_75t_R c8968(
.A(net8857),
.B(net8126),
.Y(net9014)
);

CKINVDCx12_ASAP7_75t_R c8969(
.A(net10336),
.Y(net9015)
);

FAx1_ASAP7_75t_R c8970(
.A(net9012),
.B(net6214),
.CI(net8960),
.SN(net9016)
);

SDFLx2_ASAP7_75t_R c8971(
.D(net8427),
.SE(net8154),
.SI(net9687),
.CLK(clk),
.QN(net9017)
);

MAJIxp5_ASAP7_75t_R c8972(
.A(net8840),
.B(net8941),
.C(net9919),
.Y(net9018)
);

NAND2xp5_ASAP7_75t_R c8973(
.A(net2642),
.B(net9995),
.Y(net9019)
);

MAJx2_ASAP7_75t_R c8974(
.A(net8808),
.B(net7124),
.C(net7868),
.Y(net9020)
);

MAJx3_ASAP7_75t_R c8975(
.A(net9014),
.B(net7247),
.C(net8939),
.Y(net9021)
);

NAND2xp67_ASAP7_75t_R c8976(
.A(net8121),
.B(net10307),
.Y(net9022)
);

NOR2x1_ASAP7_75t_R c8977(
.A(net8166),
.B(net9998),
.Y(net9023)
);

NAND3x1_ASAP7_75t_R c8978(
.A(net8893),
.B(net9990),
.C(net10288),
.Y(net9024)
);

NAND3x2_ASAP7_75t_R c8979(
.B(net8055),
.C(net8880),
.A(net8893),
.Y(net9025)
);

CKINVDCx14_ASAP7_75t_R c8980(
.A(net10336),
.Y(net9026)
);

NAND3xp33_ASAP7_75t_R c8981(
.A(net8126),
.B(net8203),
.C(net9017),
.Y(net9027)
);

NOR3x1_ASAP7_75t_R c8982(
.A(net7982),
.B(net8817),
.C(net8975),
.Y(net9028)
);

NOR3x2_ASAP7_75t_R c8983(
.B(net8817),
.C(net7826),
.A(net8939),
.Y(net9029)
);

NOR3xp33_ASAP7_75t_R c8984(
.A(net8186),
.B(net8927),
.C(net8888),
.Y(net9030)
);

OA21x2_ASAP7_75t_R c8985(
.A1(net8193),
.A2(net8944),
.B(net9925),
.Y(net9031)
);

NOR2x1p5_ASAP7_75t_R c8986(
.A(net8893),
.B(net9031),
.Y(net9032)
);

NAND4xp75_ASAP7_75t_R c8987(
.A(net8772),
.B(net8914),
.C(net8927),
.D(net8148),
.Y(net9033)
);

NOR2x2_ASAP7_75t_R c8988(
.A(net8121),
.B(net10060),
.Y(net9034)
);

OAI21x1_ASAP7_75t_R c8989(
.A1(net7279),
.A2(net8199),
.B(net9924),
.Y(net9035)
);

OAI21xp33_ASAP7_75t_R c8990(
.A1(net8139),
.A2(net9017),
.B(net9026),
.Y(net9036)
);

SDFLx3_ASAP7_75t_R c8991(
.D(net3442),
.SE(net8154),
.SI(net9026),
.CLK(clk),
.QN(net9037)
);

OAI21xp5_ASAP7_75t_R c8992(
.A1(net6154),
.A2(net8927),
.B(net10037),
.Y(net9038)
);

OR3x1_ASAP7_75t_R c8993(
.A(net6293),
.B(net9035),
.C(net9037),
.Y(net9039)
);

OR3x2_ASAP7_75t_R c8994(
.A(net8420),
.B(net9029),
.C(net8148),
.Y(net9040)
);

OR3x4_ASAP7_75t_R c8995(
.A(net9021),
.B(net9017),
.C(net10074),
.Y(net9041)
);

AND3x1_ASAP7_75t_R c8996(
.A(net8775),
.B(net8893),
.C(net10121),
.Y(net9042)
);

NOR4xp25_ASAP7_75t_R c8997(
.A(net8975),
.B(net8198),
.C(net9017),
.D(net7124),
.Y(net9043)
);

AND3x2_ASAP7_75t_R c8998(
.A(net8046),
.B(net9022),
.C(net8148),
.Y(net9044)
);

AND3x4_ASAP7_75t_R c8999(
.A(net8925),
.B(net7982),
.C(net9743),
.Y(net9045)
);

AO21x1_ASAP7_75t_R c9000(
.A1(net9040),
.A2(net8939),
.B(net8888),
.Y(net9046)
);

AO21x2_ASAP7_75t_R c9001(
.A1(net8744),
.A2(net9023),
.B(net8817),
.Y(net9047)
);

AOI21x1_ASAP7_75t_R c9002(
.A1(net8120),
.A2(net8944),
.B(out15),
.Y(net9048)
);

AOI21xp33_ASAP7_75t_R c9003(
.A1(net8855),
.A2(net9038),
.B(net6214),
.Y(net9049)
);

CKINVDCx16_ASAP7_75t_R c9004(
.A(net10358),
.Y(net9050)
);

CKINVDCx20_ASAP7_75t_R c9005(
.A(net10358),
.Y(net9051)
);

NOR2xp33_ASAP7_75t_R c9006(
.A(net9034),
.B(net9852),
.Y(net9052)
);

AOI21xp5_ASAP7_75t_R c9007(
.A1(net9044),
.A2(net9018),
.B(net7982),
.Y(net9053)
);

FAx1_ASAP7_75t_R c9008(
.A(net9037),
.B(net9026),
.CI(net10140),
.SN(net9054)
);

MAJIxp5_ASAP7_75t_R c9009(
.A(net7971),
.B(net9051),
.C(net9053),
.Y(net9055)
);

MAJx2_ASAP7_75t_R c9010(
.A(net9027),
.B(net9055),
.C(net9052),
.Y(net9056)
);

MAJx3_ASAP7_75t_R c9011(
.A(net8927),
.B(net9050),
.C(net10086),
.Y(net9057)
);

NAND3x1_ASAP7_75t_R c9012(
.A(net9046),
.B(net9057),
.C(net9999),
.Y(net9058)
);

NAND3x2_ASAP7_75t_R c9013(
.B(net6329),
.C(net8199),
.A(net8939),
.Y(net9059)
);

NAND3xp33_ASAP7_75t_R c9014(
.A(net8056),
.B(net8840),
.C(net9037),
.Y(net9060)
);

NOR3x1_ASAP7_75t_R c9015(
.A(net9037),
.B(net9688),
.C(net10074),
.Y(net9061)
);

AOI33xp33_ASAP7_75t_R c9016(
.A1(net9036),
.A2(net9052),
.A3(net9050),
.B1(net9060),
.B2(net9037),
.B3(net8939),
.Y(net9062)
);

NOR3x2_ASAP7_75t_R c9017(
.B(net9015),
.C(net9019),
.A(net8046),
.Y(net9063)
);

NOR3xp33_ASAP7_75t_R c9018(
.A(net9024),
.B(net9058),
.C(net9048),
.Y(net9064)
);

OA21x2_ASAP7_75t_R c9019(
.A1(net8865),
.A2(net9057),
.B(net9044),
.Y(net9065)
);

OAI21x1_ASAP7_75t_R c9020(
.A1(net9060),
.A2(net9030),
.B(net9052),
.Y(net9066)
);

OA222x2_ASAP7_75t_R c9021(
.A1(net5332),
.A2(net9065),
.B1(net9052),
.B2(net9060),
.C1(net7826),
.C2(net9037),
.Y(net9067)
);

OAI21xp33_ASAP7_75t_R c9022(
.A1(net8136),
.A2(net8851),
.B(net9048),
.Y(net9068)
);

OAI21xp5_ASAP7_75t_R c9023(
.A1(net7267),
.A2(net8888),
.B(net9060),
.Y(net9069)
);

NOR4xp75_ASAP7_75t_R c9024(
.A(net9062),
.B(net8960),
.C(net9058),
.D(net9060),
.Y(net9070)
);

OR3x1_ASAP7_75t_R c9025(
.A(net8872),
.B(net9054),
.C(net9060),
.Y(net9071)
);

OR3x2_ASAP7_75t_R c9026(
.A(net7247),
.B(net9063),
.C(net9067),
.Y(net9072)
);

OR3x4_ASAP7_75t_R c9027(
.A(net9026),
.B(net9064),
.C(net9048),
.Y(net9073)
);

AND3x1_ASAP7_75t_R c9028(
.A(net9069),
.B(net9039),
.C(net9045),
.Y(net9074)
);

AND3x2_ASAP7_75t_R c9029(
.A(net9032),
.B(net9073),
.C(net9071),
.Y(net9075)
);

AND3x4_ASAP7_75t_R c9030(
.A(net9056),
.B(net9037),
.C(out4),
.Y(net9076)
);

AO21x1_ASAP7_75t_R c9031(
.A1(net9061),
.A2(net9071),
.B(net10090),
.Y(net9077)
);

OA33x2_ASAP7_75t_R c9032(
.A1(net9066),
.A2(net8993),
.A3(net9071),
.B1(net8939),
.B2(net8148),
.B3(net9060),
.Y(net9078)
);

AO21x2_ASAP7_75t_R c9033(
.A1(net8941),
.A2(net9078),
.B(net10090),
.Y(net9079)
);

AOI21x1_ASAP7_75t_R c9034(
.A1(net9005),
.A2(net9071),
.B(net9068),
.Y(net9080)
);

AOI21xp33_ASAP7_75t_R c9035(
.A1(net9070),
.A2(net8940),
.B(net9079),
.Y(net9081)
);

AOI21xp5_ASAP7_75t_R c9036(
.A1(net8944),
.A2(net9743),
.B(net10086),
.Y(net9082)
);

FAx1_ASAP7_75t_R c9037(
.A(net9072),
.B(net9060),
.CI(net9976),
.SN(net9083)
);

MAJIxp5_ASAP7_75t_R c9038(
.A(net9079),
.B(net9083),
.C(net9082),
.Y(net9084)
);

O2A1O1Ixp33_ASAP7_75t_R c9039(
.A1(net7868),
.A2(net9077),
.B(net9688),
.C(out7)
);

O2A1O1Ixp5_ASAP7_75t_R merge9040(
.A1(net4887),
.A2(net5870),
.B(net5872),
.C(net5706),
.Y(net9085)
);

CKINVDCx5p33_ASAP7_75t_R merge9041(
.A(net10414),
.Y(net9086)
);

SDFLx4_ASAP7_75t_R merge9042(
.D(net1726),
.SE(net1606),
.SI(net1700),
.CLK(clk),
.QN(net9087)
);

DFFASRHQNx1_ASAP7_75t_R merge9043(
.D(net4654),
.RESETN(net3701),
.SETN(net3728),
.CLK(clk),
.QN(net9088)
);

ICGx5p33DC_ASAP7_75t_R merge9044(
.ENA(net848),
.SE(net825),
.CLK(clk),
.GCLK(net9089)
);

ICGx6p67DC_ASAP7_75t_R merge9045(
.ENA(net400),
.SE(net142),
.CLK(clk),
.GCLK(net9090)
);

ICGx8DC_ASAP7_75t_R merge9046(
.ENA(net6572),
.SE(net7441),
.CLK(clk),
.GCLK(net9091)
);

NOR2xp67_ASAP7_75t_R merge9047(
.A(net1467),
.B(net1474),
.Y(net9092)
);

OA211x2_ASAP7_75t_R merge9048(
.A1(net2731),
.A2(net3239),
.B(net3638),
.C(net3629),
.Y(net9093)
);

OA22x2_ASAP7_75t_R merge9049(
.A1(net7056),
.A2(net5105),
.B1(net7202),
.B2(net10288),
.Y(net9094)
);

SDFHx1_ASAP7_75t_R merge9050(
.D(net2774),
.SE(net2780),
.SI(net1875),
.CLK(clk),
.QN(net9095)
);

ICGx1_ASAP7_75t_R merge9051(
.ENA(net3076),
.SE(net3005),
.CLK(clk),
.GCLK(net9096)
);

CKINVDCx6p67_ASAP7_75t_R merge9052(
.A(net10391),
.Y(net9097)
);

OA31x2_ASAP7_75t_R merge9053(
.A1(net6273),
.A2(net7922),
.A3(net8076),
.B1(net8093),
.Y(net9098)
);

ICGx2_ASAP7_75t_R merge9054(
.ENA(net89),
.SE(net503),
.CLK(clk),
.GCLK(net9099)
);

OAI211xp5_ASAP7_75t_R merge9055(
.A1(net5105),
.A2(net6204),
.B(net5384),
.C(net5402),
.Y(net9100)
);

OAI22x1_ASAP7_75t_R merge9056(
.A1(net5240),
.A2(net5277),
.B1(net5320),
.B2(net5346),
.Y(net9101)
);

CKINVDCx8_ASAP7_75t_R merge9057(
.A(net10363),
.Y(net9102)
);

CKINVDCx9p33_ASAP7_75t_R merge9058(
.A(net10526),
.Y(net9103)
);

HB1xp67_ASAP7_75t_R merge9059(
.A(net10015),
.Y(net9104)
);

ICGx2p67DC_ASAP7_75t_R merge9060(
.ENA(net1046),
.SE(net1020),
.CLK(clk),
.GCLK(net9105)
);

OAI22xp33_ASAP7_75t_R merge9061(
.A1(net7706),
.A2(net7711),
.B1(net7727),
.B2(net7767),
.Y(net9106)
);

ICGx3_ASAP7_75t_R merge9062(
.ENA(net1856),
.SE(net2843),
.CLK(clk),
.GCLK(net9107)
);

OAI22xp5_ASAP7_75t_R merge9063(
.A1(net8776),
.A2(net8694),
.B1(net8897),
.B2(net9847),
.Y(net9108)
);

OAI31xp33_ASAP7_75t_R merge9064(
.A1(net7198),
.A2(net8934),
.A3(net8841),
.B(net8936),
.Y(net9109)
);

OAI31xp67_ASAP7_75t_R merge9065(
.A1(net8148),
.A2(net8975),
.A3(net9025),
.B(net8718),
.Y(net9110)
);

OR2x2_ASAP7_75t_R merge9066(
.A(net7957),
.B(net7393),
.Y(net9111)
);

OR4x1_ASAP7_75t_R merge9067(
.A(net7860),
.B(net7810),
.C(net7886),
.D(net7947),
.Y(net9112)
);

HB2xp67_ASAP7_75t_R merge9068(
.A(net10437),
.Y(net9113)
);

ICGx4DC_ASAP7_75t_R merge9069(
.ENA(net6526),
.SE(net4766),
.CLK(clk),
.GCLK(net9114)
);

OR4x2_ASAP7_75t_R merge9070(
.A(net8410),
.B(net8454),
.C(net8471),
.D(net8393),
.Y(net9115)
);

MAJx2_ASAP7_75t_R merge9071(
.A(net3022),
.B(net2829),
.C(net3001),
.Y(net9116)
);

HB3xp67_ASAP7_75t_R merge9072(
.A(net10493),
.Y(net9117)
);

MAJx3_ASAP7_75t_R merge9073(
.A(net535),
.B(net1476),
.C(net2131),
.Y(net9118)
);

NAND3x1_ASAP7_75t_R merge9074(
.A(net4275),
.B(net4268),
.C(net9775),
.Y(net9119)
);

HB4xp67_ASAP7_75t_R merge9075(
.A(net10426),
.Y(net9120)
);

ICGx4_ASAP7_75t_R merge9076(
.ENA(net203),
.SE(net181),
.CLK(clk),
.GCLK(net9121)
);

INVx11_ASAP7_75t_R merge9077(
.A(net10398),
.Y(net9122)
);

OR2x4_ASAP7_75t_R merge9078(
.A(net3322),
.B(net3429),
.Y(net9123)
);

NAND3x2_ASAP7_75t_R merge9079(
.B(net3173),
.C(net3992),
.A(net9860),
.Y(net9124)
);

ICGx5_ASAP7_75t_R merge9080(
.ENA(net816),
.SE(net736),
.CLK(clk),
.GCLK(net9125)
);

A2O1A1Ixp33_ASAP7_75t_R merge9081(
.A1(net8526),
.A2(net8516),
.B(net7578),
.C(net8633),
.Y(net9126)
);

AO221x2_ASAP7_75t_R merge9082(
.A1(net6412),
.A2(net6429),
.B1(net6887),
.B2(net6191),
.C(net10291),
.Y(net9127)
);

AND4x1_ASAP7_75t_R merge9083(
.A(net3642),
.B(net2707),
.C(net3624),
.D(net1785),
.Y(net9128)
);

AND4x2_ASAP7_75t_R merge9084(
.A(net8481),
.B(net8486),
.C(net8425),
.D(net8336),
.Y(net9129)
);

INVx13_ASAP7_75t_R merge9085(
.A(net10385),
.Y(net9130)
);

INVx1_ASAP7_75t_R merge9086(
.A(net10080),
.Y(net9131)
);

SDFHx2_ASAP7_75t_R merge9087(
.D(net6451),
.SE(net4177),
.SI(net6026),
.CLK(clk),
.QN(net9132)
);

ICGx5p33DC_ASAP7_75t_R merge9088(
.ENA(net983),
.SE(net1067),
.CLK(clk),
.GCLK(net9133)
);

INVx2_ASAP7_75t_R merge9089(
.A(net10389),
.Y(net9134)
);

OR2x6_ASAP7_75t_R merge9090(
.A(net208),
.B(net1088),
.Y(net9135)
);

ICGx6p67DC_ASAP7_75t_R merge9091(
.ENA(net3192),
.SE(net4135),
.CLK(clk),
.GCLK(net9136)
);

INVx3_ASAP7_75t_R merge9092(
.A(net10162),
.Y(net9137)
);

XNOR2x1_ASAP7_75t_R merge9093(
.B(net1247),
.A(net1390),
.Y(net9138)
);

OAI222xp33_ASAP7_75t_R merge9094(
.A1(net8191),
.A2(net8144),
.B1(net8244),
.B2(net7240),
.C1(net8232),
.C2(net6381),
.Y(net9139)
);

AO211x2_ASAP7_75t_R merge9095(
.A1(net8127),
.A2(net5260),
.B(net8146),
.C(net10122),
.Y(net9140)
);

AO22x1_ASAP7_75t_R merge9096(
.A1(net4289),
.A2(net4498),
.B1(net4499),
.B2(net10147),
.Y(net9141)
);

ICGx8DC_ASAP7_75t_R merge9097(
.ENA(net3765),
.SE(net3777),
.CLK(clk),
.GCLK(net9142)
);

INVx4_ASAP7_75t_R merge9098(
.A(net9197),
.Y(net9143)
);

ICGx1_ASAP7_75t_R merge9099(
.ENA(net1330),
.SE(net444),
.CLK(clk),
.GCLK(net9144)
);

INVx5_ASAP7_75t_R merge9100(
.A(net10516),
.Y(net9145)
);

XNOR2x2_ASAP7_75t_R merge9101(
.A(net490),
.B(net645),
.Y(net9146)
);

ICGx2_ASAP7_75t_R merge9102(
.ENA(net5589),
.SE(net5600),
.CLK(clk),
.GCLK(net9147)
);

ICGx2p67DC_ASAP7_75t_R merge9103(
.ENA(net7377),
.SE(net7395),
.CLK(clk),
.GCLK(net9148)
);

INVx6_ASAP7_75t_R merge9104(
.A(net9980),
.Y(net9149)
);

INVx8_ASAP7_75t_R merge9105(
.A(net10454),
.Y(net9150)
);

INVxp33_ASAP7_75t_R merge9106(
.A(net10462),
.Y(net9151)
);

SDFHx3_ASAP7_75t_R merge9107(
.D(net7767),
.SE(net5779),
.SI(net7851),
.CLK(clk),
.QN(net9152)
);

INVxp67_ASAP7_75t_R merge9108(
.A(net10429),
.Y(net9153)
);

AO22x2_ASAP7_75t_R merge9109(
.A1(net5293),
.A2(net4515),
.B1(net5442),
.B2(net5440),
.Y(net9154)
);

BUFx10_ASAP7_75t_R merge9110(
.A(net10534),
.Y(net9155)
);

XNOR2xp5_ASAP7_75t_R merge9111(
.A(net208),
.B(net335),
.Y(net9156)
);

SDFHx4_ASAP7_75t_R merge9112(
.D(net6027),
.SE(net6136),
.SI(net10270),
.CLK(clk),
.QN(net9157)
);

SDFLx1_ASAP7_75t_R merge9113(
.D(net3247),
.SE(net3234),
.SI(net10112),
.CLK(clk),
.QN(net9158)
);

AO31x2_ASAP7_75t_R merge9114(
.A1(net6728),
.A2(net7378),
.A3(net7680),
.B(net7690),
.Y(net9159)
);

BUFx12_ASAP7_75t_R merge9115(
.A(net10460),
.Y(net9160)
);

AOI211x1_ASAP7_75t_R merge9116(
.A1(net1686),
.A2(net1797),
.B(net1818),
.C(net2723),
.Y(net9161)
);

ICGx3_ASAP7_75t_R merge9117(
.ENA(net5529),
.SE(net5623),
.CLK(clk),
.GCLK(net9162)
);

AOI211xp5_ASAP7_75t_R merge9118(
.A1(net3652),
.A2(net5448),
.B(net5490),
.C(net5365),
.Y(net9163)
);

ICGx4DC_ASAP7_75t_R merge9119(
.ENA(net2831),
.SE(net1856),
.CLK(clk),
.GCLK(net9164)
);

AOI22x1_ASAP7_75t_R merge9120(
.A1(net3854),
.A2(net4901),
.B1(net4899),
.B2(net4858),
.Y(net9165)
);

AOI22xp33_ASAP7_75t_R merge9121(
.A1(net1583),
.A2(net1457),
.B1(net1588),
.B2(net1592),
.Y(net9166)
);

SDFLx2_ASAP7_75t_R merge9122(
.D(net6297),
.SE(net5359),
.SI(net3587),
.CLK(clk),
.QN(net9167)
);

XOR2x1_ASAP7_75t_R merge9123(
.A(net1867),
.B(net995),
.Y(net9168)
);

BUFx12f_ASAP7_75t_R merge9124(
.A(net10504),
.Y(net9169)
);

BUFx16f_ASAP7_75t_R merge9125(
.A(net10408),
.Y(net9170)
);

BUFx24_ASAP7_75t_R merge9126(
.A(net9199),
.Y(net9171)
);

ICGx4_ASAP7_75t_R merge9127(
.ENA(net469),
.SE(net470),
.CLK(clk),
.GCLK(net9172)
);

ICGx5_ASAP7_75t_R merge9128(
.ENA(net7386),
.SE(net6508),
.CLK(clk),
.GCLK(net9173)
);

BUFx2_ASAP7_75t_R merge9129(
.A(net10526),
.Y(net9174)
);

AOI22xp5_ASAP7_75t_R merge9130(
.A1(net7794),
.A2(net8665),
.B1(net8580),
.B2(net7574),
.Y(net9175)
);

BUFx3_ASAP7_75t_R merge9131(
.A(net10472),
.Y(net9176)
);

BUFx4_ASAP7_75t_R merge9132(
.A(net10459),
.Y(net9177)
);

AOI31xp33_ASAP7_75t_R merge9133(
.A1(net6955),
.A2(net6961),
.A3(net6113),
.B(net6758),
.Y(net9178)
);

AOI31xp67_ASAP7_75t_R merge9134(
.A1(net7921),
.A2(net8732),
.A3(net8779),
.B(net7935),
.Y(net9179)
);

NAND3xp33_ASAP7_75t_R merge9135(
.A(net3914),
.B(net4009),
.C(net3852),
.Y(net9180)
);

BUFx4f_ASAP7_75t_R merge9136(
.A(net9199),
.Y(net9181)
);

NAND4xp25_ASAP7_75t_R merge9137(
.A(net468),
.B(net4141),
.C(net4244),
.D(net3337),
.Y(net9182)
);

NOR3x1_ASAP7_75t_R merge9138(
.A(net5657),
.B(net5788),
.C(net6705),
.Y(net9183)
);

ICGx5p33DC_ASAP7_75t_R merge9139(
.ENA(net5528),
.SE(net5546),
.CLK(clk),
.GCLK(net9184)
);

BUFx5_ASAP7_75t_R merge9140(
.A(net10457),
.Y(net9185)
);

ICGx6p67DC_ASAP7_75t_R merge9141(
.ENA(net5729),
.SE(net5778),
.CLK(clk),
.GCLK(net9186)
);

SDFLx3_ASAP7_75t_R merge9142(
.D(net5574),
.SE(net8338),
.SI(net8341),
.CLK(clk),
.QN(net9187)
);

ICGx8DC_ASAP7_75t_R merge9143(
.ENA(net5900),
.SE(net5087),
.CLK(clk),
.GCLK(net9188)
);

BUFx6f_ASAP7_75t_R merge9144(
.A(net10367),
.Y(net9189)
);

ICGx1_ASAP7_75t_R merge9145(
.ENA(net982),
.SE(net979),
.CLK(clk),
.GCLK(net9190)
);

BUFx8_ASAP7_75t_R merge9146(
.A(net9970),
.Y(net9191)
);

NAND4xp75_ASAP7_75t_R merge9147(
.A(net3618),
.B(net3676),
.C(net5515),
.D(net5467),
.Y(net9192)
);

CKINVDCx10_ASAP7_75t_R merge9148(
.A(net10503),
.Y(net9193)
);

NOR4xp25_ASAP7_75t_R merge9149(
.A(net5058),
.B(net4515),
.C(net1561),
.D(net3551),
.Y(net9194)
);

CKINVDCx11_ASAP7_75t_R merge9150(
.A(net10473),
.Y(net9195)
);

NOR4xp75_ASAP7_75t_R merge9151(
.A(net8058),
.B(net7759),
.C(net6302),
.D(net4431),
.Y(net9196)
);

CKINVDCx12_ASAP7_75t_R merge9152(
.A(net9746),
.Y(net9197)
);

O2A1O1Ixp33_ASAP7_75t_R merge9153(
.A1(net6264),
.A2(net6289),
.B(net2708),
.C(net5478),
.Y(net9198)
);

SDFLx4_ASAP7_75t_R merge9154(
.D(net42),
.SE(net38),
.SI(net107),
.CLK(clk),
.QN(net9199)
);

ICGx2_ASAP7_75t_R merge9155(
.ENA(net223),
.SE(net1058),
.CLK(clk),
.GCLK(net9200)
);

CKINVDCx14_ASAP7_75t_R merge9156(
.A(net10446),
.Y(net9201)
);

CKINVDCx16_ASAP7_75t_R merge9157(
.A(net10519),
.Y(net9202)
);

ICGx2p67DC_ASAP7_75t_R merge9158(
.ENA(net5540),
.SE(net5546),
.CLK(clk),
.GCLK(net9203)
);

CKINVDCx20_ASAP7_75t_R merge9159(
.A(net10157),
.Y(net9204)
);

O2A1O1Ixp5_ASAP7_75t_R merge9160(
.A1(net4281),
.A2(net8566),
.B(net8990),
.C(net8981),
.Y(net9205)
);

OA211x2_ASAP7_75t_R merge9161(
.A1(net7974),
.A2(net4353),
.B(net7283),
.C(net7269),
.Y(net9206)
);

ICGx3_ASAP7_75t_R merge9162(
.ENA(net6492),
.SE(net6620),
.CLK(clk),
.GCLK(net9207)
);

ICGx4DC_ASAP7_75t_R merge9163(
.ENA(net4139),
.SE(net5055),
.CLK(clk),
.GCLK(net9208)
);

XOR2x2_ASAP7_75t_R merge9164(
.A(net1135),
.B(net323),
.Y(net9209)
);

CKINVDCx5p33_ASAP7_75t_R merge9165(
.A(net10395),
.Y(net9210)
);

ICGx4_ASAP7_75t_R merge9166(
.ENA(net6463),
.SE(net6505),
.CLK(clk),
.GCLK(net9211)
);

CKINVDCx6p67_ASAP7_75t_R merge9167(
.A(net10430),
.Y(net9212)
);

CKINVDCx8_ASAP7_75t_R merge9168(
.A(net10498),
.Y(net9213)
);

OA22x2_ASAP7_75t_R merge9169(
.A1(net2637),
.A2(net5097),
.B1(net6282),
.B2(net6286),
.Y(net9214)
);

OA31x2_ASAP7_75t_R merge9170(
.A1(net6313),
.A2(net7102),
.A3(net8122),
.B1(net8141),
.Y(net9215)
);

ICGx5_ASAP7_75t_R merge9171(
.ENA(net7380),
.SE(net4821),
.CLK(clk),
.GCLK(net9216)
);

ICGx5p33DC_ASAP7_75t_R merge9172(
.ENA(net8258),
.SE(net5531),
.CLK(clk),
.GCLK(net9217)
);

ICGx6p67DC_ASAP7_75t_R merge9173(
.ENA(net3817),
.SE(net3946),
.CLK(clk),
.GCLK(net9218)
);

CKINVDCx9p33_ASAP7_75t_R merge9174(
.A(net10441),
.Y(net9219)
);

XOR2xp5_ASAP7_75t_R merge9175(
.A(net181),
.B(net271),
.Y(net9220)
);

HB1xp67_ASAP7_75t_R merge9176(
.A(net10163),
.Y(net9221)
);

OAI211xp5_ASAP7_75t_R merge9177(
.A1(net7844),
.A2(net6928),
.B(net8645),
.C(net8452),
.Y(net9222)
);

HB2xp67_ASAP7_75t_R merge9178(
.A(net10160),
.Y(net9223)
);

HB3xp67_ASAP7_75t_R merge9179(
.A(net10148),
.Y(net9224)
);

HB4xp67_ASAP7_75t_R merge9180(
.A(net10541),
.Y(net9225)
);

ICGx8DC_ASAP7_75t_R merge9181(
.ENA(net6475),
.SE(net6490),
.CLK(clk),
.GCLK(net9226)
);

INVx11_ASAP7_75t_R merge9182(
.A(net10462),
.Y(net9227)
);

ICGx1_ASAP7_75t_R merge9183(
.ENA(net503),
.SE(net611),
.CLK(clk),
.GCLK(net9228)
);

INVx13_ASAP7_75t_R merge9184(
.A(net10476),
.Y(net9229)
);

ICGx2_ASAP7_75t_R merge9185(
.ENA(net3266),
.SE(net4268),
.CLK(clk),
.GCLK(net9230)
);

INVx1_ASAP7_75t_R merge9186(
.A(net10532),
.Y(net9231)
);

ICGx2p67DC_ASAP7_75t_R merge9187(
.ENA(net1877),
.SE(net155),
.CLK(clk),
.GCLK(net9232)
);

ICGx3_ASAP7_75t_R merge9188(
.ENA(net5630),
.SE(net5573),
.CLK(clk),
.GCLK(net9233)
);

AND2x2_ASAP7_75t_R merge9189(
.A(net246),
.B(net206),
.Y(net9234)
);

INVx2_ASAP7_75t_R merge9190(
.A(net10402),
.Y(net9235)
);

AND2x4_ASAP7_75t_R merge9191(
.A(net5617),
.B(net6575),
.Y(net9236)
);

OAI22x1_ASAP7_75t_R merge9192(
.A1(net7153),
.A2(net6975),
.B1(net5076),
.B2(net10142),
.Y(net9237)
);

INVx3_ASAP7_75t_R merge9193(
.A(net10515),
.Y(net9238)
);

INVx4_ASAP7_75t_R merge9194(
.A(net9746),
.Y(net9239)
);

NOR3x2_ASAP7_75t_R merge9195(
.B(net4325),
.C(net6138),
.A(net10258),
.Y(net9240)
);

DFFASRHQNx1_ASAP7_75t_R merge9196(
.D(net5973),
.RESETN(net6789),
.SETN(net6872),
.CLK(clk),
.QN(net9241)
);

ICGx4DC_ASAP7_75t_R merge9197(
.ENA(net4778),
.SE(net4812),
.CLK(clk),
.GCLK(net9242)
);

OAI22xp33_ASAP7_75t_R merge9198(
.A1(net8766),
.A2(net7466),
.B1(net7890),
.B2(net7876),
.Y(net9243)
);

ICGx4_ASAP7_75t_R merge9199(
.ENA(net979),
.SE(net988),
.CLK(clk),
.GCLK(net9244)
);

OAI22xp5_ASAP7_75t_R merge9200(
.A1(net5883),
.A2(net5305),
.B1(net4448),
.B2(net4353),
.Y(net9245)
);

INVx5_ASAP7_75t_R merge9201(
.A(net10549),
.Y(net9246)
);

ICGx5_ASAP7_75t_R merge9202(
.ENA(net5577),
.SE(net5621),
.CLK(clk),
.GCLK(net9247)
);

INVx6_ASAP7_75t_R merge9203(
.A(net10024),
.Y(net9248)
);

OAI31xp33_ASAP7_75t_R merge9204(
.A1(net7233),
.A2(net8185),
.A3(net7124),
.B(net9048),
.Y(net9249)
);

INVx8_ASAP7_75t_R merge9205(
.A(net10473),
.Y(net9250)
);

INVxp33_ASAP7_75t_R merge9206(
.A(net10505),
.Y(net9251)
);

INVxp67_ASAP7_75t_R merge9207(
.A(net10461),
.Y(net9252)
);

BUFx10_ASAP7_75t_R merge9208(
.A(net10434),
.Y(net9253)
);

NOR3xp33_ASAP7_75t_R merge9209(
.A(net6614),
.B(net8442),
.C(net6734),
.Y(net9254)
);

OAI31xp67_ASAP7_75t_R merge9210(
.A1(net3427),
.A2(net1725),
.A3(net4449),
.B(net3591),
.Y(net9255)
);

OR4x1_ASAP7_75t_R merge9211(
.A(net6806),
.B(net4911),
.C(net7741),
.D(net7721),
.Y(net9256)
);

BUFx12_ASAP7_75t_R merge9212(
.A(net9969),
.Y(net9257)
);

ICGx5p33DC_ASAP7_75t_R merge9213(
.ENA(net2825),
.SE(net3696),
.CLK(clk),
.GCLK(net9258)
);

OR4x2_ASAP7_75t_R merge9214(
.A(net7659),
.B(net7649),
.C(net7705),
.D(net7766),
.Y(net9259)
);

A2O1A1Ixp33_ASAP7_75t_R merge9215(
.A1(net5371),
.A2(net5393),
.B(net5343),
.C(net5377),
.Y(net9260)
);

BUFx12f_ASAP7_75t_R merge9216(
.A(net10426),
.Y(net9261)
);

AND4x1_ASAP7_75t_R merge9217(
.A(net1320),
.B(net3817),
.C(net3994),
.D(net2963),
.Y(net9262)
);

AND4x2_ASAP7_75t_R merge9218(
.A(net4209),
.B(net4203),
.C(net3330),
.D(net2498),
.Y(net9263)
);

BUFx16f_ASAP7_75t_R merge9219(
.A(net10466),
.Y(net9264)
);

BUFx24_ASAP7_75t_R merge9220(
.A(net10054),
.Y(net9265)
);

AO211x2_ASAP7_75t_R merge9221(
.A1(net7986),
.A2(net6198),
.B(net4456),
.C(net6122),
.Y(net9266)
);

BUFx2_ASAP7_75t_R merge9222(
.A(net10039),
.Y(net9267)
);

OA21x2_ASAP7_75t_R merge9223(
.A1(net2469),
.A2(net3506),
.B(net4353),
.Y(net9268)
);

BUFx3_ASAP7_75t_R merge9224(
.A(net10444),
.Y(net9269)
);

BUFx4_ASAP7_75t_R merge9225(
.A(net10392),
.Y(net9270)
);

ICGx6p67DC_ASAP7_75t_R merge9226(
.ENA(net390),
.SE(net611),
.CLK(clk),
.GCLK(net9271)
);

AO22x1_ASAP7_75t_R merge9227(
.A1(net4942),
.A2(net2180),
.B1(net4946),
.B2(net4099),
.Y(net9272)
);

BUFx4f_ASAP7_75t_R merge9228(
.A(net10440),
.Y(net9273)
);

AO22x2_ASAP7_75t_R merge9229(
.A1(net4441),
.A2(net4490),
.B1(net2491),
.B2(net2720),
.Y(net9274)
);

SDFHx1_ASAP7_75t_R merge9230(
.D(net5728),
.SE(net4797),
.SI(net5704),
.CLK(clk),
.QN(net9275)
);

AO31x2_ASAP7_75t_R merge9231(
.A1(net7815),
.A2(net7780),
.A3(net6906),
.B(net7767),
.Y(net9276)
);

AOI211x1_ASAP7_75t_R merge9232(
.A1(net6986),
.A2(net6972),
.B(net6096),
.C(net6099),
.Y(net9277)
);

AOI211xp5_ASAP7_75t_R merge9233(
.A1(net3466),
.A2(net3349),
.B(net1644),
.C(net2373),
.Y(net9278)
);

ICGx8DC_ASAP7_75t_R merge9234(
.ENA(net2828),
.SE(net1890),
.CLK(clk),
.GCLK(net9279)
);

SDFHx2_ASAP7_75t_R merge9235(
.D(net8013),
.SE(net7786),
.SI(net7934),
.CLK(clk),
.QN(net9280)
);

ICGx1_ASAP7_75t_R merge9236(
.ENA(net1389),
.SE(net1417),
.CLK(clk),
.GCLK(net9281)
);

ICGx2_ASAP7_75t_R merge9237(
.ENA(net6464),
.SE(net5589),
.CLK(clk),
.GCLK(net9282)
);

AND2x6_ASAP7_75t_R merge9238(
.A(net436),
.B(net1407),
.Y(net9283)
);

AOI22x1_ASAP7_75t_R merge9239(
.A1(net7068),
.A2(net5110),
.B1(net6913),
.B2(net6180),
.Y(net9284)
);

SDFHx3_ASAP7_75t_R merge9240(
.D(net1373),
.SE(net2487),
.SI(net2486),
.CLK(clk),
.QN(net9285)
);

ICGx2p67DC_ASAP7_75t_R merge9241(
.ENA(net2813),
.SE(net3696),
.CLK(clk),
.GCLK(net9286)
);

AOI22xp33_ASAP7_75t_R merge9242(
.A1(net7534),
.A2(net6624),
.B1(net6845),
.B2(net6842),
.Y(net9287)
);

ICGx3_ASAP7_75t_R merge9243(
.ENA(net7401),
.SE(net6464),
.CLK(clk),
.GCLK(net9288)
);

AOI22xp5_ASAP7_75t_R merge9244(
.A1(net2158),
.A2(net4866),
.B1(net3964),
.B2(net3914),
.Y(net9289)
);

AOI31xp33_ASAP7_75t_R merge9245(
.A1(net6967),
.A2(net6964),
.A3(net8761),
.B(net8537),
.Y(net9290)
);

BUFx5_ASAP7_75t_R merge9246(
.A(net10436),
.Y(net9291)
);

AOI31xp67_ASAP7_75t_R merge9247(
.A1(net6311),
.A2(net7241),
.A3(net5431),
.B(net5369),
.Y(net9292)
);

OAI21x1_ASAP7_75t_R merge9248(
.A1(net913),
.A2(net212),
.B(net1233),
.Y(net9293)
);

NAND4xp25_ASAP7_75t_R merge9249(
.A(net7780),
.B(net6905),
.C(net5928),
.D(net6910),
.Y(net9294)
);

NAND4xp75_ASAP7_75t_R merge9250(
.A(net1598),
.B(net1605),
.C(net3273),
.D(net3348),
.Y(net9295)
);

NOR4xp25_ASAP7_75t_R merge9251(
.A(net5309),
.B(net6151),
.C(net5338),
.D(net5306),
.Y(net9296)
);

HAxp5_ASAP7_75t_R merge9252(
.A(net6489),
.B(net5556),
.CON(net9297)
);

NOR4xp75_ASAP7_75t_R merge9253(
.A(net2339),
.B(net2242),
.C(net2131),
.D(net3006),
.Y(net9298)
);

O2A1O1Ixp33_ASAP7_75t_R merge9254(
.A1(net7033),
.A2(net6273),
.B(net8824),
.C(net8722),
.Y(net9299)
);

O2A1O1Ixp5_ASAP7_75t_R merge9255(
.A1(net5324),
.A2(net3316),
.B(net6180),
.C(net6132),
.Y(net9300)
);

OA211x2_ASAP7_75t_R merge9256(
.A1(net1604),
.A2(net1617),
.B(net710),
.C(net87),
.Y(net9301)
);

OA22x2_ASAP7_75t_R merge9257(
.A1(net7872),
.A2(net5908),
.B1(net7874),
.B2(net10285),
.Y(net9302)
);

OA31x2_ASAP7_75t_R merge9258(
.A1(net2519),
.A2(net1615),
.A3(net1634),
.B1(net10002),
.Y(net9303)
);

OAI211xp5_ASAP7_75t_R merge9259(
.A1(net4908),
.A2(net5804),
.B(net3015),
.C(net6666),
.Y(net9304)
);

OAI22x1_ASAP7_75t_R merge9260(
.A1(net6935),
.A2(net7469),
.B1(net5834),
.B2(net5135),
.Y(net9305)
);

OAI22xp33_ASAP7_75t_R merge9261(
.A1(net7994),
.A2(net8011),
.B1(net4376),
.B2(net4385),
.Y(net9306)
);

OAI22xp5_ASAP7_75t_R merge9262(
.A1(net7139),
.A2(net7226),
.B1(net7047),
.B2(net6080),
.Y(net9307)
);

OAI31xp33_ASAP7_75t_R merge9263(
.A1(net7765),
.A2(net1229),
.A3(net3955),
.B(net10166),
.Y(net9308)
);

OAI31xp67_ASAP7_75t_R merge9264(
.A1(net6508),
.A2(net6895),
.A3(net7926),
.B(net10284),
.Y(net9309)
);

ICGx4DC_ASAP7_75t_R merge9265(
.ENA(net5536),
.SE(net2828),
.CLK(clk),
.GCLK(net9310)
);

OR4x1_ASAP7_75t_R merge9266(
.A(net3449),
.B(net3429),
.C(net3478),
.D(net3175),
.Y(net9311)
);

OR4x2_ASAP7_75t_R merge9267(
.A(net6165),
.B(net4302),
.C(net7867),
.D(net7564),
.Y(net9312)
);

A2O1A1Ixp33_ASAP7_75t_R merge9268(
.A1(net5843),
.A2(net6025),
.B(net5959),
.C(net6026),
.Y(net9313)
);

AND4x1_ASAP7_75t_R merge9269(
.A(net2408),
.B(net2422),
.C(net643),
.D(net1551),
.Y(net9314)
);

SDFHx4_ASAP7_75t_R merge9270(
.D(net1946),
.SE(net1078),
.SI(net3005),
.CLK(clk),
.QN(net9315)
);

ICGx4_ASAP7_75t_R merge9271(
.ENA(net1828),
.SE(net1858),
.CLK(clk),
.GCLK(net9316)
);

AND4x2_ASAP7_75t_R merge9272(
.A(net6229),
.B(net6227),
.C(net7666),
.D(net7837),
.Y(net9317)
);

AO211x2_ASAP7_75t_R merge9273(
.A1(net4124),
.A2(net2459),
.B(net3214),
.C(net4385),
.Y(net9318)
);

AO22x1_ASAP7_75t_R merge9274(
.A1(net1645),
.A2(net1670),
.B1(net2530),
.B2(net1709),
.Y(net9319)
);

AO22x2_ASAP7_75t_R merge9275(
.A1(net6168),
.A2(net6196),
.B1(net3438),
.B2(net3432),
.Y(net9320)
);

AO31x2_ASAP7_75t_R merge9276(
.A1(net3491),
.A2(net3428),
.A3(net3492),
.B(net4360),
.Y(net9321)
);

AOI211x1_ASAP7_75t_R merge9277(
.A1(net3919),
.A2(net3908),
.B(net4852),
.C(net9663),
.Y(net9322)
);

AOI211xp5_ASAP7_75t_R merge9278(
.A1(net8038),
.A2(net4477),
.B(net5359),
.C(net9983),
.Y(net9323)
);

AOI22x1_ASAP7_75t_R merge9279(
.A1(net300),
.A2(net299),
.B1(net2930),
.B2(net2918),
.Y(net9324)
);

SDFLx1_ASAP7_75t_R merge9280(
.D(net7424),
.SE(net7549),
.SI(net5636),
.CLK(clk),
.QN(net9325)
);

AOI22xp33_ASAP7_75t_R merge9281(
.A1(net535),
.A2(net499),
.B1(net442),
.B2(net9948),
.Y(net9326)
);

AOI22xp5_ASAP7_75t_R merge9282(
.A1(net65),
.A2(net142),
.B1(net2933),
.B2(net994),
.Y(net9327)
);

AOI31xp33_ASAP7_75t_R merge9283(
.A1(net2547),
.A2(net3475),
.A3(net4378),
.B(net4264),
.Y(net9328)
);

AOI31xp67_ASAP7_75t_R merge9284(
.A1(net3852),
.A2(net3838),
.A3(net3994),
.B(net9868),
.Y(net9329)
);

NAND4xp25_ASAP7_75t_R merge9285(
.A(net724),
.B(net1662),
.C(net4393),
.D(net3504),
.Y(net9330)
);

NAND4xp75_ASAP7_75t_R merge9286(
.A(net3189),
.B(net3237),
.C(net2201),
.D(net10210),
.Y(net9331)
);

NOR4xp25_ASAP7_75t_R merge9287(
.A(net2019),
.B(net1388),
.C(net394),
.D(net331),
.Y(net9332)
);

NOR4xp75_ASAP7_75t_R merge9288(
.A(net2984),
.B(net4203),
.C(net1364),
.D(net1338),
.Y(net9333)
);

O2A1O1Ixp33_ASAP7_75t_R merge9289(
.A1(net126),
.A2(net221),
.B(net3774),
.C(net3825),
.Y(net9334)
);

O2A1O1Ixp5_ASAP7_75t_R merge9290(
.A1(net6803),
.A2(net6451),
.B(net6723),
.C(net4021),
.Y(net9335)
);

OA211x2_ASAP7_75t_R merge9291(
.A1(net1695),
.A2(net710),
.B(net792),
.C(net797),
.Y(net9336)
);

OA22x2_ASAP7_75t_R merge9292(
.A1(net1153),
.A2(net2110),
.B1(net1194),
.B2(net995),
.Y(net9337)
);

OA31x2_ASAP7_75t_R merge9293(
.A1(net3134),
.A2(net2455),
.A3(net499),
.B1(net496),
.Y(net9338)
);

OAI211xp5_ASAP7_75t_R merge9294(
.A1(net5357),
.A2(net3618),
.B(net7100),
.C(net5266),
.Y(net9339)
);

OAI22x1_ASAP7_75t_R merge9295(
.A1(net3212),
.A2(net2205),
.B1(net4168),
.B2(net3817),
.Y(net9340)
);

OAI22xp33_ASAP7_75t_R merge9296(
.A1(net6183),
.A2(net5996),
.B1(net8018),
.B2(net6132),
.Y(net9341)
);

OAI22xp5_ASAP7_75t_R merge9297(
.A1(net6295),
.A2(net5354),
.B1(net5996),
.B2(net10098),
.Y(net9342)
);

OAI31xp33_ASAP7_75t_R merge9298(
.A1(net8434),
.A2(net8422),
.A3(net8424),
.B(net9908),
.Y(net9343)
);

OAI31xp67_ASAP7_75t_R merge9299(
.A1(net6646),
.A2(net6620),
.A3(net6625),
.B(net6627),
.Y(net9344)
);

OR4x1_ASAP7_75t_R merge9300(
.A(net7095),
.B(net6940),
.C(net3987),
.D(net10284),
.Y(net9345)
);

OR4x2_ASAP7_75t_R merge9301(
.A(net3996),
.B(net4868),
.C(net4893),
.D(net9946),
.Y(net9346)
);

A2O1A1Ixp33_ASAP7_75t_R merge9302(
.A1(net4793),
.A2(net4852),
.B(net6567),
.C(net6614),
.Y(net9347)
);

AND4x1_ASAP7_75t_R merge9303(
.A(net6844),
.B(net6833),
.C(net6624),
.D(net7751),
.Y(net9348)
);

AND4x2_ASAP7_75t_R merge9304(
.A(net5702),
.B(net5704),
.C(net3701),
.D(net6702),
.Y(net9349)
);

AO211x2_ASAP7_75t_R merge9305(
.A1(net5314),
.A2(net5359),
.B(net8002),
.C(net6273),
.Y(net9350)
);

AO22x1_ASAP7_75t_R merge9306(
.A1(net3461),
.A2(net4385),
.B1(net1499),
.B2(net462),
.Y(net9351)
);

AO22x2_ASAP7_75t_R merge9307(
.A1(net5752),
.A2(net5758),
.B1(net6657),
.B2(net6620),
.Y(net9352)
);

AO31x2_ASAP7_75t_R merge9308(
.A1(net1458),
.A2(net1355),
.A3(net2407),
.B(net2403),
.Y(net9353)
);

AOI211x1_ASAP7_75t_R merge9309(
.A1(net5634),
.A2(net5657),
.B(net5548),
.C(net2877),
.Y(net9354)
);

AOI211xp5_ASAP7_75t_R merge9310(
.A1(net8355),
.A2(net8365),
.B(net6572),
.C(net6601),
.Y(net9355)
);

AOI22x1_ASAP7_75t_R merge9311(
.A1(net5612),
.A2(net3780),
.B1(net4754),
.B2(net4678),
.Y(net9356)
);

AOI22xp33_ASAP7_75t_R merge9312(
.A1(net107),
.A2(net932),
.B1(net1012),
.B2(net1043),
.Y(net9357)
);

AOI22xp5_ASAP7_75t_R merge9313(
.A1(net1781),
.A2(net1797),
.B1(net736),
.B2(net741),
.Y(net9358)
);

AOI31xp33_ASAP7_75t_R merge9314(
.A1(net4973),
.A2(net3772),
.A3(net1339),
.B(net1373),
.Y(net9359)
);

AOI31xp67_ASAP7_75t_R merge9315(
.A1(net5968),
.A2(net6891),
.A3(net7674),
.B(net10134),
.Y(net9360)
);

NAND4xp25_ASAP7_75t_R merge9316(
.A(net2540),
.B(net2553),
.C(net3436),
.D(net3315),
.Y(net9361)
);

NAND4xp75_ASAP7_75t_R merge9317(
.A(net6151),
.B(net5866),
.C(net5299),
.D(net4264),
.Y(net9362)
);

NOR4xp25_ASAP7_75t_R merge9318(
.A(net3984),
.B(net6685),
.C(net7655),
.D(net7378),
.Y(net9363)
);

NOR4xp75_ASAP7_75t_R merge9319(
.A(net440),
.B(net444),
.C(net2186),
.D(net2131),
.Y(net9364)
);

O2A1O1Ixp33_ASAP7_75t_R merge9320(
.A1(net5054),
.A2(net5084),
.B(net5081),
.C(net5843),
.Y(net9365)
);

O2A1O1Ixp5_ASAP7_75t_R merge9321(
.A1(net4985),
.A2(net6049),
.B(net6710),
.C(net5883),
.Y(net9366)
);

OA211x2_ASAP7_75t_R merge9322(
.A1(net8009),
.A2(net7883),
.B(net7112),
.C(net7115),
.Y(net9367)
);

OA22x2_ASAP7_75t_R merge9323(
.A1(net6605),
.A2(net4766),
.B1(net5633),
.B2(net5571),
.Y(net9368)
);

OA31x2_ASAP7_75t_R merge9324(
.A1(net6027),
.A2(net1477),
.A3(net534),
.B1(net9835),
.Y(net9369)
);

OAI211xp5_ASAP7_75t_R merge9325(
.A1(net6186),
.A2(net7912),
.B(net8803),
.C(net8852),
.Y(net9370)
);

OAI22x1_ASAP7_75t_R merge9326(
.A1(net2455),
.A2(net3267),
.B1(net1388),
.B2(net3411),
.Y(net9371)
);

OAI22xp33_ASAP7_75t_R merge9327(
.A1(net3555),
.A2(net3519),
.B1(net2626),
.B2(net2638),
.Y(net9372)
);

OAI22xp5_ASAP7_75t_R merge9328(
.A1(net6954),
.A2(net6211),
.B1(net6191),
.B2(net9932),
.Y(net9373)
);

OAI31xp33_ASAP7_75t_R merge9329(
.A1(net3856),
.A2(net2027),
.A3(net4798),
.B(net4828),
.Y(net9374)
);

OAI31xp67_ASAP7_75t_R merge9330(
.A1(net262),
.A2(net26),
.A3(net1895),
.B(net2027),
.Y(net9375)
);

OR4x1_ASAP7_75t_R merge9331(
.A(net5909),
.B(net5908),
.C(net1328),
.D(net3086),
.Y(net9376)
);

OR4x2_ASAP7_75t_R merge9332(
.A(net6966),
.B(net5176),
.C(net2270),
.D(net3057),
.Y(net9377)
);

A2O1A1Ixp33_ASAP7_75t_R merge9333(
.A1(net6136),
.A2(net7959),
.B(net6866),
.C(net7687),
.Y(net9378)
);

AND4x1_ASAP7_75t_R merge9334(
.A(net4809),
.B(net4824),
.C(net5567),
.D(net4849),
.Y(net9379)
);

AND4x2_ASAP7_75t_R merge9335(
.A(net4479),
.B(net4360),
.C(net5188),
.D(net5189),
.Y(net9380)
);

AO211x2_ASAP7_75t_R merge9336(
.A1(net5297),
.A2(net5312),
.B(net3647),
.C(net5466),
.Y(net9381)
);

AO22x1_ASAP7_75t_R merge9337(
.A1(net6126),
.A2(net6332),
.B1(net5267),
.B2(net10258),
.Y(net9382)
);

AO22x2_ASAP7_75t_R merge9338(
.A1(net3325),
.A2(net3283),
.B1(net564),
.B2(net529),
.Y(net9383)
);

AO31x2_ASAP7_75t_R merge9339(
.A1(net2898),
.A2(net2896),
.A3(net2974),
.B(net2967),
.Y(net9384)
);

AOI211x1_ASAP7_75t_R merge9340(
.A1(net921),
.A2(net1971),
.B(net142),
.C(net2829),
.Y(net9385)
);

AOI211xp5_ASAP7_75t_R merge9341(
.A1(net6982),
.A2(net6808),
.B(net6190),
.C(net6191),
.Y(net9386)
);

AOI22x1_ASAP7_75t_R merge9342(
.A1(net8695),
.A2(net7786),
.B1(net8751),
.B2(net8854),
.Y(net9387)
);

AOI22xp33_ASAP7_75t_R merge9343(
.A1(net1024),
.A2(net1058),
.B1(net1921),
.B2(net1971),
.Y(net9388)
);

AOI22xp5_ASAP7_75t_R merge9344(
.A1(net1138),
.A2(net4016),
.B1(net4055),
.B2(net3951),
.Y(net9389)
);

AOI31xp33_ASAP7_75t_R merge9345(
.A1(net958),
.A2(net1251),
.A3(net1060),
.B(net1239),
.Y(net9390)
);

AOI31xp67_ASAP7_75t_R merge9346(
.A1(net994),
.A2(net306),
.A3(net263),
.B(net1080),
.Y(net9391)
);

NAND4xp25_ASAP7_75t_R merge9347(
.A(net5610),
.B(net5931),
.C(net7742),
.D(net6719),
.Y(net9392)
);

NAND4xp75_ASAP7_75t_R merge9348(
.A(net4432),
.B(net5260),
.C(net4289),
.D(net4467),
.Y(net9393)
);

NOR4xp25_ASAP7_75t_R merge9349(
.A(net390),
.B(net1355),
.C(net5867),
.D(net5869),
.Y(net9394)
);

NOR4xp75_ASAP7_75t_R merge9350(
.A(net4112),
.B(net4360),
.C(net2595),
.D(net2561),
.Y(net9395)
);

O2A1O1Ixp33_ASAP7_75t_R merge9351(
.A1(net1199),
.A2(net1193),
.B(net1032),
.C(net2072),
.Y(net9396)
);

O2A1O1Ixp5_ASAP7_75t_R merge9352(
.A1(net3070),
.A2(net3076),
.B(net1211),
.C(net3943),
.Y(net9397)
);

OA211x2_ASAP7_75t_R merge9353(
.A1(net6505),
.A2(net4827),
.B(net6624),
.C(net10020),
.Y(net9398)
);

OA22x2_ASAP7_75t_R merge9354(
.A1(net6200),
.A2(net6046),
.B1(net2495),
.B2(net3326),
.Y(net9399)
);

OA31x2_ASAP7_75t_R merge9355(
.A1(net7566),
.A2(net8366),
.A3(net8454),
.B1(net8424),
.Y(net9400)
);

OAI211xp5_ASAP7_75t_R merge9356(
.A1(net7395),
.A2(net3825),
.B(net6696),
.C(net6694),
.Y(net9401)
);

OAI22x1_ASAP7_75t_R merge9357(
.A1(net2383),
.A2(net2365),
.B1(net3286),
.B2(net3134),
.Y(net9402)
);

OAI22xp33_ASAP7_75t_R merge9358(
.A1(net3450),
.A2(net2591),
.B1(net2612),
.B2(net10062),
.Y(net9403)
);

OAI22xp5_ASAP7_75t_R merge9359(
.A1(net1939),
.A2(net1856),
.B1(net1993),
.B2(net1088),
.Y(net9404)
);

OAI31xp33_ASAP7_75t_R merge9360(
.A1(net3395),
.A2(net3383),
.A3(net4207),
.B(net4324),
.Y(net9405)
);

OAI31xp67_ASAP7_75t_R merge9361(
.A1(net6585),
.A2(net6612),
.A3(net5616),
.B(net5630),
.Y(net9406)
);

OR4x1_ASAP7_75t_R merge9362(
.A(net5022),
.B(net5870),
.C(net2298),
.D(net2297),
.Y(net9407)
);

OR4x2_ASAP7_75t_R merge9363(
.A(net1662),
.B(net1658),
.C(net3464),
.D(net3448),
.Y(net9408)
);

A2O1A1Ixp33_ASAP7_75t_R merge9364(
.A1(net4770),
.A2(net3901),
.B(net5708),
.C(net5704),
.Y(net9409)
);

AND4x1_ASAP7_75t_R merge9365(
.A(net1732),
.B(net2600),
.C(net863),
.D(net884),
.Y(net9410)
);

AND4x2_ASAP7_75t_R merge9366(
.A(net4953),
.B(net7740),
.C(net8614),
.D(net9989),
.Y(net9411)
);

AO211x2_ASAP7_75t_R merge9367(
.A1(net462),
.A2(net641),
.B(net3364),
.C(net2335),
.Y(net9412)
);

AO22x1_ASAP7_75t_R merge9368(
.A1(net5887),
.A2(net5928),
.B1(net5026),
.B2(net4901),
.Y(net9413)
);

AO22x2_ASAP7_75t_R merge9369(
.A1(net6157),
.A2(net6153),
.B1(net7112),
.B2(net10114),
.Y(net9414)
);

AO31x2_ASAP7_75t_R merge9370(
.A1(net400),
.A2(net835),
.A3(net3390),
.B(net3266),
.Y(net9415)
);

AOI211x1_ASAP7_75t_R merge9371(
.A1(net4262),
.A2(net5215),
.B(net5245),
.C(net6080),
.Y(net9416)
);

AOI211xp5_ASAP7_75t_R merge9372(
.A1(net3085),
.A2(net1280),
.B(net396),
.C(net440),
.Y(net9417)
);

AOI22x1_ASAP7_75t_R merge9373(
.A1(net5154),
.A2(net4217),
.B1(net2365),
.B2(net2235),
.Y(net9418)
);

AOI22xp33_ASAP7_75t_R merge9374(
.A1(net4693),
.A2(net4832),
.B1(net5616),
.B2(net10264),
.Y(net9419)
);

AOI22xp5_ASAP7_75t_R merge9375(
.A1(net7151),
.A2(net7139),
.B1(net7076),
.B2(net7123),
.Y(net9420)
);

AOI31xp33_ASAP7_75t_R merge9376(
.A1(net2284),
.A2(net2298),
.A3(net4312),
.B(net4257),
.Y(net9421)
);

AOI31xp67_ASAP7_75t_R merge9377(
.A1(net4203),
.A2(net6080),
.A3(net7906),
.B(net7892),
.Y(net9422)
);

NAND4xp25_ASAP7_75t_R merge9378(
.A(net5255),
.B(net6174),
.C(net6748),
.D(net5908),
.Y(net9423)
);

NAND4xp75_ASAP7_75t_R merge9379(
.A(net6647),
.B(net6688),
.C(net6474),
.D(net6589),
.Y(net9424)
);

NOR4xp25_ASAP7_75t_R merge9380(
.A(net5921),
.B(net6029),
.C(net7817),
.D(net5836),
.Y(net9425)
);

NOR4xp75_ASAP7_75t_R merge9381(
.A(net1391),
.B(net1353),
.C(net1531),
.D(net2518),
.Y(net9426)
);

O2A1O1Ixp33_ASAP7_75t_R merge9382(
.A1(net8854),
.A2(net5262),
.B(net5336),
.C(net9639),
.Y(net9427)
);

O2A1O1Ixp5_ASAP7_75t_R merge9383(
.A1(net5897),
.A2(net5866),
.B(net7106),
.C(net7095),
.Y(net9428)
);

OA211x2_ASAP7_75t_R merge9384(
.A1(net2077),
.A2(net1135),
.B(net995),
.C(net9849),
.Y(net9429)
);

OA22x2_ASAP7_75t_R merge9385(
.A1(net2511),
.A2(net2518),
.B1(net2249),
.B2(net2248),
.Y(net9430)
);

OA31x2_ASAP7_75t_R merge9386(
.A1(net7811),
.A2(net7841),
.A3(net6142),
.B1(net5866),
.Y(net9431)
);

OAI211xp5_ASAP7_75t_R merge9387(
.A1(net261),
.A2(net280),
.B(net2926),
.C(net2907),
.Y(net9432)
);

OAI22x1_ASAP7_75t_R merge9388(
.A1(net5250),
.A2(net5266),
.B1(net4257),
.B2(net5105),
.Y(net9433)
);

OAI22xp33_ASAP7_75t_R merge9389(
.A1(net3337),
.A2(net5116),
.B1(net5386),
.B2(net2637),
.Y(net9434)
);

OAI22xp5_ASAP7_75t_R merge9390(
.A1(net2198),
.A2(net2208),
.B1(net206),
.B2(net1058),
.Y(net9435)
);

OAI31xp33_ASAP7_75t_R merge9391(
.A1(net7561),
.A2(net7374),
.A3(net5736),
.B(net6673),
.Y(net9436)
);

OAI31xp67_ASAP7_75t_R merge9392(
.A1(net2861),
.A2(net2975),
.A3(net2998),
.B(net2914),
.Y(net9437)
);

OR4x1_ASAP7_75t_R merge9393(
.A(net2301),
.B(net3162),
.C(net3244),
.D(net3250),
.Y(net9438)
);

OR4x2_ASAP7_75t_R merge9394(
.A(net7580),
.B(net7523),
.C(net8468),
.D(net8318),
.Y(net9439)
);

A2O1A1Ixp33_ASAP7_75t_R merge9395(
.A1(net5798),
.A2(net5788),
.B(net3989),
.C(net4937),
.Y(net9440)
);

AND4x1_ASAP7_75t_R merge9396(
.A(net3162),
.B(net3183),
.C(net3381),
.D(net4325),
.Y(net9441)
);

AND4x2_ASAP7_75t_R merge9397(
.A(net3459),
.B(net2383),
.C(net3469),
.D(net2582),
.Y(net9442)
);

AO211x2_ASAP7_75t_R merge9398(
.A1(net2502),
.A2(net3438),
.B(net4453),
.C(net1526),
.Y(net9443)
);

AO22x1_ASAP7_75t_R merge9399(
.A1(net4792),
.A2(net4852),
.B1(net1402),
.B2(net3245),
.Y(net9444)
);

AO22x2_ASAP7_75t_R merge9400(
.A1(net5939),
.A2(net4981),
.B1(net5032),
.B2(net5001),
.Y(net9445)
);

AO31x2_ASAP7_75t_R merge9401(
.A1(net3884),
.A2(net3856),
.A3(net3855),
.B(net3731),
.Y(net9446)
);

AOI211x1_ASAP7_75t_R merge9402(
.A1(net3908),
.A2(net5656),
.B(net7571),
.C(net7578),
.Y(net9447)
);

AOI211xp5_ASAP7_75t_R merge9403(
.A1(net433),
.A2(net428),
.B(net5003),
.C(net5870),
.Y(net9448)
);

AOI22x1_ASAP7_75t_R merge9404(
.A1(net6742),
.A2(net6866),
.B1(net6680),
.B2(net6678),
.Y(net9449)
);

AOI22xp33_ASAP7_75t_R merge9405(
.A1(net5013),
.A2(net5880),
.B1(net5024),
.B2(net5056),
.Y(net9450)
);

AOI22xp5_ASAP7_75t_R merge9406(
.A1(net7050),
.A2(net6198),
.B1(net8492),
.B2(net8506),
.Y(net9451)
);

AOI31xp33_ASAP7_75t_R merge9407(
.A1(net529),
.A2(net534),
.A3(net536),
.B(net1365),
.Y(net9452)
);

AOI31xp67_ASAP7_75t_R merge9408(
.A1(net1435),
.A2(net606),
.A3(net1532),
.B(net1504),
.Y(net9453)
);

NAND4xp25_ASAP7_75t_R merge9409(
.A(net4322),
.B(net6165),
.C(net6221),
.D(net5260),
.Y(net9454)
);

NAND4xp75_ASAP7_75t_R merge9410(
.A(net4583),
.B(net5198),
.C(net3334),
.D(net3400),
.Y(net9455)
);

NOR4xp25_ASAP7_75t_R merge9411(
.A(net3863),
.B(net3856),
.C(net3896),
.D(net3880),
.Y(net9456)
);

NOR4xp75_ASAP7_75t_R merge9412(
.A(net728),
.B(net730),
.C(net1655),
.D(net1561),
.Y(net9457)
);

O2A1O1Ixp33_ASAP7_75t_R merge9413(
.A1(net3069),
.A2(net4324),
.B(net10207),
.C(net10243),
.Y(net9458)
);

O2A1O1Ixp5_ASAP7_75t_R merge9414(
.A1(net2966),
.A2(net3929),
.B(net4882),
.C(net4857),
.Y(net9459)
);

OA211x2_ASAP7_75t_R merge9415(
.A1(net3949),
.A2(net3033),
.B(net4001),
.C(net4893),
.Y(net9460)
);

OAI21xp33_ASAP7_75t_R merge9416(
.A1(net1172),
.A2(net3014),
.B(net3942),
.Y(net9461)
);

OA22x2_ASAP7_75t_R merge9417(
.A1(net5540),
.A2(net5545),
.B1(net5680),
.B2(net10266),
.Y(net9462)
);

OA31x2_ASAP7_75t_R merge9418(
.A1(net1654),
.A2(net2529),
.A3(net2385),
.B1(net2518),
.Y(net9463)
);

OAI211xp5_ASAP7_75t_R merge9419(
.A1(net1491),
.A2(net4283),
.B(net3266),
.C(net10211),
.Y(net9464)
);

OAI22x1_ASAP7_75t_R merge9420(
.A1(net5868),
.A2(net7674),
.B1(net10224),
.B2(net10296),
.Y(net9465)
);

OAI22xp33_ASAP7_75t_R merge9421(
.A1(net1067),
.A2(net2919),
.B1(net3002),
.B2(net3950),
.Y(net9466)
);

SDFLx2_ASAP7_75t_R merge9422(
.D(net4410),
.SE(net1627),
.SI(net3438),
.CLK(clk),
.QN(net9467)
);

OAI22xp5_ASAP7_75t_R merge9423(
.A1(net2276),
.A2(net2361),
.B1(net487),
.B2(net1227),
.Y(net9468)
);

SDFLx3_ASAP7_75t_R merge9424(
.D(net3057),
.SE(net407),
.SI(net3180),
.CLK(clk),
.QN(net9469)
);

OAI31xp33_ASAP7_75t_R merge9425(
.A1(net3886),
.A2(net2938),
.A3(net3943),
.B(net4055),
.Y(net9470)
);

OAI31xp67_ASAP7_75t_R merge9426(
.A1(net1869),
.A2(net2951),
.A3(net3835),
.B(net2874),
.Y(net9471)
);

OR4x1_ASAP7_75t_R merge9427(
.A(net3739),
.B(net4691),
.C(net3834),
.D(net4700),
.Y(net9472)
);

OR4x2_ASAP7_75t_R merge9428(
.A(net6678),
.B(net6701),
.C(net5994),
.D(net6038),
.Y(net9473)
);

A2O1A1Ixp33_ASAP7_75t_R merge9429(
.A1(net1699),
.A2(net1693),
.B(net3489),
.C(net4375),
.Y(net9474)
);

AND4x1_ASAP7_75t_R merge9430(
.A(net5835),
.B(net5853),
.C(net6743),
.D(net6703),
.Y(net9475)
);

AND4x2_ASAP7_75t_R merge9431(
.A(net6772),
.B(net6791),
.C(net4941),
.D(net4985),
.Y(net9476)
);

AO211x2_ASAP7_75t_R merge9432(
.A1(net5099),
.A2(net2393),
.B(net647),
.C(net689),
.Y(net9477)
);

AO22x1_ASAP7_75t_R merge9433(
.A1(net5076),
.A2(net7802),
.B1(net7886),
.B2(net10147),
.Y(net9478)
);

AO22x2_ASAP7_75t_R merge9434(
.A1(net348),
.A2(net384),
.B1(net1251),
.B2(net1301),
.Y(net9479)
);

AO31x2_ASAP7_75t_R merge9435(
.A1(net4122),
.A2(net4293),
.A3(net4332),
.B(net4325),
.Y(net9480)
);

AOI211x1_ASAP7_75t_R merge9436(
.A1(net3256),
.A2(net534),
.B(net1605),
.C(net1597),
.Y(net9481)
);

AOI211xp5_ASAP7_75t_R merge9437(
.A1(net2072),
.A2(net1947),
.B(net2070),
.C(net1971),
.Y(net9482)
);

AOI22x1_ASAP7_75t_R merge9438(
.A1(net564),
.A2(net879),
.B1(net850),
.B2(net10179),
.Y(net9483)
);

AOI22xp33_ASAP7_75t_R merge9439(
.A1(net4046),
.A2(net4063),
.B1(net467),
.B2(net444),
.Y(net9484)
);

AOI22xp5_ASAP7_75t_R merge9440(
.A1(net3136),
.A2(net3134),
.B1(net4043),
.B2(net3943),
.Y(net9485)
);

AOI31xp33_ASAP7_75t_R merge9441(
.A1(net2951),
.A2(net2758),
.A3(net3890),
.B(net2014),
.Y(net9486)
);

AOI31xp67_ASAP7_75t_R merge9442(
.A1(net2993),
.A2(net2942),
.A3(net4720),
.B(net4692),
.Y(net9487)
);

NAND4xp25_ASAP7_75t_R merge9443(
.A(net2705),
.B(net2726),
.C(net3551),
.D(net9733),
.Y(net9488)
);

NAND4xp75_ASAP7_75t_R merge9444(
.A(net2431),
.B(net1572),
.C(net4315),
.D(net4330),
.Y(net9489)
);

NOR4xp25_ASAP7_75t_R merge9445(
.A(net4515),
.B(net5418),
.C(net5125),
.D(net4994),
.Y(net9490)
);

NOR4xp75_ASAP7_75t_R merge9446(
.A(net2323),
.B(net1540),
.C(net6358),
.D(net9708),
.Y(net9491)
);

O2A1O1Ixp33_ASAP7_75t_R merge9447(
.A1(net4231),
.A2(net4293),
.B(net3419),
.C(net5240),
.Y(net9492)
);

O2A1O1Ixp5_ASAP7_75t_R merge9448(
.A1(net7527),
.A2(net8438),
.B(net5636),
.C(net7435),
.Y(net9493)
);

OA211x2_ASAP7_75t_R merge9449(
.A1(net5847),
.A2(net5827),
.B(net7518),
.C(net7484),
.Y(net9494)
);

OA22x2_ASAP7_75t_R merge9450(
.A1(net6970),
.A2(net6987),
.B1(net2436),
.B2(net622),
.Y(net9495)
);

OA31x2_ASAP7_75t_R merge9451(
.A1(net4031),
.A2(net5028),
.A3(net5082),
.B1(net4981),
.Y(net9496)
);

OAI211xp5_ASAP7_75t_R merge9452(
.A1(net462),
.A2(net1571),
.B(net1537),
.C(net643),
.Y(net9497)
);

OAI22x1_ASAP7_75t_R merge9453(
.A1(net263),
.A2(net261),
.B1(net2280),
.B2(net3025),
.Y(net9498)
);

OAI22xp33_ASAP7_75t_R merge9454(
.A1(net7750),
.A2(net4963),
.B1(net3294),
.B2(net1336),
.Y(net9499)
);

OAI22xp5_ASAP7_75t_R merge9455(
.A1(net7848),
.A2(net7885),
.B1(net7585),
.B2(net8433),
.Y(net9500)
);

OAI31xp33_ASAP7_75t_R merge9456(
.A1(net7045),
.A2(net6027),
.A3(net5945),
.B(net6053),
.Y(net9501)
);

OAI31xp67_ASAP7_75t_R merge9457(
.A1(net1224),
.A2(net1247),
.A3(net3290),
.B(net3316),
.Y(net9502)
);

OR4x1_ASAP7_75t_R merge9458(
.A(net6732),
.B(net6652),
.C(net5823),
.D(net5806),
.Y(net9503)
);

OR4x2_ASAP7_75t_R merge9459(
.A(net4834),
.B(net4539),
.C(net7923),
.D(net5197),
.Y(net9504)
);

A2O1A1Ixp33_ASAP7_75t_R merge9460(
.A1(net7432),
.A2(net7522),
.B(net7605),
.C(net4852),
.Y(net9505)
);

AND4x1_ASAP7_75t_R merge9461(
.A(net1602),
.B(net1605),
.C(net3348),
.D(net3447),
.Y(net9506)
);

AND4x2_ASAP7_75t_R merge9462(
.A(net3604),
.B(net3437),
.C(net3262),
.D(net9986),
.Y(net9507)
);

AO211x2_ASAP7_75t_R merge9463(
.A1(net155),
.A2(net1081),
.B(net3788),
.C(net3743),
.Y(net9508)
);

AO22x1_ASAP7_75t_R merge9464(
.A1(net2037),
.A2(net2049),
.B1(net3714),
.B2(net3731),
.Y(net9509)
);

AO22x2_ASAP7_75t_R merge9465(
.A1(net1032),
.A2(net983),
.B1(net967),
.B2(net988),
.Y(net9510)
);

AO31x2_ASAP7_75t_R merge9466(
.A1(net1264),
.A2(net1270),
.A3(net4188),
.B(net4195),
.Y(net9511)
);

AOI211x1_ASAP7_75t_R merge9467(
.A1(net5886),
.A2(net3859),
.B(net1358),
.C(net1367),
.Y(net9512)
);

AOI211xp5_ASAP7_75t_R merge9468(
.A1(net7245),
.A2(net6329),
.B(net4968),
.C(net5423),
.Y(net9513)
);

AOI22x1_ASAP7_75t_R merge9469(
.A1(net6490),
.A2(net6578),
.B1(net7657),
.B2(net7624),
.Y(net9514)
);

AOI22xp33_ASAP7_75t_R merge9470(
.A1(net4678),
.A2(net4701),
.B1(net4649),
.B2(net4700),
.Y(net9515)
);

AOI22xp5_ASAP7_75t_R merge9471(
.A1(net3412),
.A2(net3404),
.B1(net5999),
.B2(net5245),
.Y(net9516)
);

AOI31xp33_ASAP7_75t_R merge9472(
.A1(net6483),
.A2(net6856),
.A3(net7426),
.B(net6694),
.Y(net9517)
);

AOI31xp67_ASAP7_75t_R merge9473(
.A1(net1663),
.A2(net1673),
.A3(net5247),
.B(net5276),
.Y(net9518)
);

NAND4xp25_ASAP7_75t_R merge9474(
.A(net4157),
.B(net3163),
.C(net2951),
.D(net4800),
.Y(net9519)
);

NAND4xp75_ASAP7_75t_R merge9475(
.A(net1352),
.B(net589),
.C(net3310),
.D(net3290),
.Y(net9520)
);

NOR4xp25_ASAP7_75t_R merge9476(
.A(net2594),
.B(net2474),
.C(net782),
.D(net742),
.Y(net9521)
);

NOR4xp75_ASAP7_75t_R merge9477(
.A(net3105),
.B(net3176),
.C(net4784),
.D(net4797),
.Y(net9522)
);

O2A1O1Ixp33_ASAP7_75t_R merge9478(
.A1(net6052),
.A2(net5980),
.B(net610),
.C(net558),
.Y(net9523)
);

O2A1O1Ixp5_ASAP7_75t_R merge9479(
.A1(net279),
.A2(net283),
.B(net6668),
.C(net6683),
.Y(net9524)
);

OA211x2_ASAP7_75t_R merge9480(
.A1(net138),
.A2(net1852),
.B(net271),
.C(net1259),
.Y(net9525)
);

OA22x2_ASAP7_75t_R merge9481(
.A1(net3027),
.A2(net2990),
.B1(net1708),
.B2(net1736),
.Y(net9526)
);

OA31x2_ASAP7_75t_R merge9482(
.A1(net6488),
.A2(net6702),
.A3(net7607),
.B1(net5772),
.Y(net9527)
);

OAI211xp5_ASAP7_75t_R merge9483(
.A1(net1459),
.A2(net4203),
.B(net2995),
.C(net2036),
.Y(net9528)
);

OAI22x1_ASAP7_75t_R merge9484(
.A1(net3041),
.A2(net3014),
.B1(net5115),
.B2(net7012),
.Y(net9529)
);

OAI22xp33_ASAP7_75t_R merge9485(
.A1(net4880),
.A2(net7732),
.B1(net10091),
.B2(net10143),
.Y(net9530)
);

OAI22xp5_ASAP7_75t_R merge9486(
.A1(net3575),
.A2(net3570),
.B1(net845),
.B2(net831),
.Y(net9531)
);

OAI31xp33_ASAP7_75t_R merge9487(
.A1(net255),
.A2(net294),
.A3(net3343),
.B(net2475),
.Y(net9532)
);

OAI31xp67_ASAP7_75t_R merge9488(
.A1(net2235),
.A2(net2253),
.A3(net3264),
.B(net1337),
.Y(net9533)
);

OR4x1_ASAP7_75t_R merge9489(
.A(net3098),
.B(net4131),
.C(net404),
.D(net1328),
.Y(net9534)
);

OR4x2_ASAP7_75t_R merge9490(
.A(net4171),
.B(net4086),
.C(net7674),
.D(net10283),
.Y(net9535)
);

A2O1A1Ixp33_ASAP7_75t_R merge9491(
.A1(net7558),
.A2(net7374),
.B(net8408),
.C(net7578),
.Y(net9536)
);

AND4x1_ASAP7_75t_R merge9492(
.A(net880),
.B(net850),
.C(net6112),
.D(net5934),
.Y(net9537)
);

AND4x2_ASAP7_75t_R merge9493(
.A(net115),
.B(net2973),
.C(net3200),
.D(net3167),
.Y(net9538)
);

AO211x2_ASAP7_75t_R merge9494(
.A1(net3309),
.A2(net3282),
.B(net281),
.C(net2860),
.Y(net9539)
);

AO22x1_ASAP7_75t_R merge9495(
.A1(net3504),
.A2(net4406),
.B1(net4309),
.B2(net4355),
.Y(net9540)
);

AO22x2_ASAP7_75t_R merge9496(
.A1(net2114),
.A2(net1179),
.B1(net3025),
.B2(net10067),
.Y(net9541)
);

AO31x2_ASAP7_75t_R merge9497(
.A1(net770),
.A2(net765),
.A3(net6816),
.B(net6164),
.Y(net9542)
);

AOI211x1_ASAP7_75t_R merge9498(
.A1(net4324),
.A2(net5172),
.B(net534),
.C(net3421),
.Y(net9543)
);

AOI211xp5_ASAP7_75t_R merge9499(
.A1(net3244),
.A2(net2386),
.B(net4872),
.C(net4880),
.Y(net9544)
);

AOI22x1_ASAP7_75t_R merge9500(
.A1(net5112),
.A2(net5016),
.B1(net1059),
.B2(net2400),
.Y(net9545)
);

AOI22xp33_ASAP7_75t_R merge9501(
.A1(net4836),
.A2(net3234),
.B1(net4167),
.B2(net4170),
.Y(net9546)
);

AOI22xp5_ASAP7_75t_R merge9502(
.A1(net4287),
.A2(net4289),
.B1(net8592),
.B2(net8566),
.Y(net9547)
);

AOI31xp33_ASAP7_75t_R merge9503(
.A1(net2952),
.A2(net223),
.A3(net2268),
.B(net10195),
.Y(net9548)
);

AOI31xp67_ASAP7_75t_R merge9504(
.A1(net5232),
.A2(net5216),
.A3(net7028),
.B(net5197),
.Y(net9549)
);

NAND4xp25_ASAP7_75t_R merge9505(
.A(net3425),
.B(net2502),
.C(net3992),
.D(net4845),
.Y(net9550)
);

NAND4xp75_ASAP7_75t_R merge9506(
.A(net4805),
.B(net3864),
.C(net3996),
.D(net3940),
.Y(net9551)
);

NOR4xp25_ASAP7_75t_R merge9507(
.A(net8539),
.B(net8521),
.C(net8370),
.D(net7670),
.Y(net9552)
);

NOR4xp75_ASAP7_75t_R merge9508(
.A(net2412),
.B(net2359),
.C(net151),
.D(net271),
.Y(net9553)
);

O2A1O1Ixp33_ASAP7_75t_R merge9509(
.A1(net6809),
.A2(net6026),
.B(net6334),
.C(net6297),
.Y(net9554)
);

O2A1O1Ixp5_ASAP7_75t_R merge9510(
.A1(net2733),
.A2(net3604),
.B(net6076),
.C(net5076),
.Y(net9555)
);

OA211x2_ASAP7_75t_R merge9511(
.A1(net2411),
.A2(net2034),
.B(net264),
.C(net261),
.Y(net9556)
);

OA22x2_ASAP7_75t_R merge9512(
.A1(net6144),
.A2(net1481),
.B1(net1622),
.B2(net10270),
.Y(net9557)
);

OA31x2_ASAP7_75t_R merge9513(
.A1(net1273),
.A2(net3085),
.A3(net3063),
.B1(net3066),
.Y(net9558)
);

OAI211xp5_ASAP7_75t_R merge9514(
.A1(net1150),
.A2(net2063),
.B(net2920),
.C(net1010),
.Y(net9559)
);

OAI22x1_ASAP7_75t_R merge9515(
.A1(net5632),
.A2(net5636),
.B1(net2173),
.B2(net2180),
.Y(net9560)
);

OAI22xp33_ASAP7_75t_R merge9516(
.A1(net884),
.A2(net738),
.B1(net4309),
.B2(net9795),
.Y(net9561)
);

OAI22xp5_ASAP7_75t_R merge9517(
.A1(net3912),
.A2(net3893),
.B1(net4967),
.B2(net5033),
.Y(net9562)
);

OAI31xp33_ASAP7_75t_R merge9518(
.A1(net3877),
.A2(net4955),
.A3(net5674),
.B(net5617),
.Y(net9563)
);

OAI31xp67_ASAP7_75t_R merge9519(
.A1(net5821),
.A2(net5883),
.A3(net4044),
.B(net6508),
.Y(net9564)
);

OR4x1_ASAP7_75t_R merge9520(
.A(net4354),
.B(net4333),
.C(net4609),
.D(net5004),
.Y(net9565)
);

OR4x2_ASAP7_75t_R merge9521(
.A(net7642),
.B(net7742),
.C(net4286),
.D(net5257),
.Y(net9566)
);

A2O1A1Ixp33_ASAP7_75t_R merge9522(
.A1(net7716),
.A2(net7710),
.B(net6046),
.C(net4408),
.Y(net9567)
);

AND4x1_ASAP7_75t_R merge9523(
.A(net727),
.B(net2345),
.C(net3345),
.D(net10214),
.Y(net9568)
);

AND4x2_ASAP7_75t_R merge9524(
.A(net5178),
.B(net5118),
.C(net2643),
.D(net891),
.Y(net9569)
);

AO211x2_ASAP7_75t_R merge9525(
.A1(net4267),
.A2(net5043),
.B(net3049),
.C(net6919),
.Y(net9570)
);

AO22x1_ASAP7_75t_R merge9526(
.A1(net6547),
.A2(net6620),
.B1(net1393),
.B2(net1417),
.Y(net9571)
);

AO22x2_ASAP7_75t_R merge9527(
.A1(net6026),
.A2(net7012),
.B1(net5030),
.B2(net2381),
.Y(net9572)
);

AO31x2_ASAP7_75t_R merge9528(
.A1(net1809),
.A2(net2675),
.A3(net5234),
.B(net5229),
.Y(net9573)
);

AOI211x1_ASAP7_75t_R merge9529(
.A1(net1341),
.A2(net444),
.B(net3960),
.C(net4131),
.Y(net9574)
);

AOI211xp5_ASAP7_75t_R merge9530(
.A1(net8551),
.A2(net8548),
.B(net4016),
.C(net1160),
.Y(net9575)
);

AOI22x1_ASAP7_75t_R merge9531(
.A1(net6119),
.A2(net5217),
.B1(net656),
.B2(net490),
.Y(net9576)
);

AOI22xp33_ASAP7_75t_R merge9532(
.A1(net7032),
.A2(net6931),
.B1(net5249),
.B2(net5240),
.Y(net9577)
);

AOI22xp5_ASAP7_75t_R merge9533(
.A1(net2568),
.A2(net2558),
.B1(net3078),
.B2(net2110),
.Y(net9578)
);

AOI31xp33_ASAP7_75t_R merge9534(
.A1(net323),
.A2(net314),
.A3(net3800),
.B(net3812),
.Y(net9579)
);

AOI31xp67_ASAP7_75t_R merge9535(
.A1(net5001),
.A2(net7720),
.A3(net7705),
.B(net10103),
.Y(net9580)
);

NAND4xp25_ASAP7_75t_R merge9536(
.A(net5306),
.B(net5362),
.C(net468),
.D(net835),
.Y(net9581)
);

NAND4xp75_ASAP7_75t_R merge9537(
.A(net5967),
.B(net5990),
.C(net5062),
.D(net4177),
.Y(net9582)
);

NOR4xp25_ASAP7_75t_R merge9538(
.A(net3007),
.B(net3025),
.C(net2589),
.D(net1709),
.Y(net9583)
);

NOR4xp75_ASAP7_75t_R merge9539(
.A(net5118),
.B(net4985),
.C(net4246),
.D(net3400),
.Y(net9584)
);

O2A1O1Ixp33_ASAP7_75t_R merge9540(
.A1(net2346),
.A2(net2442),
.B(net6195),
.C(net6199),
.Y(net9585)
);

O2A1O1Ixp5_ASAP7_75t_R merge9541(
.A1(net838),
.A2(net4539),
.B(net5162),
.C(net5185),
.Y(net9586)
);

OA211x2_ASAP7_75t_R merge9542(
.A1(net3234),
.A2(net4047),
.B(net6882),
.C(net5928),
.Y(net9587)
);

OA22x2_ASAP7_75t_R merge9543(
.A1(net3176),
.A2(net4229),
.B1(net1631),
.B2(net1635),
.Y(net9588)
);

OA31x2_ASAP7_75t_R merge9544(
.A1(net1605),
.A2(net1592),
.A3(net6940),
.B1(net9711),
.Y(net9589)
);

OAI211xp5_ASAP7_75t_R merge9545(
.A1(net7459),
.A2(net7475),
.B(net220),
.C(net209),
.Y(net9590)
);

OAI22x1_ASAP7_75t_R merge9546(
.A1(net6908),
.A2(net6910),
.B1(net7797),
.B2(net5959),
.Y(net9591)
);

OAI22xp33_ASAP7_75t_R merge9547(
.A1(net5866),
.A2(net7912),
.B1(net6031),
.B2(net5848),
.Y(net9592)
);

OAI22xp5_ASAP7_75t_R merge9548(
.A1(net7758),
.A2(net8603),
.B1(net3243),
.B2(net4077),
.Y(net9593)
);

OAI31xp33_ASAP7_75t_R merge9549(
.A1(net2503),
.A2(net2593),
.A3(net554),
.B(net549),
.Y(net9594)
);

OAI31xp67_ASAP7_75t_R merge9550(
.A1(net5610),
.A2(net1915),
.A3(net3943),
.B(net10115),
.Y(net9595)
);

OR4x1_ASAP7_75t_R merge9551(
.A(net3476),
.B(net2459),
.C(net3948),
.D(net3946),
.Y(net9596)
);

OR4x2_ASAP7_75t_R merge9552(
.A(net5884),
.B(net5821),
.C(net6802),
.D(net6791),
.Y(net9597)
);

A2O1A1Ixp33_ASAP7_75t_R merge9553(
.A1(net3962),
.A2(net3887),
.B(net3781),
.C(net3772),
.Y(net9598)
);

AND4x1_ASAP7_75t_R merge9554(
.A(net197),
.B(net177),
.C(net3124),
.D(net3943),
.Y(net9599)
);

AND4x2_ASAP7_75t_R merge9555(
.A(net5801),
.B(net4867),
.C(net3482),
.D(net3524),
.Y(net9600)
);

AO211x2_ASAP7_75t_R merge9556(
.A1(net5756),
.A2(net5719),
.B(net7390),
.C(net7426),
.Y(net9601)
);

AO22x1_ASAP7_75t_R merge9557(
.A1(net3893),
.A2(net3896),
.B1(net219),
.B2(net203),
.Y(net9602)
);

AO22x2_ASAP7_75t_R merge9558(
.A1(net5661),
.A2(net6545),
.B1(net5820),
.B2(net5853),
.Y(net9603)
);

AO31x2_ASAP7_75t_R merge9559(
.A1(net1730),
.A2(net2589),
.A3(net7159),
.B(net7130),
.Y(net9604)
);

AOI211x1_ASAP7_75t_R merge9560(
.A1(net5028),
.A2(net4978),
.B(net5032),
.C(net9913),
.Y(net9605)
);

AOI211xp5_ASAP7_75t_R merge9561(
.A1(net1663),
.A2(net1737),
.B(net3503),
.C(net2474),
.Y(net9606)
);

AOI22x1_ASAP7_75t_R merge9562(
.A1(net7385),
.A2(net7476),
.B1(net8368),
.B2(net7393),
.Y(net9607)
);

AOI22xp33_ASAP7_75t_R merge9563(
.A1(net3261),
.A2(net3218),
.B1(net4814),
.B2(net4828),
.Y(net9608)
);

AOI22xp5_ASAP7_75t_R merge9564(
.A1(net2494),
.A2(net2577),
.B1(net4880),
.B2(net9806),
.Y(net9609)
);

AOI31xp33_ASAP7_75t_R merge9565(
.A1(net1233),
.A2(net2145),
.A3(net2877),
.B(net6577),
.Y(net9610)
);

AOI31xp67_ASAP7_75t_R merge9566(
.A1(net3003),
.A2(net3992),
.A3(net3808),
.B(net2877),
.Y(net9611)
);

NAND4xp25_ASAP7_75t_R merge9567(
.A(net468),
.B(net1420),
.C(net3291),
.D(net9964),
.Y(net9612)
);

NAND4xp75_ASAP7_75t_R merge9568(
.A(net493),
.B(net468),
.C(net4816),
.D(net4811),
.Y(net9613)
);

NOR4xp25_ASAP7_75t_R merge9569(
.A(net5942),
.B(net6842),
.C(net2076),
.D(net2067),
.Y(net9614)
);

NOR4xp75_ASAP7_75t_R merge9570(
.A(net6701),
.B(net6964),
.C(net5111),
.D(net6168),
.Y(net9615)
);

O2A1O1Ixp33_ASAP7_75t_R merge9571(
.A1(net3463),
.A2(net2600),
.B(net3577),
.C(net3571),
.Y(net9616)
);

O2A1O1Ixp5_ASAP7_75t_R merge9572(
.A1(net4167),
.A2(net3204),
.B(net2017),
.C(net2807),
.Y(net9617)
);

OA211x2_ASAP7_75t_R merge9573(
.A1(net3768),
.A2(net3880),
.B(net2999),
.C(net3919),
.Y(net9618)
);

OA22x2_ASAP7_75t_R merge9574(
.A1(net221),
.A2(net1080),
.B1(net2143),
.B2(net3077),
.Y(net9619)
);

OA31x2_ASAP7_75t_R merge9575(
.A1(net3525),
.A2(net2569),
.A3(net2298),
.B1(net9996),
.Y(net9620)
);

OAI211xp5_ASAP7_75t_R merge9576(
.A1(net4392),
.A2(net2637),
.B(net7699),
.C(net7506),
.Y(net9621)
);

OAI22x1_ASAP7_75t_R merge9577(
.A1(net1976),
.A2(net2018),
.B1(net5712),
.B2(net5704),
.Y(net9622)
);

OAI22xp33_ASAP7_75t_R merge9578(
.A1(net3017),
.A2(net2829),
.B1(net2842),
.B2(net4884),
.Y(net9623)
);

OAI22xp5_ASAP7_75t_R merge9579(
.A1(net1278),
.A2(net1334),
.B1(net6080),
.B2(net7136),
.Y(net9624)
);

OAI31xp33_ASAP7_75t_R merge9580(
.A1(net7968),
.A2(net7893),
.A3(net2638),
.B(net5296),
.Y(net9625)
);

OAI31xp67_ASAP7_75t_R merge9581(
.A1(net6127),
.A2(net6122),
.A3(net8649),
.B(net7759),
.Y(net9626)
);

OR4x1_ASAP7_75t_R merge9582(
.A(net1635),
.B(net2453),
.C(net2455),
.D(net10078),
.Y(net9627)
);

OR4x2_ASAP7_75t_R merge9583(
.A(net1120),
.B(net1108),
.C(net2370),
.D(net1473),
.Y(net9628)
);

A2O1A1Ixp33_ASAP7_75t_R merge9584(
.A1(net6286),
.A2(net6285),
.B(net4955),
.C(net34),
.Y(net9629)
);

AND4x1_ASAP7_75t_R merge9585(
.A(net6792),
.B(net6791),
.C(net8596),
.D(net8366),
.Y(net9630)
);

AND4x2_ASAP7_75t_R merge9586(
.A(net5618),
.B(net2877),
.C(net3817),
.D(net3769),
.Y(net9631)
);

AO211x2_ASAP7_75t_R merge9587(
.A1(net4710),
.A2(net5636),
.B(net3793),
.C(net6505),
.Y(net9632)
);

NAND2x1_ASAP7_75t_R merge9588(
.A(net3188),
.B(net3206),
.Y(net9633)
);

ICGx5_ASAP7_75t_R merge9589(
.ENA(net3387),
.SE(net3401),
.CLK(clk),
.GCLK(net9634)
);

NAND2x1p5_ASAP7_75t_R merge9590(
.A(net1335),
.B(net1369),
.Y(net9635)
);

ICGx5p33DC_ASAP7_75t_R merge9591(
.ENA(net405),
.SE(net431),
.CLK(clk),
.GCLK(net9636)
);

ICGx6p67DC_ASAP7_75t_R merge9592(
.ENA(net7325),
.SE(net7356),
.CLK(clk),
.GCLK(net9637)
);

ICGx8DC_ASAP7_75t_R merge9593(
.ENA(net8209),
.SE(net8250),
.CLK(clk),
.GCLK(net9638)
);

ICGx1_ASAP7_75t_R merge9594(
.ENA(net8837),
.SE(net8829),
.CLK(clk),
.GCLK(net9639)
);

ICGx2_ASAP7_75t_R merge9595(
.ENA(net7738),
.SE(net7768),
.CLK(clk),
.GCLK(net9640)
);

ICGx2p67DC_ASAP7_75t_R merge9596(
.ENA(net5388),
.SE(net5430),
.CLK(clk),
.GCLK(net9641)
);

ICGx3_ASAP7_75t_R merge9597(
.ENA(net7479),
.SE(net7483),
.CLK(clk),
.GCLK(net9642)
);

NAND2x2_ASAP7_75t_R merge9598(
.A(net1624),
.B(net1636),
.Y(net9643)
);

ICGx4DC_ASAP7_75t_R merge9599(
.ENA(net2443),
.SE(net2458),
.CLK(clk),
.GCLK(net9644)
);

NAND2xp33_ASAP7_75t_R merge9600(
.A(net4126),
.B(net4127),
.Y(net9645)
);

NAND2xp5_ASAP7_75t_R merge9601(
.A(net7888),
.B(net7949),
.Y(net9646)
);

ICGx4_ASAP7_75t_R merge9602(
.ENA(net3526),
.SE(net3583),
.CLK(clk),
.GCLK(net9647)
);

ICGx5_ASAP7_75t_R merge9603(
.ENA(net302),
.GCLK(net308),
.CLK(clk)
);

ICGx5p33DC_ASAP7_75t_R merge9604(
.ENA(net1841),
.SE(net1855),
.CLK(clk),
.GCLK(net9649)
);

ICGx6p67DC_ASAP7_75t_R merge9605(
.ENA(net62),
.SE(net93),
.CLK(clk),
.GCLK(net9650)
);

ICGx8DC_ASAP7_75t_R merge9606(
.ENA(net2695),
.SE(net2749),
.CLK(clk),
.GCLK(net9651)
);

ICGx1_ASAP7_75t_R merge9607(
.ENA(net1169),
.SE(net1176),
.CLK(clk),
.GCLK(net9652)
);

NAND2xp67_ASAP7_75t_R merge9608(
.A(net704),
.B(net729),
.Y(net9653)
);

ICGx2_ASAP7_75t_R merge9609(
.ENA(net8676),
.SE(net8757),
.CLK(clk),
.GCLK(net9654)
);

NOR2x1_ASAP7_75t_R merge9610(
.A(net8143),
.B(net8176),
.Y(net9655)
);

ICGx2p67DC_ASAP7_75t_R merge9611(
.ENA(net5228),
.SE(net5241),
.CLK(clk),
.GCLK(net9656)
);

ICGx3_ASAP7_75t_R merge9612(
.ENA(net811),
.SE(net772),
.CLK(clk),
.GCLK(net9657)
);

ICGx4DC_ASAP7_75t_R merge9613(
.ENA(net7389),
.SE(net7381),
.CLK(clk),
.GCLK(net9658)
);

ICGx4_ASAP7_75t_R merge9614(
.ENA(net8328),
.GCLK(net8332),
.CLK(clk)
);

ICGx5_ASAP7_75t_R merge9615(
.ENA(net6518),
.SE(net9297),
.CLK(clk),
.GCLK(net9660)
);

ICGx5p33DC_ASAP7_75t_R merge9616(
.ENA(net8671),
.SE(net8655),
.CLK(clk),
.GCLK(net9661)
);

ICGx6p67DC_ASAP7_75t_R merge9617(
.ENA(net8041),
.SE(net8107),
.CLK(clk),
.GCLK(net9662)
);

ICGx8DC_ASAP7_75t_R merge9618(
.ENA(net4815),
.SE(net4822),
.CLK(clk),
.GCLK(net9663)
);

NOR2x1p5_ASAP7_75t_R merge9619(
.A(net4199),
.B(net4265),
.Y(net9664)
);

ICGx1_ASAP7_75t_R merge9620(
.ENA(net5587),
.SE(net5594),
.CLK(clk),
.GCLK(net9665)
);

ICGx2_ASAP7_75t_R merge9621(
.ENA(net828),
.SE(net867),
.CLK(clk),
.GCLK(net9666)
);

ICGx2p67DC_ASAP7_75t_R merge9622(
.ENA(net7562),
.SE(net7568),
.CLK(clk),
.GCLK(net9667)
);

NOR2x2_ASAP7_75t_R merge9623(
.A(net1820),
.B(net1751),
.Y(net9668)
);

NOR2xp33_ASAP7_75t_R merge9624(
.A(net620),
.B(net642),
.Y(net9669)
);

ICGx3_ASAP7_75t_R merge9625(
.ENA(net4972),
.SE(net4975),
.CLK(clk),
.GCLK(net9670)
);

ICGx4DC_ASAP7_75t_R merge9626(
.ENA(net7129),
.SE(net7156),
.CLK(clk),
.GCLK(net9671)
);

ICGx4_ASAP7_75t_R merge9627(
.ENA(net5155),
.SE(net5174),
.CLK(clk),
.GCLK(net9672)
);

NOR2xp67_ASAP7_75t_R merge9628(
.A(net8917),
.B(net8915),
.Y(net9673)
);

OR2x2_ASAP7_75t_R merge9629(
.A(net2005),
.B(net2008),
.Y(net9674)
);

ICGx5_ASAP7_75t_R merge9630(
.ENA(net6633),
.SE(net6661),
.CLK(clk),
.GCLK(net9675)
);

OR2x4_ASAP7_75t_R merge9631(
.A(net6716),
.B(net6784),
.Y(net9676)
);

ICGx5p33DC_ASAP7_75t_R merge9632(
.ENA(net5619),
.SE(net5690),
.CLK(clk),
.GCLK(net9677)
);

ICGx6p67DC_ASAP7_75t_R merge9633(
.ENA(net6054),
.SE(net6115),
.CLK(clk),
.GCLK(net9678)
);

ICGx8DC_ASAP7_75t_R merge9634(
.ENA(net2510),
.SE(net2513),
.CLK(clk),
.GCLK(net9679)
);

OR2x6_ASAP7_75t_R merge9635(
.A(net3299),
.B(net3302),
.Y(net9680)
);

ICGx1_ASAP7_75t_R merge9636(
.ENA(net377),
.SE(net378),
.CLK(clk),
.GCLK(net9681)
);

ICGx2_ASAP7_75t_R merge9637(
.ENA(net9118),
.SE(net9298),
.CLK(clk),
.GCLK(net9682)
);

ICGx2p67DC_ASAP7_75t_R merge9638(
.ENA(net1739),
.SE(net1689),
.CLK(clk),
.GCLK(net9683)
);

ICGx3_ASAP7_75t_R merge9639(
.ENA(net4771),
.SE(net4739),
.CLK(clk),
.GCLK(net9684)
);

ICGx4DC_ASAP7_75t_R merge9640(
.ENA(net4557),
.SE(net4588),
.CLK(clk),
.GCLK(net9685)
);

ICGx4_ASAP7_75t_R merge9641(
.ENA(net7999),
.SE(net7995),
.CLK(clk),
.GCLK(net9686)
);

ICGx5_ASAP7_75t_R merge9642(
.ENA(net8930),
.SE(net9009),
.CLK(clk),
.GCLK(net9687)
);

ICGx5p33DC_ASAP7_75t_R merge9643(
.ENA(net9011),
.SE(net9084),
.CLK(clk),
.GCLK(net9688)
);

ICGx6p67DC_ASAP7_75t_R merge9644(
.ENA(net7845),
.SE(net7866),
.CLK(clk),
.GCLK(net9689)
);

ICGx8DC_ASAP7_75t_R merge9645(
.ENA(net5956),
.SE(net5987),
.CLK(clk),
.GCLK(net9690)
);

XNOR2x1_ASAP7_75t_R merge9646(
.B(net3479),
.A(net3501),
.Y(net9691)
);

XNOR2x2_ASAP7_75t_R merge9647(
.A(net1414),
.B(net1471),
.Y(net9692)
);

ICGx1_ASAP7_75t_R merge9648(
.ENA(net2922),
.SE(net2968),
.CLK(clk),
.GCLK(net9693)
);

XNOR2xp5_ASAP7_75t_R merge9649(
.A(net5904),
.B(net5924),
.Y(net9694)
);

XOR2x1_ASAP7_75t_R merge9650(
.A(net3956),
.B(net3961),
.Y(net9695)
);

ICGx2_ASAP7_75t_R merge9651(
.ENA(net4359),
.SE(net4436),
.CLK(clk),
.GCLK(net9696)
);

ICGx2p67DC_ASAP7_75t_R merge9652(
.ENA(net4488),
.SE(net4489),
.CLK(clk),
.GCLK(net9697)
);

ICGx3_ASAP7_75t_R merge9653(
.ENA(net6549),
.SE(net6562),
.CLK(clk),
.GCLK(net9698)
);

XOR2x2_ASAP7_75t_R merge9654(
.A(net6235),
.B(net6259),
.Y(net9699)
);

XOR2xp5_ASAP7_75t_R merge9655(
.A(net7676),
.B(net7682),
.Y(net9700)
);

AND2x2_ASAP7_75t_R merge9656(
.A(net2628),
.B(net2644),
.Y(net9701)
);

ICGx4DC_ASAP7_75t_R merge9657(
.ENA(net1965),
.SE(net1992),
.CLK(clk),
.GCLK(net9702)
);

AND2x4_ASAP7_75t_R merge9658(
.A(net4886),
.B(net4892),
.Y(net9703)
);

ICGx4_ASAP7_75t_R merge9659(
.ENA(net972),
.SE(net973),
.CLK(clk),
.GCLK(net9704)
);

ICGx5_ASAP7_75t_R merge9660(
.ENA(net8525),
.SE(net8584),
.CLK(clk),
.GCLK(net9705)
);

ICGx5p33DC_ASAP7_75t_R merge9661(
.ENA(net8429),
.SE(net8491),
.CLK(clk),
.GCLK(net9706)
);

ICGx6p67DC_ASAP7_75t_R merge9662(
.ENA(net5453),
.SE(net5465),
.CLK(clk),
.GCLK(net9707)
);

ICGx8DC_ASAP7_75t_R merge9663(
.ENA(net6317),
.SE(net6327),
.CLK(clk),
.GCLK(net9708)
);

ICGx1_ASAP7_75t_R merge9664(
.ENA(net4030),
.SE(net4037),
.CLK(clk),
.GCLK(net9709)
);

ICGx2_ASAP7_75t_R merge9665(
.ENA(net5280),
.SE(net5301),
.CLK(clk),
.GCLK(net9710)
);

ICGx2p67DC_ASAP7_75t_R merge9666(
.ENA(net6896),
.SE(net6921),
.CLK(clk),
.GCLK(net9711)
);

ICGx3_ASAP7_75t_R merge9667(
.ENA(net205),
.SE(net211),
.CLK(clk),
.GCLK(net9712)
);

ICGx4DC_ASAP7_75t_R merge9668(
.ENA(net3684),
.SE(net3688),
.CLK(clk),
.GCLK(net9713)
);

AND2x6_ASAP7_75t_R merge9669(
.A(net5826),
.B(net5845),
.Y(net9714)
);

HAxp5_ASAP7_75t_R merge9670(
.A(net6985),
.B(net6984),
.CON(net9715)
);

NAND2x1_ASAP7_75t_R merge9671(
.A(net1535),
.B(net1541),
.Y(net9716)
);

ICGx4_ASAP7_75t_R merge9672(
.ENA(net2834),
.SE(net2799),
.CLK(clk),
.GCLK(net9717)
);

NAND2x1p5_ASAP7_75t_R merge9673(
.A(net7040),
.B(net7048),
.Y(net9718)
);

ICGx5_ASAP7_75t_R merge9674(
.ENA(net5760),
.SE(net5765),
.CLK(clk),
.GCLK(net9719)
);

ICGx5p33DC_ASAP7_75t_R merge9675(
.ENA(net7242),
.SE(net7244),
.CLK(clk),
.GCLK(net9720)
);

NAND2x2_ASAP7_75t_R merge9676(
.A(net3101),
.B(net3172),
.Y(net9721)
);

ICGx6p67DC_ASAP7_75t_R merge9677(
.ENA(net6139),
.SE(net6185),
.CLK(clk),
.GCLK(net9722)
);

NAND2xp33_ASAP7_75t_R merge9678(
.A(net2085),
.B(net2118),
.Y(net9723)
);

NAND2xp5_ASAP7_75t_R merge9679(
.A(net3904),
.B(net3865),
.Y(net9724)
);

ICGx8DC_ASAP7_75t_R merge9680(
.ENA(net2856),
.SE(net2872),
.CLK(clk),
.GCLK(net9725)
);

ICGx1_ASAP7_75t_R merge9681(
.ENA(net2266),
.SE(net2254),
.CLK(clk),
.GCLK(net9726)
);

ICGx2_ASAP7_75t_R merge9682(
.ENA(net4669),
.SE(net4674),
.CLK(clk),
.GCLK(net9727)
);

NAND2xp67_ASAP7_75t_R merge9683(
.A(net1141),
.B(net1143),
.Y(net9728)
);

ICGx2p67DC_ASAP7_75t_R merge9684(
.ENA(net3775),
.SE(net3795),
.CLK(clk),
.GCLK(net9729)
);

NOR2x1_ASAP7_75t_R merge9685(
.A(net991),
.B(net1063),
.Y(net9730)
);

ICGx3_ASAP7_75t_R merge9686(
.ENA(net6799),
.SE(net6841),
.CLK(clk),
.GCLK(net9731)
);

NOR2x1p5_ASAP7_75t_R merge9687(
.A(net3031),
.B(net3019),
.Y(net9732)
);

ICGx4DC_ASAP7_75t_R merge9688(
.ENA(net3601),
.SE(net3597),
.CLK(clk),
.GCLK(net9733)
);

NOR2x2_ASAP7_75t_R merge9689(
.A(net5050),
.B(net5107),
.Y(net9734)
);

ICGx4_ASAP7_75t_R merge9690(
.ENA(net4270),
.SE(net4295),
.CLK(clk),
.GCLK(net9735)
);

ICGx5_ASAP7_75t_R merge9691(
.ENA(net6415),
.SE(net6440),
.CLK(clk),
.GCLK(net9736)
);

ICGx5p33DC_ASAP7_75t_R merge9692(
.ENA(net8362),
.SE(net8417),
.CLK(clk),
.GCLK(net9737)
);

ICGx6p67DC_ASAP7_75t_R merge9693(
.ENA(net518),
.SE(net521),
.CLK(clk),
.GCLK(net9738)
);

NOR2xp33_ASAP7_75t_R merge9694(
.A(net1276),
.B(net1286),
.Y(net9739)
);

NOR2xp67_ASAP7_75t_R merge9695(
.A(net2189),
.B(net2206),
.Y(net9740)
);

ICGx8DC_ASAP7_75t_R merge9696(
.ENA(net3826),
.SE(net2987),
.CLK(clk),
.GCLK(net9741)
);

OR2x2_ASAP7_75t_R merge9697(
.A(net4250),
.B(net3225),
.Y(net9742)
);

ICGx1_ASAP7_75t_R merge9698(
.ENA(net9033),
.SE(net9076),
.CLK(clk),
.GCLK(net9743)
);

ICGx2_ASAP7_75t_R merge9699(
.ENA(net1908),
.SE(net1049),
.CLK(clk),
.GCLK(net9744)
);

ICGx2p67DC_ASAP7_75t_R merge9700(
.ENA(net4007),
.SE(net3841),
.CLK(clk),
.GCLK(net9745)
);

ICGx3_ASAP7_75t_R merge9701(
.ENA(net1144),
.SE(net9525),
.CLK(clk),
.GCLK(net9746)
);

ICGx4DC_ASAP7_75t_R merge9702(
.ENA(net1566),
.SE(net1560),
.CLK(clk),
.GCLK(net9747)
);

ICGx4_ASAP7_75t_R merge9703(
.ENA(net1880),
.SE(net1903),
.CLK(clk),
.GCLK(net9748)
);

OR2x4_ASAP7_75t_R merge9704(
.A(net2500),
.B(net1465),
.Y(net9749)
);

OR2x6_ASAP7_75t_R merge9705(
.A(net3569),
.B(net2662),
.Y(net9750)
);

XNOR2x1_ASAP7_75t_R merge9706(
.B(net1440),
.A(net1487),
.Y(net9751)
);

ICGx5_ASAP7_75t_R merge9707(
.ENA(net985),
.SE(net9730),
.CLK(clk),
.GCLK(net9752)
);

XNOR2x2_ASAP7_75t_R merge9708(
.A(net3088),
.B(net2150),
.Y(net9753)
);

ICGx5p33DC_ASAP7_75t_R merge9709(
.ENA(net4519),
.SE(net4590),
.CLK(clk),
.GCLK(net9754)
);

XNOR2xp5_ASAP7_75t_R merge9710(
.A(net3236),
.B(net3038),
.Y(net9755)
);

ICGx6p67DC_ASAP7_75t_R merge9711(
.ENA(net1862),
.SE(net2916),
.CLK(clk),
.GCLK(net9756)
);

ICGx8DC_ASAP7_75t_R merge9712(
.ENA(net8128),
.SE(net8145),
.CLK(clk),
.GCLK(net9757)
);

ICGx1_ASAP7_75t_R merge9713(
.ENA(net3690),
.SE(net3843),
.CLK(clk),
.GCLK(net9758)
);

ICGx2_ASAP7_75t_R merge9714(
.ENA(net7940),
.SE(net8036),
.CLK(clk),
.GCLK(net9759)
);

ICGx2p67DC_ASAP7_75t_R merge9715(
.ENA(net9047),
.SE(net8227),
.CLK(clk),
.GCLK(out4)
);

ICGx3_ASAP7_75t_R merge9716(
.ENA(net7089),
.SE(net6946),
.CLK(clk),
.GCLK(net9760)
);

ICGx4DC_ASAP7_75t_R merge9717(
.ENA(net8017),
.SE(net8090),
.CLK(clk),
.GCLK(net9761)
);

ICGx4_ASAP7_75t_R merge9718(
.ENA(net7313),
.SE(net8125),
.CLK(clk),
.GCLK(net9762)
);

ICGx5_ASAP7_75t_R merge9719(
.ENA(net3338),
.SE(net3230),
.CLK(clk),
.GCLK(net9763)
);

ICGx5p33DC_ASAP7_75t_R merge9720(
.ENA(net3268),
.SE(net2329),
.CLK(clk),
.GCLK(net9764)
);

XOR2x1_ASAP7_75t_R merge9721(
.A(net3998),
.B(net2129),
.Y(net9765)
);

ICGx6p67DC_ASAP7_75t_R merge9722(
.ENA(net5626),
.SE(net6606),
.CLK(clk),
.GCLK(net9766)
);

XOR2x2_ASAP7_75t_R merge9723(
.A(net6726),
.B(net6785),
.Y(net9767)
);

XOR2xp5_ASAP7_75t_R merge9724(
.A(net2146),
.B(net3040),
.Y(net9768)
);

ICGx8DC_ASAP7_75t_R merge9725(
.ENA(net6780),
.SE(net6745),
.CLK(clk),
.GCLK(net9769)
);

AND2x2_ASAP7_75t_R merge9726(
.A(net2247),
.B(net3332),
.Y(net9770)
);

AND2x4_ASAP7_75t_R merge9727(
.A(net3762),
.B(net4767),
.Y(net9771)
);

ICGx1_ASAP7_75t_R merge9728(
.ENA(net3670),
.SE(net4537),
.CLK(clk),
.GCLK(net9772)
);

ICGx2_ASAP7_75t_R merge9729(
.ENA(net7278),
.SE(net7303),
.CLK(clk),
.GCLK(net9773)
);

ICGx2p67DC_ASAP7_75t_R merge9730(
.ENA(net7714),
.SE(net8560),
.CLK(clk),
.GCLK(net9774)
);

ICGx3_ASAP7_75t_R merge9731(
.ENA(net5083),
.SE(net4334),
.CLK(clk),
.GCLK(net9775)
);

ICGx4DC_ASAP7_75t_R merge9732(
.ENA(net5665),
.SE(net7448),
.CLK(clk),
.GCLK(net9776)
);

ICGx4_ASAP7_75t_R merge9733(
.ENA(net4927),
.SE(net4085),
.CLK(clk),
.GCLK(net9777)
);

ICGx5_ASAP7_75t_R merge9734(
.ENA(net7773),
.SE(net6850),
.CLK(clk),
.GCLK(net9778)
);

ICGx5p33DC_ASAP7_75t_R merge9735(
.ENA(net6445),
.SE(net5433),
.CLK(clk),
.GCLK(net9779)
);

AND2x6_ASAP7_75t_R merge9736(
.A(net7024),
.B(net7897),
.Y(net9780)
);

HAxp5_ASAP7_75t_R merge9737(
.A(net2041),
.B(net1231),
.CON(net9781)
);

ICGx6p67DC_ASAP7_75t_R merge9738(
.ENA(net1801),
.SE(net1812),
.CLK(clk),
.GCLK(net9782)
);

ICGx8DC_ASAP7_75t_R merge9739(
.ENA(net450),
.SE(net1405),
.CLK(clk),
.GCLK(net9783)
);

NAND2x1_ASAP7_75t_R merge9740(
.A(net2300),
.B(net2170),
.Y(net9784)
);

ICGx1_ASAP7_75t_R merge9741(
.ENA(net8448),
.SE(net7599),
.CLK(clk),
.GCLK(net9785)
);

ICGx2_ASAP7_75t_R merge9742(
.ENA(net3828),
.SE(net3807),
.CLK(clk),
.GCLK(net9786)
);

ICGx2p67DC_ASAP7_75t_R merge9743(
.ENA(net8771),
.SE(net8839),
.CLK(clk),
.GCLK(net9787)
);

ICGx3_ASAP7_75t_R merge9744(
.ENA(net5008),
.SE(net3158),
.CLK(clk),
.GCLK(net9788)
);

ICGx4DC_ASAP7_75t_R merge9745(
.ENA(net7691),
.SE(net8415),
.CLK(clk),
.GCLK(net9789)
);

ICGx4_ASAP7_75t_R merge9746(
.ENA(net7091),
.SE(net5342),
.CLK(clk),
.GCLK(net9790)
);

ICGx5_ASAP7_75t_R merge9747(
.ENA(net1804),
.SE(net896),
.CLK(clk),
.GCLK(net9791)
);

NAND2x1p5_ASAP7_75t_R merge9748(
.A(net1793),
.B(net889),
.Y(net9792)
);

NAND2x2_ASAP7_75t_R merge9749(
.A(net2211),
.B(net2246),
.Y(net9793)
);

ICGx5p33DC_ASAP7_75t_R merge9750(
.ENA(net4531),
.SE(net6397),
.CLK(clk),
.GCLK(net9794)
);

ICGx6p67DC_ASAP7_75t_R merge9751(
.ENA(net4342),
.SE(net4366),
.CLK(clk),
.GCLK(net9795)
);

NAND2xp33_ASAP7_75t_R merge9752(
.A(net1226),
.B(net2050),
.Y(net9796)
);

NAND2xp5_ASAP7_75t_R merge9753(
.A(net2542),
.B(net2583),
.Y(net9797)
);

NAND2xp67_ASAP7_75t_R merge9754(
.A(net8028),
.B(net6360),
.Y(net9798)
);

NOR2x1_ASAP7_75t_R merge9755(
.A(net1444),
.B(net1394),
.Y(net9799)
);

ICGx8DC_ASAP7_75t_R merge9756(
.ENA(net8416),
.SE(net6617),
.CLK(clk),
.GCLK(net9800)
);

ICGx1_ASAP7_75t_R merge9757(
.ENA(net2704),
.SE(net2741),
.CLK(clk),
.GCLK(net9801)
);

ICGx2_ASAP7_75t_R merge9758(
.ENA(net6028),
.SE(net6077),
.CLK(clk),
.GCLK(net9802)
);

NOR2x1p5_ASAP7_75t_R merge9759(
.A(net2051),
.B(net1318),
.Y(net9803)
);

NOR2x2_ASAP7_75t_R merge9760(
.A(net7201),
.B(net7105),
.Y(net9804)
);

ICGx2p67DC_ASAP7_75t_R merge9761(
.ENA(net3613),
.SE(net4415),
.CLK(clk),
.GCLK(net9805)
);

ICGx3_ASAP7_75t_R merge9762(
.ENA(net3973),
.SE(net4012),
.CLK(clk),
.GCLK(net9806)
);

ICGx4DC_ASAP7_75t_R merge9763(
.ENA(net4744),
.SE(net3928),
.CLK(clk),
.GCLK(net9807)
);

NOR2xp33_ASAP7_75t_R merge9764(
.A(net4301),
.B(net6039),
.Y(net9808)
);

NOR2xp67_ASAP7_75t_R merge9765(
.A(net5073),
.B(net4909),
.Y(net9809)
);

OR2x2_ASAP7_75t_R merge9766(
.A(net4421),
.B(net2535),
.Y(net9810)
);

ICGx4_ASAP7_75t_R merge9767(
.ENA(net6105),
.SE(net5098),
.CLK(clk),
.GCLK(net9811)
);

ICGx5_ASAP7_75t_R merge9768(
.ENA(net895),
.SE(net1819),
.CLK(clk),
.GCLK(net9812)
);

ICGx5p33DC_ASAP7_75t_R merge9769(
.ENA(net2496),
.SE(net3333),
.CLK(clk),
.GCLK(net9813)
);

ICGx6p67DC_ASAP7_75t_R merge9770(
.ENA(net8163),
.SE(net8142),
.CLK(clk),
.GCLK(net9814)
);

ICGx8DC_ASAP7_75t_R merge9771(
.ENA(net4602),
.SE(net6261),
.CLK(clk),
.GCLK(net9815)
);

OR2x4_ASAP7_75t_R merge9772(
.A(net5989),
.B(net6741),
.Y(net9816)
);

ICGx1_ASAP7_75t_R merge9773(
.ENA(net8334),
.SE(net8412),
.CLK(clk),
.GCLK(net9817)
);

ICGx2_ASAP7_75t_R merge9774(
.ENA(net6568),
.SE(net7536),
.CLK(clk),
.GCLK(net9818)
);

ICGx2p67DC_ASAP7_75t_R merge9775(
.ENA(net8810),
.SE(net8040),
.CLK(clk),
.GCLK(net9819)
);

OR2x6_ASAP7_75t_R merge9776(
.A(net7870),
.B(net8639),
.Y(net9820)
);

ICGx3_ASAP7_75t_R merge9777(
.ENA(net2059),
.SE(net2906),
.CLK(clk),
.GCLK(net9821)
);

XNOR2x1_ASAP7_75t_R merge9778(
.B(net4311),
.A(net5351),
.Y(net9822)
);

ICGx4DC_ASAP7_75t_R merge9779(
.ENA(net6345),
.SE(net6120),
.CLK(clk),
.GCLK(net9823)
);

XNOR2x2_ASAP7_75t_R merge9780(
.A(net4388),
.B(net2565),
.Y(net9824)
);

ICGx4_ASAP7_75t_R merge9781(
.ENA(net1209),
.SE(net9334),
.CLK(clk),
.GCLK(net9825)
);

ICGx5_ASAP7_75t_R merge9782(
.ENA(net6739),
.SE(net5861),
.CLK(clk),
.GCLK(net9826)
);

ICGx5p33DC_ASAP7_75t_R merge9783(
.ENA(net6574),
.SE(net4748),
.CLK(clk),
.GCLK(net9827)
);

ICGx6p67DC_ASAP7_75t_R merge9784(
.ENA(net386),
.SE(net9234),
.CLK(clk),
.GCLK(net9828)
);

XNOR2xp5_ASAP7_75t_R merge9785(
.A(net3043),
.B(net3084),
.Y(net9829)
);

ICGx8DC_ASAP7_75t_R merge9786(
.ENA(net6609),
.SE(net8411),
.CLK(clk),
.GCLK(net9830)
);

ICGx1_ASAP7_75t_R merge9787(
.ENA(net6449),
.SE(net7254),
.CLK(clk),
.GCLK(net9831)
);

ICGx2_ASAP7_75t_R merge9788(
.ENA(net1377),
.SE(net1305),
.CLK(clk),
.GCLK(net9832)
);

XOR2x1_ASAP7_75t_R merge9789(
.A(net6953),
.B(net8662),
.Y(net9833)
);

XOR2x2_ASAP7_75t_R merge9790(
.A(net8500),
.B(net8617),
.Y(net9834)
);

ICGx2p67DC_ASAP7_75t_R merge9791(
.ENA(net5261),
.SE(net6073),
.CLK(clk),
.GCLK(net9835)
);

ICGx3_ASAP7_75t_R merge9792(
.ENA(net4555),
.SE(net5470),
.CLK(clk),
.GCLK(net9836)
);

XOR2xp5_ASAP7_75t_R merge9793(
.A(net8650),
.B(net6923),
.Y(net9837)
);

AND2x2_ASAP7_75t_R merge9794(
.A(net1442),
.B(net1469),
.Y(net9838)
);

AND2x4_ASAP7_75t_R merge9795(
.A(net4929),
.B(net4008),
.Y(net9839)
);

AND2x6_ASAP7_75t_R merge9796(
.A(net6023),
.B(net4979),
.Y(net9840)
);

ICGx4DC_ASAP7_75t_R merge9797(
.ENA(net6720),
.SE(net7590),
.CLK(clk),
.GCLK(net9841)
);

ICGx4_ASAP7_75t_R merge9798(
.ENA(net3579),
.SE(net2579),
.CLK(clk),
.GCLK(net9842)
);

ICGx5_ASAP7_75t_R merge9799(
.ENA(net8147),
.SE(net8189),
.CLK(clk),
.GCLK(net9843)
);

ICGx5p33DC_ASAP7_75t_R merge9800(
.ENA(net2123),
.SE(net2330),
.CLK(clk),
.GCLK(net9844)
);

ICGx6p67DC_ASAP7_75t_R merge9801(
.ENA(net4833),
.SE(net6753),
.CLK(clk),
.GCLK(net9845)
);

HAxp5_ASAP7_75t_R merge9802(
.A(net4823),
.B(net5944),
.CON(net9846)
);

ICGx8DC_ASAP7_75t_R merge9803(
.ENA(net8904),
.SE(net7274),
.CLK(clk),
.GCLK(net9847)
);

NAND2x1_ASAP7_75t_R merge9804(
.A(net7785),
.B(net7694),
.Y(net9848)
);

ICGx1_ASAP7_75t_R merge9805(
.ENA(net1894),
.SE(net1930),
.CLK(clk),
.GCLK(net9849)
);

NAND2x1p5_ASAP7_75t_R merge9806(
.A(net7613),
.B(net6687),
.Y(net9850)
);

ICGx2_ASAP7_75t_R merge9807(
.ENA(net8707),
.SE(net8724),
.CLK(clk),
.GCLK(net9851)
);

ICGx2p67DC_ASAP7_75t_R merge9808(
.ENA(net9007),
.SE(net6395),
.CLK(clk),
.GCLK(net9852)
);

NAND2x2_ASAP7_75t_R merge9809(
.A(net4903),
.B(net4242),
.Y(net9853)
);

ICGx3_ASAP7_75t_R merge9810(
.ENA(net2278),
.SE(net1542),
.CLK(clk),
.GCLK(net9854)
);

ICGx4DC_ASAP7_75t_R merge9811(
.ENA(net4331),
.SE(net3422),
.CLK(clk),
.GCLK(net9855)
);

ICGx4_ASAP7_75t_R merge9812(
.ENA(net1790),
.SE(net3664),
.CLK(clk),
.GCLK(net9856)
);

ICGx5_ASAP7_75t_R merge9813(
.ENA(net3749),
.SE(net3748),
.CLK(clk),
.GCLK(net9857)
);

ICGx5p33DC_ASAP7_75t_R merge9814(
.ENA(net2728),
.SE(net4578),
.CLK(clk),
.GCLK(net9858)
);

ICGx6p67DC_ASAP7_75t_R merge9815(
.ENA(net5074),
.SE(net7037),
.CLK(clk),
.GCLK(net9859)
);

ICGx8DC_ASAP7_75t_R merge9816(
.ENA(net4005),
.SE(net3090),
.CLK(clk),
.GCLK(net9860)
);

NAND2xp33_ASAP7_75t_R merge9817(
.A(net5768),
.B(net8436),
.Y(net9861)
);

ICGx1_ASAP7_75t_R merge9818(
.ENA(net5640),
.SE(net5682),
.CLK(clk),
.GCLK(net9862)
);

ICGx2_ASAP7_75t_R merge9819(
.ENA(net7035),
.SE(net8577),
.CLK(clk),
.GCLK(net9863)
);

ICGx2p67DC_ASAP7_75t_R merge9820(
.ENA(net9388),
.SE(net9599),
.CLK(clk),
.GCLK(net9864)
);

NAND2xp5_ASAP7_75t_R merge9821(
.A(net6686),
.B(net6698),
.Y(net9865)
);

NAND2xp67_ASAP7_75t_R merge9822(
.A(net8466),
.B(net7598),
.Y(net9866)
);

ICGx3_ASAP7_75t_R merge9823(
.ENA(net7703),
.SE(net6768),
.CLK(clk),
.GCLK(net9867)
);

ICGx4DC_ASAP7_75t_R merge9824(
.ENA(net4162),
.SE(net4006),
.CLK(clk),
.GCLK(net9868)
);

ICGx4_ASAP7_75t_R merge9825(
.ENA(net4504),
.SE(net4381),
.CLK(clk),
.GCLK(net9869)
);

ICGx5_ASAP7_75t_R merge9826(
.ENA(net4708),
.SE(net4854),
.CLK(clk),
.GCLK(net9870)
);

ICGx5p33DC_ASAP7_75t_R merge9827(
.ENA(net5482),
.SE(net3606),
.CLK(clk),
.GCLK(net9871)
);

NOR2x1_ASAP7_75t_R merge9828(
.A(net4848),
.B(net5020),
.Y(net9872)
);

NOR2x1p5_ASAP7_75t_R merge9829(
.A(net5850),
.B(net4922),
.Y(net9873)
);

NOR2x2_ASAP7_75t_R merge9830(
.A(net3516),
.B(net3238),
.Y(net9874)
);

ICGx6p67DC_ASAP7_75t_R merge9831(
.ENA(net8793),
.SE(net8641),
.CLK(clk),
.GCLK(net9875)
);

ICGx8DC_ASAP7_75t_R merge9832(
.ENA(net7701),
.SE(net4919),
.CLK(clk),
.GCLK(net9876)
);

ICGx1_ASAP7_75t_R merge9833(
.ENA(net8172),
.SE(net8958),
.CLK(clk),
.GCLK(net9877)
);

NOR2xp33_ASAP7_75t_R merge9834(
.A(net2223),
.B(net2216),
.Y(net9878)
);

NOR2xp67_ASAP7_75t_R merge9835(
.A(net8985),
.B(net9008),
.Y(net9879)
);

OR2x2_ASAP7_75t_R merge9836(
.A(net5268),
.B(net6017),
.Y(net9880)
);

ICGx2_ASAP7_75t_R merge9837(
.ENA(net6729),
.SE(net6735),
.CLK(clk),
.GCLK(net9881)
);

ICGx2p67DC_ASAP7_75t_R merge9838(
.ENA(net7946),
.SE(net6182),
.CLK(clk),
.GCLK(net9882)
);

OR2x4_ASAP7_75t_R merge9839(
.A(net8472),
.B(net8407),
.Y(net9883)
);

ICGx3_ASAP7_75t_R merge9840(
.ENA(net5684),
.SE(net5997),
.CLK(clk),
.GCLK(net9884)
);

OR2x6_ASAP7_75t_R merge9841(
.A(net8453),
.B(net8651),
.Y(net9885)
);

ICGx4DC_ASAP7_75t_R merge9842(
.ENA(net8547),
.SE(net8624),
.CLK(clk),
.GCLK(net9886)
);

XNOR2x1_ASAP7_75t_R merge9843(
.B(net4998),
.A(net4254),
.Y(net9887)
);

ICGx4_ASAP7_75t_R merge9844(
.ENA(net1765),
.SE(net1786),
.CLK(clk),
.GCLK(net9888)
);

ICGx5_ASAP7_75t_R merge9845(
.ENA(net1975),
.SE(net9220),
.CLK(clk),
.GCLK(net9889)
);

XNOR2x2_ASAP7_75t_R merge9846(
.A(net4187),
.B(net4094),
.Y(net9890)
);

XNOR2xp5_ASAP7_75t_R merge9847(
.A(net8905),
.B(net8194),
.Y(net9891)
);

ICGx5p33DC_ASAP7_75t_R merge9848(
.ENA(net8204),
.SE(net4597),
.CLK(clk),
.GCLK(net9892)
);

ICGx6p67DC_ASAP7_75t_R merge9849(
.ENA(net6417),
.SE(net6431),
.CLK(clk),
.GCLK(net9893)
);

ICGx8DC_ASAP7_75t_R merge9850(
.ENA(net8032),
.SE(net8104),
.CLK(clk),
.GCLK(net9894)
);

ICGx1_ASAP7_75t_R merge9851(
.ENA(net5491),
.SE(net8184),
.CLK(clk),
.GCLK(net9895)
);

ICGx2_ASAP7_75t_R merge9852(
.ENA(net392),
.SE(net2155),
.CLK(clk),
.GCLK(net9896)
);

ICGx2p67DC_ASAP7_75t_R merge9853(
.ENA(net2665),
.SE(net6407),
.CLK(clk),
.GCLK(net9897)
);

ICGx3_ASAP7_75t_R merge9854(
.ENA(net2560),
.SE(net2556),
.CLK(clk),
.GCLK(net9898)
);

ICGx4DC_ASAP7_75t_R merge9855(
.ENA(net3658),
.SE(net4204),
.CLK(clk),
.GCLK(net9899)
);

ICGx4_ASAP7_75t_R merge9856(
.ENA(net4018),
.SE(net4097),
.CLK(clk),
.GCLK(net9900)
);

ICGx5_ASAP7_75t_R merge9857(
.ENA(net6425),
.SE(net5345),
.CLK(clk),
.GCLK(net9901)
);

ICGx5p33DC_ASAP7_75t_R merge9858(
.ENA(net7158),
.SE(net8903),
.CLK(clk),
.GCLK(net9902)
);

ICGx6p67DC_ASAP7_75t_R merge9859(
.ENA(net8867),
.SE(net8735),
.CLK(clk),
.GCLK(net9903)
);

ICGx8DC_ASAP7_75t_R merge9860(
.ENA(net9803),
.SE(net2042),
.CLK(clk),
.GCLK(net9904)
);

XOR2x1_ASAP7_75t_R merge9861(
.A(net6854),
.B(net6939),
.Y(net9905)
);

ICGx1_ASAP7_75t_R merge9862(
.ENA(net8135),
.SE(net9002),
.CLK(clk),
.GCLK(net9906)
);

ICGx2_ASAP7_75t_R merge9863(
.ENA(net3221),
.SE(net9327),
.CLK(clk),
.GCLK(net9907)
);

ICGx2p67DC_ASAP7_75t_R merge9864(
.ENA(net8475),
.SE(net7531),
.CLK(clk),
.GCLK(net9908)
);

ICGx3_ASAP7_75t_R merge9865(
.ENA(net4830),
.SE(net4847),
.CLK(clk),
.GCLK(net9909)
);

ICGx4DC_ASAP7_75t_R merge9866(
.ENA(net4395),
.SE(net5075),
.CLK(clk),
.GCLK(net9910)
);

ICGx4_ASAP7_75t_R merge9867(
.ENA(net5510),
.SE(net4387),
.CLK(clk),
.GCLK(net9911)
);

ICGx5_ASAP7_75t_R merge9868(
.ENA(net8572),
.SE(net8623),
.CLK(clk),
.GCLK(net9912)
);

ICGx5p33DC_ASAP7_75t_R merge9869(
.ENA(net5067),
.SE(net8674),
.CLK(clk),
.GCLK(net9913)
);

ICGx6p67DC_ASAP7_75t_R merge9870(
.ENA(net6103),
.SE(net7197),
.CLK(clk),
.GCLK(net9914)
);

ICGx8DC_ASAP7_75t_R merge9871(
.ENA(net8747),
.SE(net8709),
.CLK(clk),
.GCLK(net9915)
);

ICGx1_ASAP7_75t_R merge9872(
.ENA(net4509),
.SE(net6022),
.CLK(clk),
.GCLK(net9916)
);

ICGx2_ASAP7_75t_R merge9873(
.ENA(net3321),
.SE(net3314),
.CLK(clk),
.GCLK(net9917)
);

ICGx2p67DC_ASAP7_75t_R merge9874(
.ENA(net6179),
.SE(net6088),
.CLK(clk),
.GCLK(net9918)
);

ICGx3_ASAP7_75t_R merge9875(
.ENA(net8998),
.SE(net8928),
.CLK(clk),
.GCLK(net9919)
);

ICGx4DC_ASAP7_75t_R merge9876(
.ENA(net2721),
.SE(net1746),
.CLK(clk),
.GCLK(net9920)
);

ICGx4_ASAP7_75t_R merge9877(
.ENA(net7294),
.SE(net6448),
.CLK(clk),
.GCLK(net9921)
);

ICGx5_ASAP7_75t_R merge9878(
.ENA(net7292),
.SE(net9043),
.CLK(clk),
.GCLK(out15)
);

ICGx5p33DC_ASAP7_75t_R merge9879(
.ENA(net1811),
.SE(net3675),
.CLK(clk),
.GCLK(net9922)
);

XOR2x2_ASAP7_75t_R merge9880(
.A(net6279),
.B(net5447),
.Y(net9923)
);

ICGx6p67DC_ASAP7_75t_R merge9881(
.ENA(net9010),
.SE(net7359),
.CLK(clk),
.GCLK(net9924)
);

ICGx8DC_ASAP7_75t_R merge9882(
.ENA(net8131),
.SE(net9013),
.CLK(clk),
.GCLK(net9925)
);

ICGx1_ASAP7_75t_R merge9883(
.ENA(net9532),
.SE(net9622),
.CLK(clk),
.GCLK(net9926)
);

ICGx2_ASAP7_75t_R merge9884(
.ENA(net9749),
.SE(net9716),
.CLK(clk),
.GCLK(net9927)
);

ICGx2p67DC_ASAP7_75t_R merge9885(
.ENA(net8836),
.SE(net7896),
.CLK(clk),
.GCLK(net9928)
);

ICGx3_ASAP7_75t_R merge9886(
.ENA(net8562),
.SE(net5672),
.CLK(clk),
.GCLK(net9929)
);

ICGx4DC_ASAP7_75t_R merge9887(
.ENA(net5685),
.SE(net9462),
.CLK(clk),
.GCLK(net9930)
);

XOR2xp5_ASAP7_75t_R merge9888(
.A(net4350),
.B(net5061),
.Y(net9931)
);

ICGx4_ASAP7_75t_R merge9889(
.ENA(net6766),
.SE(net6938),
.CLK(clk),
.GCLK(net9932)
);

ICGx5_ASAP7_75t_R merge9890(
.ENA(net9574),
.SE(net460),
.CLK(clk),
.GCLK(net9933)
);

ICGx5p33DC_ASAP7_75t_R merge9891(
.ENA(net628),
.SE(net9556),
.CLK(clk),
.GCLK(net9934)
);

ICGx6p67DC_ASAP7_75t_R merge9892(
.ENA(net9515),
.SE(net9771),
.CLK(clk),
.GCLK(net9935)
);

ICGx8DC_ASAP7_75t_R merge9893(
.ENA(net6060),
.SE(net5947),
.CLK(clk),
.GCLK(net9936)
);

ICGx1_ASAP7_75t_R merge9894(
.ENA(net4569),
.SE(net4564),
.CLK(clk),
.GCLK(net9937)
);

ICGx2_ASAP7_75t_R merge9895(
.ENA(net8563),
.SE(net8519),
.CLK(clk),
.GCLK(net9938)
);

ICGx2p67DC_ASAP7_75t_R merge9896(
.ENA(net7782),
.SE(net7913),
.CLK(clk),
.GCLK(net9939)
);

AND2x2_ASAP7_75t_R merge9897(
.A(net8670),
.B(net8736),
.Y(net9940)
);

ICGx3_ASAP7_75t_R merge9898(
.ENA(net9330),
.SE(net3508),
.CLK(clk),
.GCLK(net9941)
);

ICGx4DC_ASAP7_75t_R merge9899(
.ENA(net8599),
.SE(net8660),
.CLK(clk),
.GCLK(net9942)
);

ICGx4_ASAP7_75t_R merge9900(
.ENA(net6430),
.SE(net5517),
.CLK(clk),
.GCLK(net9943)
);

AND2x4_ASAP7_75t_R merge9901(
.A(net8901),
.B(net8987),
.Y(net9944)
);

ICGx5_ASAP7_75t_R merge9902(
.ENA(net4327),
.SE(net4518),
.CLK(clk),
.GCLK(net9945)
);

ICGx5p33DC_ASAP7_75t_R merge9903(
.ENA(net9839),
.SE(net9739),
.CLK(clk),
.GCLK(net9946)
);

ICGx6p67DC_ASAP7_75t_R merge9904(
.ENA(net8530),
.SE(net8590),
.CLK(clk),
.GCLK(net9947)
);

ICGx8DC_ASAP7_75t_R merge9905(
.ENA(net545),
.SE(net9394),
.CLK(clk),
.GCLK(net9948)
);

ICGx1_ASAP7_75t_R merge9906(
.ENA(net6339),
.SE(net5439),
.CLK(clk),
.GCLK(net9949)
);

ICGx2_ASAP7_75t_R merge9907(
.ENA(net9324),
.SE(net9674),
.CLK(clk),
.GCLK(net9950)
);

ICGx2p67DC_ASAP7_75t_R merge9908(
.ENA(net6602),
.SE(net9354),
.CLK(clk),
.GCLK(net9951)
);

ICGx3_ASAP7_75t_R merge9909(
.ENA(net9403),
.SE(net9521),
.CLK(clk),
.GCLK(net9952)
);

ICGx4DC_ASAP7_75t_R merge9910(
.ENA(net9628),
.SE(net278),
.CLK(clk),
.GCLK(net9953)
);

ICGx4_ASAP7_75t_R merge9911(
.ENA(net9598),
.SE(net9479),
.CLK(clk),
.GCLK(net9954)
);

ICGx5_ASAP7_75t_R merge9912(
.ENA(net9545),
.SE(net9092),
.CLK(clk),
.GCLK(net9955)
);

ICGx5p33DC_ASAP7_75t_R merge9913(
.ENA(net9878),
.SE(net1482),
.CLK(clk),
.GCLK(net9956)
);

ICGx6p67DC_ASAP7_75t_R merge9914(
.ENA(net9408),
.SE(net9792),
.CLK(clk),
.GCLK(net9957)
);

AND2x6_ASAP7_75t_R merge9915(
.A(net6274),
.B(net6175),
.Y(net9958)
);

ICGx8DC_ASAP7_75t_R merge9916(
.ENA(net8029),
.SE(net8797),
.CLK(clk),
.GCLK(net9959)
);

ICGx1_ASAP7_75t_R merge9917(
.ENA(net6438),
.SE(net8913),
.CLK(clk),
.GCLK(net9960)
);

ICGx2_ASAP7_75t_R merge9918(
.ENA(net9558),
.SE(net9740),
.CLK(clk),
.GCLK(net9961)
);

ICGx2p67DC_ASAP7_75t_R merge9919(
.ENA(net4554),
.SE(net4533),
.CLK(clk),
.GCLK(net9962)
);

ICGx3_ASAP7_75t_R merge9920(
.ENA(net9293),
.SE(net9610),
.CLK(clk),
.GCLK(net9963)
);

ICGx4DC_ASAP7_75t_R merge9921(
.ENA(net1416),
.SE(net9751),
.CLK(clk),
.GCLK(net9964)
);

ICGx4_ASAP7_75t_R merge9922(
.ENA(net8470),
.SE(net8602),
.CLK(clk),
.GCLK(net9965)
);

ICGx5_ASAP7_75t_R merge9923(
.ENA(net9522),
.SE(net9326),
.CLK(clk),
.GCLK(net9966)
);

ICGx5p33DC_ASAP7_75t_R merge9924(
.ENA(net6152),
.SE(net9262),
.CLK(clk),
.GCLK(net9967)
);

ICGx6p67DC_ASAP7_75t_R merge9925(
.ENA(net8215),
.SE(net8157),
.CLK(clk),
.GCLK(net9968)
);

ICGx8DC_ASAP7_75t_R merge9926(
.ENA(net9135),
.SE(net9471),
.CLK(clk),
.GCLK(net9969)
);

ICGx1_ASAP7_75t_R merge9927(
.ENA(net9570),
.SE(net2462),
.CLK(clk),
.GCLK(net9970)
);

ICGx2_ASAP7_75t_R merge9928(
.ENA(net6371),
.SE(net6363),
.CLK(clk),
.GCLK(net9971)
);

ICGx2p67DC_ASAP7_75t_R merge9929(
.ENA(net7121),
.SE(net7031),
.CLK(clk),
.GCLK(net9972)
);

ICGx3_ASAP7_75t_R merge9930(
.ENA(net9723),
.SE(net9529),
.CLK(clk),
.GCLK(net9973)
);

ICGx4DC_ASAP7_75t_R merge9931(
.ENA(net8746),
.SE(net8713),
.CLK(clk),
.GCLK(net9974)
);

ICGx4_ASAP7_75t_R merge9932(
.ENA(net8578),
.SE(net8405),
.CLK(clk),
.GCLK(net9975)
);

ICGx5_ASAP7_75t_R merge9933(
.ENA(net6447),
.SE(net9080),
.CLK(clk),
.GCLK(net9976)
);

ICGx5p33DC_ASAP7_75t_R merge9934(
.ENA(net9765),
.SE(net5854),
.CLK(clk),
.GCLK(net9977)
);

ICGx6p67DC_ASAP7_75t_R merge9935(
.ENA(net4747),
.SE(net3842),
.CLK(clk),
.GCLK(net9978)
);

ICGx8DC_ASAP7_75t_R merge9936(
.ENA(net7695),
.SE(net7697),
.CLK(clk),
.GCLK(net9979)
);

ICGx1_ASAP7_75t_R merge9937(
.ENA(net9437),
.SE(net9446),
.CLK(clk),
.GCLK(net9980)
);

HAxp5_ASAP7_75t_R merge9938(
.A(net7584),
.B(net8441),
.CON(net9981)
);

ICGx2_ASAP7_75t_R merge9939(
.ENA(net2200),
.SE(net9485),
.CLK(clk),
.GCLK(net9982)
);

ICGx2p67DC_ASAP7_75t_R merge9940(
.ENA(net7324),
.SE(net8060),
.CLK(clk),
.GCLK(net9983)
);

ICGx3_ASAP7_75t_R merge9941(
.ENA(net779),
.SE(net2664),
.CLK(clk),
.GCLK(net9984)
);

ICGx4DC_ASAP7_75t_R merge9942(
.ENA(net1397),
.SE(net9421),
.CLK(clk),
.GCLK(net9985)
);

ICGx4_ASAP7_75t_R merge9943(
.ENA(net3454),
.SE(net9691),
.CLK(clk),
.GCLK(net9986)
);

ICGx5_ASAP7_75t_R merge9944(
.ENA(net6355),
.SE(net1553),
.CLK(clk),
.GCLK(net9987)
);

ICGx5p33DC_ASAP7_75t_R merge9945(
.ENA(net8763),
.SE(net7310),
.CLK(clk),
.GCLK(net9988)
);

ICGx6p67DC_ASAP7_75t_R merge9946(
.ENA(net8638),
.SE(net7925),
.CLK(clk),
.GCLK(net9989)
);

ICGx8DC_ASAP7_75t_R merge9947(
.ENA(net9016),
.SE(net8825),
.CLK(clk),
.GCLK(net9990)
);

ICGx1_ASAP7_75t_R merge9948(
.ENA(net8720),
.SE(net8544),
.CLK(clk),
.GCLK(net9991)
);

ICGx2_ASAP7_75t_R merge9949(
.ENA(net9486),
.SE(net9728),
.CLK(clk),
.GCLK(net9992)
);

ICGx2p67DC_ASAP7_75t_R merge9950(
.ENA(net9601),
.SE(net1181),
.CLK(clk),
.GCLK(net9993)
);

ICGx3_ASAP7_75t_R merge9951(
.ENA(net9361),
.SE(net9123),
.CLK(clk),
.GCLK(net9994)
);

ICGx4DC_ASAP7_75t_R merge9952(
.ENA(net9006),
.SE(net8937),
.CLK(clk),
.GCLK(net9995)
);

ICGx4_ASAP7_75t_R merge9953(
.ENA(net6406),
.SE(net6435),
.CLK(clk),
.GCLK(out5)
);

ICGx5_ASAP7_75t_R merge9954(
.ENA(net9755),
.SE(net9784),
.CLK(clk),
.GCLK(net9996)
);

ICGx5p33DC_ASAP7_75t_R merge9955(
.ENA(net8200),
.SE(net8826),
.CLK(clk),
.GCLK(net9997)
);

ICGx6p67DC_ASAP7_75t_R merge9956(
.ENA(net9001),
.SE(net8948),
.CLK(clk),
.GCLK(net9998)
);

ICGx8DC_ASAP7_75t_R merge9957(
.ENA(net7288),
.SE(net7264),
.CLK(clk),
.GCLK(net9999)
);

NAND2x1_ASAP7_75t_R merge9958(
.A(net8860),
.B(net8789),
.Y(net10000)
);

ICGx1_ASAP7_75t_R merge9959(
.ENA(net8759),
.SE(net8105),
.CLK(clk),
.GCLK(net10001)
);

ICGx2_ASAP7_75t_R merge9960(
.ENA(net3471),
.SE(net2533),
.CLK(clk),
.GCLK(net10002)
);

ICGx2p67DC_ASAP7_75t_R merge9961(
.ENA(net9311),
.SE(net9589),
.CLK(clk),
.GCLK(net10003)
);

ICGx3_ASAP7_75t_R merge9962(
.ENA(net8091),
.SE(net8908),
.CLK(clk),
.GCLK(net10004)
);

ICGx4DC_ASAP7_75t_R merge9963(
.ENA(net8226),
.SE(net7345),
.CLK(clk),
.GCLK(net10005)
);

ICGx4_ASAP7_75t_R merge9964(
.ENA(net1220),
.SE(net9337),
.CLK(clk),
.GCLK(net10006)
);

NAND2x1p5_ASAP7_75t_R merge9965(
.A(net8627),
.B(net8654),
.Y(net10007)
);

ICGx5_ASAP7_75t_R merge9966(
.ENA(net8223),
.SE(net7336),
.CLK(clk),
.GCLK(net10008)
);

ICGx5p33DC_ASAP7_75t_R merge9967(
.ENA(net8634),
.SE(net8469),
.CLK(clk),
.GCLK(net10009)
);

ICGx6p67DC_ASAP7_75t_R merge9968(
.ENA(net7364),
.SE(net7308),
.CLK(clk),
.GCLK(net10010)
);

ICGx8DC_ASAP7_75t_R merge9969(
.ENA(net7368),
.SE(net7905),
.CLK(clk),
.GCLK(net10011)
);

ICGx1_ASAP7_75t_R merge9970(
.ENA(net424),
.SE(net3122),
.CLK(clk),
.GCLK(net10012)
);

ICGx2_ASAP7_75t_R merge9971(
.ENA(net9846),
.SE(net9432),
.CLK(clk),
.GCLK(net10013)
);

ICGx2p67DC_ASAP7_75t_R merge9972(
.ENA(net8467),
.SE(net8625),
.CLK(clk),
.GCLK(net10014)
);

ICGx3_ASAP7_75t_R merge9973(
.ENA(net9518),
.SE(net3468),
.CLK(clk),
.GCLK(net10015)
);

ICGx4DC_ASAP7_75t_R merge9974(
.ENA(net3900),
.SE(net9724),
.CLK(clk),
.GCLK(net10016)
);

ICGx4_ASAP7_75t_R merge9975(
.ENA(net9182),
.SE(net637),
.CLK(clk),
.GCLK(net10017)
);

ICGx5_ASAP7_75t_R merge9976(
.ENA(net7871),
.SE(net8886),
.CLK(clk),
.GCLK(net10018)
);

ICGx5p33DC_ASAP7_75t_R merge9977(
.ENA(net3971),
.SE(net9289),
.CLK(clk),
.GCLK(net10019)
);

ICGx6p67DC_ASAP7_75t_R merge9978(
.ENA(net5852),
.SE(net9473),
.CLK(clk),
.GCLK(net10020)
);

ICGx8DC_ASAP7_75t_R merge9979(
.ENA(net8061),
.SE(net8087),
.CLK(clk),
.GCLK(net10021)
);

ICGx1_ASAP7_75t_R merge9980(
.ENA(net9824),
.SE(net9606),
.CLK(clk),
.GCLK(net10022)
);

ICGx2_ASAP7_75t_R merge9981(
.ENA(net9695),
.SE(net5851),
.CLK(clk),
.GCLK(net10023)
);

ICGx2p67DC_ASAP7_75t_R merge9982(
.ENA(net9468),
.SE(net9544),
.CLK(clk),
.GCLK(net10024)
);

ICGx3_ASAP7_75t_R merge9983(
.ENA(net8900),
.SE(net8743),
.CLK(clk),
.GCLK(net10025)
);

ICGx4DC_ASAP7_75t_R merge9984(
.ENA(net8721),
.SE(net8703),
.CLK(clk),
.GCLK(net10026)
);

ICGx4_ASAP7_75t_R merge9985(
.ENA(net7367),
.SE(net7335),
.CLK(clk),
.GCLK(net10027)
);

ICGx5_ASAP7_75t_R merge9986(
.ENA(net9850),
.SE(net3060),
.CLK(clk),
.GCLK(net10028)
);

ICGx5p33DC_ASAP7_75t_R merge9987(
.ENA(net8856),
.SE(net8100),
.CLK(clk),
.GCLK(net10029)
);

ICGx6p67DC_ASAP7_75t_R merge9988(
.ENA(net7225),
.SE(net7256),
.CLK(clk),
.GCLK(net10030)
);

ICGx8DC_ASAP7_75t_R merge9989(
.ENA(net9168),
.SE(net9498),
.CLK(clk),
.GCLK(net10031)
);

ICGx1_ASAP7_75t_R merge9990(
.ENA(net8812),
.SE(net9694),
.CLK(clk),
.GCLK(net10032)
);

ICGx2_ASAP7_75t_R merge9991(
.ENA(net8149),
.SE(net8991),
.CLK(clk),
.GCLK(net10033)
);

ICGx2p67DC_ASAP7_75t_R merge9992(
.ENA(net9653),
.SE(net2548),
.CLK(clk),
.GCLK(net10034)
);

ICGx3_ASAP7_75t_R merge9993(
.ENA(net9138),
.SE(net9438),
.CLK(clk),
.GCLK(net10035)
);

ICGx4DC_ASAP7_75t_R merge9994(
.ENA(net9703),
.SE(net9591),
.CLK(clk),
.GCLK(net10036)
);

ICGx4_ASAP7_75t_R merge9995(
.ENA(net9028),
.SE(net8994),
.CLK(clk),
.GCLK(net10037)
);

ICGx5_ASAP7_75t_R merge9996(
.ENA(net9511),
.SE(net4024),
.CLK(clk),
.GCLK(net10038)
);

ICGx5p33DC_ASAP7_75t_R merge9997(
.ENA(net9374),
.SE(net9444),
.CLK(clk),
.GCLK(net10039)
);

NAND2x2_ASAP7_75t_R merge9998(
.A(net8931),
.B(net8052),
.Y(net10040)
);

ICGx6p67DC_ASAP7_75t_R merge9999(
.ENA(net7259),
.SE(net7343),
.CLK(clk),
.GCLK(net10041)
);

ICGx8DC_ASAP7_75t_R merge10000(
.ENA(net9380),
.SE(net9260),
.CLK(clk),
.GCLK(net10042)
);

ICGx1_ASAP7_75t_R merge10001(
.ENA(net7357),
.SE(net8988),
.CLK(clk),
.GCLK(net10043)
);

ICGx2_ASAP7_75t_R merge10002(
.ENA(net4420),
.SE(net5337),
.CLK(clk),
.GCLK(net10044)
);

ICGx2p67DC_ASAP7_75t_R merge10003(
.ENA(net9635),
.SE(net9458),
.CLK(clk),
.GCLK(net10045)
);

ICGx3_ASAP7_75t_R merge10004(
.ENA(net8138),
.SE(net9000),
.CLK(clk),
.GCLK(net10046)
);

ICGx4DC_ASAP7_75t_R merge10005(
.ENA(net2046),
.SE(net225),
.CLK(clk),
.GCLK(net10047)
);

ICGx4_ASAP7_75t_R merge10006(
.ENA(net8037),
.SE(net9809),
.CLK(clk),
.GCLK(net10048)
);

ICGx5_ASAP7_75t_R merge10007(
.ENA(net9673),
.SE(net7361),
.CLK(clk),
.GCLK(net10049)
);

ICGx5p33DC_ASAP7_75t_R merge10008(
.ENA(net8432),
.SE(net7587),
.CLK(clk),
.GCLK(net10050)
);

ICGx6p67DC_ASAP7_75t_R merge10009(
.ENA(net3154),
.SE(net1310),
.CLK(clk),
.GCLK(net10051)
);

ICGx8DC_ASAP7_75t_R merge10010(
.ENA(net6640),
.SE(net7591),
.CLK(clk),
.GCLK(net10052)
);

ICGx1_ASAP7_75t_R merge10011(
.ENA(net9159),
.SE(net9129),
.CLK(clk),
.GCLK(net10053)
);

ICGx2_ASAP7_75t_R merge10012(
.ENA(net9581),
.SE(net9874),
.CLK(clk),
.GCLK(net10054)
);

ICGx2p67DC_ASAP7_75t_R merge10013(
.ENA(net8932),
.SE(net8095),
.CLK(clk),
.GCLK(net10055)
);

ICGx3_ASAP7_75t_R merge10014(
.ENA(net9166),
.SE(net9506),
.CLK(clk),
.GCLK(net10056)
);

ICGx4DC_ASAP7_75t_R merge10015(
.ENA(net8874),
.SE(net8916),
.CLK(clk),
.GCLK(net10057)
);

ICGx4_ASAP7_75t_R merge10016(
.ENA(net9004),
.SE(net8201),
.CLK(clk),
.GCLK(net10058)
);

ICGx5_ASAP7_75t_R merge10017(
.ENA(net7795),
.SE(net9820),
.CLK(clk),
.GCLK(net10059)
);

ICGx5p33DC_ASAP7_75t_R merge10018(
.ENA(net7351),
.SE(net9020),
.CLK(clk),
.GCLK(net10060)
);

ICGx6p67DC_ASAP7_75t_R merge10019(
.ENA(net8153),
.SE(net9240),
.CLK(clk),
.GCLK(net10061)
);

ICGx8DC_ASAP7_75t_R merge10020(
.ENA(net3502),
.SE(net9668),
.CLK(clk),
.GCLK(net10062)
);

ICGx1_ASAP7_75t_R merge10021(
.ENA(net9541),
.SE(net9732),
.CLK(clk),
.GCLK(net10063)
);

ICGx2_ASAP7_75t_R merge10022(
.ENA(net9538),
.SE(net2040),
.CLK(clk),
.GCLK(net10064)
);

ICGx2p67DC_ASAP7_75t_R merge10023(
.ENA(net8213),
.SE(net8218),
.CLK(clk),
.GCLK(out23)
);

ICGx3_ASAP7_75t_R merge10024(
.ENA(net1325),
.SE(net3185),
.CLK(clk),
.GCLK(net10065)
);

ICGx4DC_ASAP7_75t_R merge10025(
.ENA(net9397),
.SE(net9459),
.CLK(clk),
.GCLK(net10066)
);

ICGx4_ASAP7_75t_R merge10026(
.ENA(net9829),
.SE(net9853),
.CLK(clk),
.GCLK(net10067)
);

NAND2xp33_ASAP7_75t_R merge10027(
.A(net8956),
.B(net8979),
.Y(net10068)
);

ICGx5_ASAP7_75t_R merge10028(
.ENA(net8243),
.SE(net8220),
.CLK(clk),
.GCLK(net10069)
);

ICGx5p33DC_ASAP7_75t_R merge10029(
.ENA(net9460),
.SE(net5862),
.CLK(clk),
.GCLK(net10070)
);

ICGx6p67DC_ASAP7_75t_R merge10030(
.ENA(net9332),
.SE(net9617),
.CLK(clk),
.GCLK(net10071)
);

ICGx8DC_ASAP7_75t_R merge10031(
.ENA(net7355),
.SE(net7358),
.CLK(clk),
.GCLK(net10072)
);

ICGx1_ASAP7_75t_R merge10032(
.ENA(net9645),
.SE(net9633),
.CLK(clk),
.GCLK(net10073)
);

ICGx2_ASAP7_75t_R merge10033(
.ENA(net9049),
.SE(net8978),
.CLK(clk),
.GCLK(net10074)
);

ICGx2p67DC_ASAP7_75t_R merge10034(
.ENA(net8246),
.SE(net8224),
.CLK(clk),
.GCLK(net10075)
);

ICGx3_ASAP7_75t_R merge10035(
.ENA(net9405),
.SE(net9770),
.CLK(clk),
.GCLK(net10076)
);

NAND2xp5_ASAP7_75t_R merge10036(
.A(net9041),
.B(net8230),
.Y(net10077)
);

ICGx4DC_ASAP7_75t_R merge10037(
.ENA(net9643),
.SE(net9443),
.CLK(clk),
.GCLK(net10078)
);

ICGx4_ASAP7_75t_R merge10038(
.ENA(net9551),
.SE(net9329),
.CLK(clk),
.GCLK(net10079)
);

ICGx5_ASAP7_75t_R merge10039(
.ENA(net9721),
.SE(net9502),
.CLK(clk),
.GCLK(net10080)
);

ICGx5p33DC_ASAP7_75t_R merge10040(
.ENA(net8219),
.GCLK(net8225),
.CLK(clk)
);

ICGx6p67DC_ASAP7_75t_R merge10041(
.ENA(net9905),
.SE(net6867),
.CLK(clk),
.GCLK(net10081)
);

ICGx8DC_ASAP7_75t_R merge10042(
.ENA(net1470),
.SE(net9838),
.CLK(clk),
.GCLK(net10082)
);

ICGx1_ASAP7_75t_R merge10043(
.ENA(net9883),
.SE(net9116),
.CLK(clk),
.GCLK(net10083)
);

ICGx2_ASAP7_75t_R merge10044(
.ENA(net9734),
.SE(net4149),
.CLK(clk),
.GCLK(net10084)
);

ICGx2p67DC_ASAP7_75t_R merge10045(
.ENA(net9530),
.SE(net9873),
.CLK(clk),
.GCLK(net10085)
);

ICGx3_ASAP7_75t_R merge10046(
.ENA(net9042),
.SE(net9059),
.CLK(clk),
.GCLK(net10086)
);

ICGx4DC_ASAP7_75t_R merge10047(
.ENA(net9410),
.SE(net9616),
.CLK(clk),
.GCLK(net10087)
);

ICGx4_ASAP7_75t_R merge10048(
.ENA(net8228),
.SE(net8229),
.CLK(clk),
.GCLK(out10)
);

ICGx5_ASAP7_75t_R merge10049(
.ENA(net2111),
.SE(net9602),
.CLK(clk),
.GCLK(net10088)
);

ICGx5p33DC_ASAP7_75t_R merge10050(
.ENA(net4072),
.SE(net9793),
.CLK(clk),
.GCLK(net10089)
);

ICGx6p67DC_ASAP7_75t_R merge10051(
.ENA(net9074),
.SE(net9075),
.CLK(clk),
.GCLK(net10090)
);

ICGx8DC_ASAP7_75t_R merge10052(
.ENA(net9461),
.SE(net4889),
.CLK(clk),
.GCLK(net10091)
);

ICGx1_ASAP7_75t_R merge10053(
.ENA(net9081),
.SE(net8231),
.CLK(clk),
.GCLK(out7)
);

ICGx2_ASAP7_75t_R merge10054(
.ENA(net10007),
.SE(net9126),
.CLK(clk),
.GCLK(net10092)
);

ICGx2p67DC_ASAP7_75t_R merge10055(
.ENA(net9344),
.SE(net9254),
.CLK(clk),
.GCLK(net10093)
);

ICGx3_ASAP7_75t_R merge10056(
.ENA(net9370),
.SE(net9423),
.CLK(clk),
.GCLK(net10094)
);

ICGx4DC_ASAP7_75t_R merge10057(
.ENA(net9209),
.SE(net9768),
.CLK(clk),
.GCLK(net10095)
);

ICGx4_ASAP7_75t_R merge10058(
.ENA(net9470),
.SE(net2038),
.CLK(clk),
.GCLK(net10096)
);

ICGx5_ASAP7_75t_R merge10059(
.ENA(net9319),
.SE(net3588),
.CLK(clk),
.GCLK(net10097)
);

ICGx5p33DC_ASAP7_75t_R merge10060(
.ENA(net10040),
.SE(net6337),
.CLK(clk),
.GCLK(net10098)
);

ICGx6p67DC_ASAP7_75t_R merge10061(
.ENA(net9753),
.SE(net9816),
.CLK(clk),
.GCLK(net10099)
);

ICGx8DC_ASAP7_75t_R merge10062(
.ENA(net9481),
.SE(net9822),
.CLK(clk),
.GCLK(net10100)
);

ICGx1_ASAP7_75t_R merge10063(
.ENA(net9840),
.SE(net1409),
.CLK(clk),
.GCLK(net10101)
);

ICGx2_ASAP7_75t_R merge10064(
.ENA(net9372),
.SE(net2614),
.CLK(clk),
.GCLK(net10102)
);

ICGx2p67DC_ASAP7_75t_R merge10065(
.ENA(net9887),
.SE(net9392),
.CLK(clk),
.GCLK(net10103)
);

ICGx3_ASAP7_75t_R merge10066(
.ENA(net9626),
.SE(net6149),
.CLK(clk),
.GCLK(net10104)
);

ICGx4DC_ASAP7_75t_R merge10067(
.ENA(net9750),
.SE(net9701),
.CLK(clk),
.GCLK(net10105)
);

ICGx4_ASAP7_75t_R merge10068(
.ENA(net9124),
.SE(net2240),
.CLK(clk),
.GCLK(net10106)
);

ICGx5_ASAP7_75t_R merge10069(
.ENA(net9351),
.SE(net9797),
.CLK(clk),
.GCLK(net10107)
);

ICGx5p33DC_ASAP7_75t_R merge10070(
.ENA(net289),
.SE(net9796),
.CLK(clk),
.GCLK(net10108)
);

ICGx6p67DC_ASAP7_75t_R merge10071(
.ENA(net9255),
.SE(net9154),
.CLK(clk),
.GCLK(net10109)
);

ICGx8DC_ASAP7_75t_R merge10072(
.ENA(net6916),
.SE(net9605),
.CLK(clk),
.GCLK(net10110)
);

ICGx1_ASAP7_75t_R merge10073(
.ENA(net454),
.SE(net9426),
.CLK(clk),
.GCLK(net10111)
);

ICGx2_ASAP7_75t_R merge10074(
.ENA(net9680),
.SE(net9353),
.CLK(clk),
.GCLK(net10112)
);

ICGx2p67DC_ASAP7_75t_R merge10075(
.ENA(net4106),
.SE(net2053),
.CLK(clk),
.GCLK(net10113)
);

ICGx3_ASAP7_75t_R merge10076(
.ENA(net9206),
.SE(net9804),
.CLK(clk),
.GCLK(net10114)
);

ICGx4DC_ASAP7_75t_R merge10077(
.ENA(net9885),
.SE(net9343),
.CLK(clk),
.GCLK(net10115)
);

ICGx4_ASAP7_75t_R merge10078(
.ENA(net9236),
.SE(net9865),
.CLK(clk),
.GCLK(net10116)
);

ICGx5_ASAP7_75t_R merge10079(
.ENA(net9594),
.SE(net9621),
.CLK(clk),
.GCLK(net10117)
);

ICGx5p33DC_ASAP7_75t_R merge10080(
.ENA(net9296),
.SE(net9312),
.CLK(clk),
.GCLK(net10118)
);

ICGx6p67DC_ASAP7_75t_R merge10081(
.ENA(net9373),
.SE(net9313),
.CLK(clk),
.GCLK(net10119)
);

ICGx8DC_ASAP7_75t_R merge10082(
.ENA(net5011),
.SE(net9448),
.CLK(clk),
.GCLK(net10120)
);

ICGx1_ASAP7_75t_R merge10083(
.ENA(net9451),
.SE(net10077),
.CLK(clk),
.GCLK(net10121)
);

ICGx2_ASAP7_75t_R merge10084(
.ENA(net9362),
.SE(net7175),
.CLK(clk),
.GCLK(net10122)
);

ICGx2p67DC_ASAP7_75t_R merge10085(
.ENA(net9505),
.SE(net9866),
.CLK(clk),
.GCLK(net10123)
);

ICGx3_ASAP7_75t_R merge10086(
.ENA(net9931),
.SE(net9457),
.CLK(clk),
.GCLK(net10124)
);

ICGx4DC_ASAP7_75t_R merge10087(
.ENA(net9944),
.SE(net8883),
.CLK(clk),
.GCLK(net10125)
);

ICGx4_ASAP7_75t_R merge10088(
.ENA(net9781),
.SE(net9692),
.CLK(clk),
.GCLK(net10126)
);

ICGx5_ASAP7_75t_R merge10089(
.ENA(net6187),
.SE(net5930),
.CLK(clk),
.GCLK(net10127)
);

ICGx5p33DC_ASAP7_75t_R merge10090(
.ENA(net9503),
.SE(net9360),
.CLK(clk),
.GCLK(net10128)
);

ICGx6p67DC_ASAP7_75t_R merge10091(
.ENA(net9317),
.SE(net9101),
.CLK(clk),
.GCLK(net10129)
);

ICGx8DC_ASAP7_75t_R merge10092(
.ENA(net9156),
.SE(net4098),
.CLK(clk),
.GCLK(net10130)
);

ICGx1_ASAP7_75t_R merge10093(
.ENA(net9283),
.SE(net1434),
.CLK(clk),
.GCLK(net10131)
);

ICGx2_ASAP7_75t_R merge10094(
.ENA(net9534),
.SE(net9940),
.CLK(clk),
.GCLK(net10132)
);

ICGx2p67DC_ASAP7_75t_R merge10095(
.ENA(net9699),
.SE(net9321),
.CLK(clk),
.GCLK(net10133)
);

ICGx3_ASAP7_75t_R merge10096(
.ENA(net9767),
.SE(net9700),
.CLK(clk),
.GCLK(net10134)
);

ICGx4DC_ASAP7_75t_R merge10097(
.ENA(net9577),
.SE(net7039),
.CLK(clk),
.GCLK(net10135)
);

ICGx4_ASAP7_75t_R merge10098(
.ENA(net9385),
.SE(net9456),
.CLK(clk),
.GCLK(net10136)
);

ICGx5_ASAP7_75t_R merge10099(
.ENA(net9489),
.SE(net9492),
.CLK(clk),
.GCLK(net10137)
);

ICGx5p33DC_ASAP7_75t_R merge10100(
.ENA(net3909),
.SE(net9872),
.CLK(clk),
.GCLK(net10138)
);

ICGx6p67DC_ASAP7_75t_R merge10101(
.ENA(net9452),
.SE(net9799),
.CLK(clk),
.GCLK(net10139)
);

ICGx8DC_ASAP7_75t_R merge10102(
.ENA(net10000),
.SE(net8926),
.CLK(clk),
.GCLK(net10140)
);

ICGx1_ASAP7_75t_R merge10103(
.ENA(net9098),
.SE(net9879),
.CLK(clk),
.GCLK(net10141)
);

ICGx2_ASAP7_75t_R merge10104(
.ENA(net9367),
.SE(net9718),
.CLK(clk),
.GCLK(net10142)
);

ICGx2p67DC_ASAP7_75t_R merge10105(
.ENA(net9646),
.SE(net7903),
.CLK(clk),
.GCLK(net10143)
);

ICGx3_ASAP7_75t_R merge10106(
.ENA(net7864),
.SE(net9833),
.CLK(clk),
.GCLK(net10144)
);

ICGx4DC_ASAP7_75t_R merge10107(
.ENA(net5855),
.SE(net9676),
.CLK(clk),
.GCLK(net10145)
);

ICGx4_ASAP7_75t_R merge10108(
.ENA(net9837),
.SE(net9848),
.CLK(clk),
.GCLK(net10146)
);

ICGx5_ASAP7_75t_R merge10109(
.ENA(net9880),
.SE(net9808),
.CLK(clk),
.GCLK(net10147)
);

ICGx5p33DC_ASAP7_75t_R merge10110(
.ENA(net9549),
.SE(net9415),
.CLK(clk),
.GCLK(net10148)
);

ICGx6p67DC_ASAP7_75t_R merge10111(
.ENA(net9715),
.SE(net9655),
.CLK(clk),
.GCLK(net10149)
);

ICGx8DC_ASAP7_75t_R merge10112(
.ENA(net9119),
.SE(net9146),
.CLK(clk),
.GCLK(net10150)
);

ICGx1_ASAP7_75t_R merge10113(
.ENA(net9891),
.SE(net9798),
.CLK(clk),
.GCLK(net10151)
);

ICGx2_ASAP7_75t_R merge10114(
.ENA(net9669),
.SE(net9268),
.CLK(clk),
.GCLK(net10152)
);

ICGx2p67DC_ASAP7_75t_R merge10115(
.ENA(net9810),
.SE(net9958),
.CLK(clk),
.GCLK(net10153)
);

ICGx3_ASAP7_75t_R merge10116(
.ENA(net7869),
.SE(net9175),
.CLK(clk),
.GCLK(net10154)
);

ICGx4DC_ASAP7_75t_R merge10117(
.ENA(net9141),
.SE(net9198),
.CLK(clk),
.GCLK(net10155)
);

ICGx4_ASAP7_75t_R merge10118(
.ENA(net9366),
.SE(net9664),
.CLK(clk),
.GCLK(net10156)
);

ICGx5_ASAP7_75t_R merge10119(
.ENA(net9584),
.SE(net9535),
.CLK(clk),
.GCLK(net10157)
);

ICGx5p33DC_ASAP7_75t_R merge10120(
.ENA(net9180),
.SE(net6771),
.CLK(clk),
.GCLK(net10158)
);

ICGx6p67DC_ASAP7_75t_R merge10121(
.ENA(net9323),
.SE(net10068),
.CLK(clk),
.GCLK(net10159)
);

ICGx8DC_ASAP7_75t_R merge10122(
.ENA(net3568),
.SE(net9442),
.CLK(clk),
.GCLK(net10160)
);

ICGx1_ASAP7_75t_R merge10123(
.ENA(net2152),
.SE(net9890),
.CLK(clk),
.GCLK(net10161)
);

ICGx2_ASAP7_75t_R merge10124(
.ENA(net9923),
.SE(net9542),
.CLK(clk),
.GCLK(out0)
);

ICGx2p67DC_ASAP7_75t_R merge10125(
.ENA(net9318),
.SE(net2576),
.CLK(clk),
.GCLK(net10162)
);

ICGx3_ASAP7_75t_R merge10126(
.ENA(net9619),
.SE(net9466),
.CLK(clk),
.GCLK(net10163)
);

ICGx4DC_ASAP7_75t_R merge10127(
.ENA(net9183),
.SE(net9714),
.CLK(clk),
.GCLK(net10164)
);

ICGx4_ASAP7_75t_R merge10128(
.ENA(net9571),
.SE(net9742),
.CLK(clk),
.GCLK(net10165)
);

ICGx5_ASAP7_75t_R merge10129(
.ENA(net9365),
.SE(net9834),
.CLK(clk),
.GCLK(net10166)
);

ICGx5p33DC_ASAP7_75t_R merge10130(
.ENA(net9780),
.SE(net7027),
.CLK(clk),
.GCLK(net10167)
);

ICGx6p67DC_ASAP7_75t_R merge10131(
.ENA(net5007),
.SE(net9407),
.CLK(clk),
.GCLK(net10168)
);

ICGx8DC_ASAP7_75t_R merge10132(
.ENA(net4430),
.SE(net9433),
.CLK(clk),
.GCLK(net10169)
);

ICGx1_ASAP7_75t_R merge10133(
.ENA(net9111),
.SE(net9376),
.CLK(clk),
.GCLK(net10170)
);

ICGx2_ASAP7_75t_R merge10134(
.ENA(net9861),
.SE(net9981),
.CLK(clk),
.GCLK(net10171)
);

ICGx2p67DC_ASAP7_75t_R merge10135(
.ENA(net6276),
.SE(net9540),
.CLK(clk),
.GCLK(net10172)
);

DFFHQNx1_ASAP7_75t_R s10136(
.D(net136),
.CLK(clk),
.QN(net10173)
);

DFFHQNx2_ASAP7_75t_R s10137(
.D(net139),
.CLK(clk),
.QN(net10174)
);

DFFHQNx3_ASAP7_75t_R s10138(
.D(net217),
.CLK(clk),
.QN(net10175)
);

DFFHQx4_ASAP7_75t_R s10139(
.D(net301),
.CLK(clk),
.Q(net10176)
);

DFFLQNx1_ASAP7_75t_R s10140(
.D(net309),
.CLK(clk),
.QN(net10177)
);

DFFLQNx2_ASAP7_75t_R s10141(
.D(net391),
.CLK(clk),
.QN(net10178)
);

DFFLQNx3_ASAP7_75t_R s10142(
.D(net473),
.CLK(clk),
.QN(net10179)
);

DFFLQx4_ASAP7_75t_R s10143(
.D(net539),
.CLK(clk),
.Q(net10180)
);

DHLx1_ASAP7_75t_R s10144(
.D(net542),
.CLK(clk),
.Q(net10181)
);

DHLx2_ASAP7_75t_R s10145(
.D(net562),
.CLK(clk),
.Q(net10182)
);

DHLx3_ASAP7_75t_R s10146(
.D(net563),
.CLK(clk),
.Q(net10183)
);

DLLx1_ASAP7_75t_R s10147(
.D(net712),
.CLK(clk),
.Q(net10184)
);

DLLx2_ASAP7_75t_R s10148(
.D(net815),
.CLK(clk),
.Q(net10185)
);

DLLx3_ASAP7_75t_R s10149(
.D(net1009),
.CLK(clk),
.Q(net10186)
);

DFFHQNx1_ASAP7_75t_R s10150(
.D(net1062),
.CLK(clk),
.QN(net10187)
);

DFFHQNx2_ASAP7_75t_R s10151(
.D(net1065),
.CLK(clk),
.QN(net10188)
);

DFFHQNx3_ASAP7_75t_R s10152(
.D(net1066),
.CLK(clk),
.QN(net10189)
);

DFFHQx4_ASAP7_75t_R s10153(
.D(net1151),
.CLK(clk),
.Q(net10190)
);

DFFLQNx1_ASAP7_75t_R s10154(
.D(net1271),
.CLK(clk),
.QN(net10191)
);

DFFLQNx2_ASAP7_75t_R s10155(
.D(net1300),
.CLK(clk),
.QN(net10192)
);

DFFLQNx3_ASAP7_75t_R s10156(
.D(net1375),
.CLK(clk),
.QN(net10193)
);

DFFLQx4_ASAP7_75t_R s10157(
.D(net1396),
.CLK(clk),
.Q(net10194)
);

DHLx1_ASAP7_75t_R s10158(
.D(net1399),
.CLK(clk),
.Q(net10195)
);

DHLx2_ASAP7_75t_R s10159(
.D(net1463),
.CLK(clk),
.Q(net10196)
);

DHLx3_ASAP7_75t_R s10160(
.D(net1555),
.CLK(clk),
.Q(net10197)
);

DLLx1_ASAP7_75t_R s10161(
.D(net1562),
.CLK(clk),
.Q(net10198)
);

DLLx2_ASAP7_75t_R s10162(
.D(net1563),
.CLK(clk),
.Q(net10199)
);

DLLx3_ASAP7_75t_R s10163(
.D(net1679),
.CLK(clk),
.Q(net10200)
);

DFFHQNx1_ASAP7_75t_R s10164(
.D(net1762),
.CLK(clk),
.QN(net10201)
);

DFFHQNx2_ASAP7_75t_R s10165(
.D(net1770),
.CLK(clk),
.QN(net10202)
);

DFFHQNx3_ASAP7_75t_R s10166(
.D(net1799),
.CLK(clk),
.QN(net10203)
);

DFFHQx4_ASAP7_75t_R s10167(
.D(net1906),
.CLK(clk),
.Q(net10204)
);

DFFLQNx1_ASAP7_75t_R s10168(
.D(net2047),
.CLK(clk),
.QN(net10205)
);

DFFLQNx2_ASAP7_75t_R s10169(
.D(net2213),
.CLK(clk),
.QN(net10206)
);

DFFLQNx3_ASAP7_75t_R s10170(
.D(net2215),
.CLK(clk),
.QN(net10207)
);

DFFLQx4_ASAP7_75t_R s10171(
.D(net2222),
.CLK(clk),
.Q(net10208)
);

DHLx1_ASAP7_75t_R s10172(
.D(net2322),
.CLK(clk),
.Q(net10209)
);

DHLx2_ASAP7_75t_R s10173(
.D(net2324),
.CLK(clk),
.Q(net10210)
);

DHLx3_ASAP7_75t_R s10174(
.D(net2326),
.CLK(clk),
.Q(net10211)
);

DLLx1_ASAP7_75t_R s10175(
.D(net2331),
.CLK(clk),
.Q(net10212)
);

DLLx2_ASAP7_75t_R s10176(
.D(net2406),
.CLK(clk),
.Q(net10213)
);

DLLx3_ASAP7_75t_R s10177(
.D(net2489),
.CLK(clk),
.Q(net10214)
);

DFFHQNx1_ASAP7_75t_R s10178(
.D(net2651),
.CLK(clk),
.QN(net10215)
);

DFFHQNx2_ASAP7_75t_R s10179(
.D(net2718),
.CLK(clk),
.QN(net10216)
);

DFFHQNx3_ASAP7_75t_R s10180(
.D(net2737),
.CLK(clk),
.QN(net10217)
);

DFFHQx4_ASAP7_75t_R s10181(
.D(net2753),
.CLK(clk),
.Q(net10218)
);

DFFLQNx1_ASAP7_75t_R s10182(
.D(net2835),
.CLK(clk),
.QN(net10219)
);

DFFLQNx2_ASAP7_75t_R s10183(
.D(net2895),
.CLK(clk),
.QN(net10220)
);

DFFLQNx3_ASAP7_75t_R s10184(
.D(net3050),
.CLK(clk),
.QN(net10221)
);

DFFLQx4_ASAP7_75t_R s10185(
.D(net3072),
.CLK(clk),
.Q(net10222)
);

DHLx1_ASAP7_75t_R s10186(
.D(net3081),
.CLK(clk),
.Q(net10223)
);

DHLx2_ASAP7_75t_R s10187(
.D(net3123),
.CLK(clk),
.Q(net10224)
);

DHLx3_ASAP7_75t_R s10188(
.D(net3308),
.CLK(clk),
.Q(net10225)
);

DLLx1_ASAP7_75t_R s10189(
.D(net3328),
.CLK(clk),
.Q(net10226)
);

DLLx2_ASAP7_75t_R s10190(
.D(net3488),
.CLK(clk),
.Q(net10227)
);

DLLx3_ASAP7_75t_R s10191(
.D(net3507),
.CLK(clk),
.Q(net10228)
);

DFFHQNx1_ASAP7_75t_R s10192(
.D(net3590),
.CLK(clk),
.QN(net10229)
);

DFFHQNx2_ASAP7_75t_R s10193(
.D(net3659),
.CLK(clk),
.QN(net10230)
);

DFFHQNx3_ASAP7_75t_R s10194(
.D(net3661),
.CLK(clk),
.QN(net10231)
);

DFFHQx4_ASAP7_75t_R s10195(
.D(net3665),
.CLK(clk),
.Q(net10232)
);

DFFLQNx1_ASAP7_75t_R s10196(
.D(net3668),
.CLK(clk),
.QN(net10233)
);

DFFLQNx2_ASAP7_75t_R s10197(
.D(net3671),
.CLK(clk),
.QN(net10234)
);

DFFLQNx3_ASAP7_75t_R s10198(
.D(net3737),
.CLK(clk),
.QN(net10235)
);

DFFLQx4_ASAP7_75t_R s10199(
.D(net3818),
.CLK(clk),
.Q(net10236)
);

DHLx1_ASAP7_75t_R s10200(
.D(net3823),
.CLK(clk),
.Q(net10237)
);

DHLx2_ASAP7_75t_R s10201(
.D(net3918),
.CLK(clk),
.Q(net10238)
);

DHLx3_ASAP7_75t_R s10202(
.D(net3953),
.CLK(clk),
.Q(net10239)
);

DLLx1_ASAP7_75t_R s10203(
.D(net4090),
.CLK(clk),
.Q(net10240)
);

DLLx2_ASAP7_75t_R s10204(
.D(net4100),
.CLK(clk),
.Q(net10241)
);

DLLx3_ASAP7_75t_R s10205(
.D(net4292),
.CLK(clk),
.Q(net10242)
);

DFFHQNx1_ASAP7_75t_R s10206(
.D(net4316),
.CLK(clk),
.QN(net10243)
);

DFFHQNx2_ASAP7_75t_R s10207(
.D(net4338),
.CLK(clk),
.QN(net10244)
);

DFFHQNx3_ASAP7_75t_R s10208(
.D(net4516),
.CLK(clk),
.QN(net10245)
);

DFFHQx4_ASAP7_75t_R s10209(
.D(net4559),
.CLK(clk),
.Q(net10246)
);

DFFLQNx1_ASAP7_75t_R s10210(
.D(net4570),
.CLK(clk),
.QN(net10247)
);

DFFLQNx2_ASAP7_75t_R s10211(
.D(net4582),
.CLK(clk),
.QN(net10248)
);

DFFLQNx3_ASAP7_75t_R s10212(
.D(net4675),
.CLK(clk),
.QN(net10249)
);

DFFLQx4_ASAP7_75t_R s10213(
.D(net4682),
.CLK(clk),
.Q(net10250)
);

DHLx1_ASAP7_75t_R s10214(
.D(net4683),
.CLK(clk),
.Q(net10251)
);

DHLx2_ASAP7_75t_R s10215(
.D(net4689),
.CLK(clk),
.Q(net10252)
);

DHLx3_ASAP7_75t_R s10216(
.D(net4772),
.CLK(clk),
.Q(net10253)
);

DLLx1_ASAP7_75t_R s10217(
.D(net4910),
.CLK(clk),
.Q(net10254)
);

DLLx2_ASAP7_75t_R s10218(
.D(net4997),
.CLK(clk),
.Q(net10255)
);

DLLx3_ASAP7_75t_R s10219(
.D(net5144),
.CLK(clk),
.Q(net10256)
);

DFFHQNx1_ASAP7_75t_R s10220(
.D(net5161),
.CLK(clk),
.QN(net10257)
);

DFFHQNx2_ASAP7_75t_R s10221(
.D(net5270),
.CLK(clk),
.QN(net10258)
);

DFFHQNx3_ASAP7_75t_R s10222(
.D(net5272),
.CLK(clk),
.QN(net10259)
);

DFFHQx4_ASAP7_75t_R s10223(
.D(net5434),
.CLK(clk),
.Q(net10260)
);

DFFLQNx1_ASAP7_75t_R s10224(
.D(net5451),
.CLK(clk),
.QN(net10261)
);

DFFLQNx2_ASAP7_75t_R s10225(
.D(net5524),
.CLK(clk),
.QN(net10262)
);

DFFLQNx3_ASAP7_75t_R s10226(
.D(net5601),
.CLK(clk),
.QN(net10263)
);

DFFLQx4_ASAP7_75t_R s10227(
.D(net5606),
.CLK(clk),
.Q(net10264)
);

DHLx1_ASAP7_75t_R s10228(
.D(net5611),
.CLK(clk),
.Q(net10265)
);

DHLx2_ASAP7_75t_R s10229(
.D(net5679),
.CLK(clk),
.Q(net10266)
);

DHLx3_ASAP7_75t_R s10230(
.D(net5694),
.CLK(clk),
.Q(net10267)
);

DLLx1_ASAP7_75t_R s10231(
.D(net5695),
.CLK(clk),
.Q(net10268)
);

DLLx2_ASAP7_75t_R s10232(
.D(net5781),
.CLK(clk),
.Q(net10269)
);

DLLx3_ASAP7_75t_R s10233(
.D(net5946),
.CLK(clk),
.Q(net10270)
);

DFFHQNx1_ASAP7_75t_R s10234(
.D(net6092),
.CLK(clk),
.QN(net10271)
);

DFFHQNx2_ASAP7_75t_R s10235(
.D(net6111),
.CLK(clk),
.QN(net10272)
);

DFFHQNx3_ASAP7_75t_R s10236(
.D(net6280),
.CLK(clk),
.QN(net10273)
);

DFFHQx4_ASAP7_75t_R s10237(
.D(net6320),
.CLK(clk),
.Q(net10274)
);

DFFLQNx1_ASAP7_75t_R s10238(
.D(net6392),
.CLK(clk),
.QN(net10275)
);

DFFLQNx2_ASAP7_75t_R s10239(
.D(net6524),
.CLK(clk),
.QN(net10276)
);

DFFLQNx3_ASAP7_75t_R s10240(
.D(net6530),
.CLK(clk),
.QN(net10277)
);

DFFLQx4_ASAP7_75t_R s10241(
.D(net6544),
.CLK(clk),
.Q(net10278)
);

DHLx1_ASAP7_75t_R s10242(
.D(net6593),
.CLK(clk),
.Q(net10279)
);

DHLx2_ASAP7_75t_R s10243(
.D(net6762),
.CLK(clk),
.Q(net10280)
);

DHLx3_ASAP7_75t_R s10244(
.D(net6793),
.CLK(clk),
.Q(net10281)
);

DLLx1_ASAP7_75t_R s10245(
.D(net6860),
.CLK(clk),
.Q(net10282)
);

DLLx2_ASAP7_75t_R s10246(
.D(net6862),
.CLK(clk),
.Q(net10283)
);

DLLx3_ASAP7_75t_R s10247(
.D(net6992),
.CLK(clk),
.Q(net10284)
);

DFFHQNx1_ASAP7_75t_R s10248(
.D(net7036),
.CLK(clk),
.QN(net10285)
);

DFFHQNx2_ASAP7_75t_R s10249(
.D(net7143),
.CLK(clk),
.QN(net10286)
);

DFFHQNx3_ASAP7_75t_R s10250(
.D(net7144),
.CLK(clk),
.QN(net10287)
);

DFFHQx4_ASAP7_75t_R s10251(
.D(net7204),
.CLK(clk),
.Q(net10288)
);

DFFLQNx1_ASAP7_75t_R s10252(
.D(net7280),
.CLK(clk),
.QN(net10289)
);

DFFLQNx2_ASAP7_75t_R s10253(
.D(net7317),
.CLK(clk),
.QN(net10290)
);

DFFLQNx3_ASAP7_75t_R s10254(
.D(net7330),
.CLK(clk),
.QN(net10291)
);

DFFLQx4_ASAP7_75t_R s10255(
.D(net7366),
.CLK(clk),
.Q(net10292)
);

DHLx1_ASAP7_75t_R s10256(
.D(net7433),
.CLK(clk),
.Q(net10293)
);

DHLx2_ASAP7_75t_R s10257(
.D(net7440),
.CLK(clk),
.Q(net10294)
);

DHLx3_ASAP7_75t_R s10258(
.D(net7447),
.CLK(clk),
.Q(net10295)
);

DLLx1_ASAP7_75t_R s10259(
.D(net7521),
.CLK(clk),
.Q(net10296)
);

DLLx2_ASAP7_75t_R s10260(
.D(net7535),
.CLK(clk),
.Q(net10297)
);

DLLx3_ASAP7_75t_R s10261(
.D(net7612),
.CLK(clk),
.Q(net10298)
);

DFFHQNx1_ASAP7_75t_R s10262(
.D(net7684),
.CLK(clk),
.QN(net10299)
);

DFFHQNx2_ASAP7_75t_R s10263(
.D(net7702),
.CLK(clk),
.QN(net10300)
);

DFFHQNx3_ASAP7_75t_R s10264(
.D(net7779),
.CLK(clk),
.QN(net10301)
);

DFFHQx4_ASAP7_75t_R s10265(
.D(net7819),
.CLK(clk),
.Q(net10302)
);

DFFLQNx1_ASAP7_75t_R s10266(
.D(net7917),
.CLK(clk),
.QN(net10303)
);

DFFLQNx2_ASAP7_75t_R s10267(
.D(net7920),
.CLK(clk),
.QN(net10304)
);

DFFLQNx3_ASAP7_75t_R s10268(
.D(net7931),
.CLK(clk),
.QN(net10305)
);

DFFLQx4_ASAP7_75t_R s10269(
.D(net8023),
.CLK(clk),
.Q(net10306)
);

DHLx1_ASAP7_75t_R s10270(
.D(net8034),
.CLK(clk),
.Q(net10307)
);

DHLx2_ASAP7_75t_R s10271(
.D(net8035),
.CLK(clk),
.Q(net10308)
);

DHLx3_ASAP7_75t_R s10272(
.D(net8089),
.CLK(clk),
.Q(net10309)
);

DLLx1_ASAP7_75t_R s10273(
.D(net8216),
.CLK(clk),
.Q(net10310)
);

DLLx2_ASAP7_75t_R s10274(
.D(net8321),
.CLK(clk),
.Q(net10311)
);

DLLx3_ASAP7_75t_R s10275(
.D(net8335),
.CLK(clk),
.Q(net10312)
);

DFFHQNx1_ASAP7_75t_R s10276(
.D(net8413),
.CLK(clk),
.QN(net10313)
);

DFFHQNx2_ASAP7_75t_R s10277(
.D(net8418),
.CLK(clk),
.QN(net10314)
);

DFFHQNx3_ASAP7_75t_R s10278(
.D(net8462),
.CLK(clk),
.QN(net10315)
);

DFFHQx4_ASAP7_75t_R s10279(
.D(net8464),
.CLK(clk),
.Q(net10316)
);

DFFLQNx1_ASAP7_75t_R s10280(
.D(net8501),
.CLK(clk),
.QN(net10317)
);

DFFLQNx2_ASAP7_75t_R s10281(
.D(net8502),
.CLK(clk),
.QN(net10318)
);

DFFLQNx3_ASAP7_75t_R s10282(
.D(net8657),
.CLK(clk),
.QN(net10319)
);

DFFLQx4_ASAP7_75t_R s10283(
.D(net8698),
.CLK(clk),
.Q(net10320)
);

DHLx1_ASAP7_75t_R s10284(
.D(net8750),
.CLK(clk),
.Q(net10321)
);

DHLx2_ASAP7_75t_R s10285(
.D(net8780),
.CLK(clk),
.Q(net10322)
);

DHLx3_ASAP7_75t_R s10286(
.D(net8802),
.CLK(clk),
.Q(net10323)
);

DLLx1_ASAP7_75t_R s10287(
.D(net8834),
.CLK(clk),
.Q(net10324)
);

DLLx2_ASAP7_75t_R s10288(
.D(net8876),
.CLK(clk),
.Q(net10325)
);

DLLx3_ASAP7_75t_R s10289(
.D(net8921),
.CLK(clk),
.Q(net10326)
);

DFFHQNx1_ASAP7_75t_R s10290(
.D(net8976),
.CLK(clk),
.QN(net10327)
);

DFFHQNx2_ASAP7_75t_R s10291(
.D(net8999),
.CLK(clk),
.QN(net10328)
);

DFFHQNx3_ASAP7_75t_R s10292(
.D(net9085),
.CLK(clk),
.QN(net10329)
);

DFFHQx4_ASAP7_75t_R s10293(
.D(net9093),
.CLK(clk),
.Q(net10330)
);

DFFLQNx1_ASAP7_75t_R s10294(
.D(net9094),
.CLK(clk),
.QN(net10331)
);

DFFLQNx2_ASAP7_75t_R s10295(
.D(net9100),
.CLK(clk),
.QN(net10332)
);

DFFLQNx3_ASAP7_75t_R s10296(
.D(net9106),
.CLK(clk),
.QN(net10333)
);

DFFLQx4_ASAP7_75t_R s10297(
.D(net9108),
.CLK(clk),
.Q(net10334)
);

DHLx1_ASAP7_75t_R s10298(
.D(net9109),
.CLK(clk),
.Q(net10335)
);

DHLx2_ASAP7_75t_R s10299(
.D(net9110),
.CLK(clk),
.Q(net10336)
);

DHLx3_ASAP7_75t_R s10300(
.D(net9112),
.CLK(clk),
.Q(net10337)
);

DLLx1_ASAP7_75t_R s10301(
.D(net9115),
.CLK(clk),
.Q(net10338)
);

DLLx2_ASAP7_75t_R s10302(
.D(net9127),
.CLK(clk),
.Q(net10339)
);

DLLx3_ASAP7_75t_R s10303(
.D(net9128),
.CLK(clk),
.Q(net10340)
);

DFFHQNx1_ASAP7_75t_R s10304(
.D(net9139),
.CLK(clk),
.QN(net10341)
);

DFFHQNx2_ASAP7_75t_R s10305(
.D(net9140),
.CLK(clk),
.QN(net10342)
);

DFFHQNx3_ASAP7_75t_R s10306(
.D(net9161),
.CLK(clk),
.QN(net10343)
);

DFFHQx4_ASAP7_75t_R s10307(
.D(net9163),
.CLK(clk),
.Q(net10344)
);

DFFLQNx1_ASAP7_75t_R s10308(
.D(net9165),
.CLK(clk),
.QN(net10345)
);

DFFLQNx2_ASAP7_75t_R s10309(
.D(net9178),
.CLK(clk),
.QN(net10346)
);

DFFLQNx3_ASAP7_75t_R s10310(
.D(net9179),
.CLK(clk),
.QN(net10347)
);

DFFLQx4_ASAP7_75t_R s10311(
.D(net9192),
.CLK(clk),
.Q(net10348)
);

DHLx1_ASAP7_75t_R s10312(
.D(net9194),
.CLK(clk),
.Q(net10349)
);

DHLx2_ASAP7_75t_R s10313(
.D(net9196),
.CLK(clk),
.Q(net10350)
);

DHLx3_ASAP7_75t_R s10314(
.D(net9205),
.CLK(clk),
.Q(net10351)
);

DLLx1_ASAP7_75t_R s10315(
.D(net9214),
.CLK(clk),
.Q(net10352)
);

DLLx2_ASAP7_75t_R s10316(
.D(net9215),
.CLK(clk),
.Q(net10353)
);

DLLx3_ASAP7_75t_R s10317(
.D(net9222),
.CLK(clk),
.Q(net10354)
);

DFFHQNx1_ASAP7_75t_R s10318(
.D(net9237),
.CLK(clk),
.QN(net10355)
);

DFFHQNx2_ASAP7_75t_R s10319(
.D(net9243),
.CLK(clk),
.QN(net10356)
);

DFFHQNx3_ASAP7_75t_R s10320(
.D(net9245),
.CLK(clk),
.QN(net10357)
);

DFFHQx4_ASAP7_75t_R s10321(
.D(net9249),
.CLK(clk),
.Q(net10358)
);

DFFLQNx1_ASAP7_75t_R s10322(
.D(net9256),
.CLK(clk),
.QN(net10359)
);

DFFLQNx2_ASAP7_75t_R s10323(
.D(net9259),
.CLK(clk),
.QN(net10360)
);

DFFLQNx3_ASAP7_75t_R s10324(
.D(net9263),
.CLK(clk),
.QN(net10361)
);

DFFLQx4_ASAP7_75t_R s10325(
.D(net9266),
.CLK(clk),
.Q(net10362)
);

DHLx1_ASAP7_75t_R s10326(
.D(net9272),
.CLK(clk),
.Q(net10363)
);

DHLx2_ASAP7_75t_R s10327(
.D(net9274),
.CLK(clk),
.Q(net10364)
);

DHLx3_ASAP7_75t_R s10328(
.D(net9276),
.CLK(clk),
.Q(net10365)
);

DLLx1_ASAP7_75t_R s10329(
.D(net9277),
.CLK(clk),
.Q(net10366)
);

DLLx2_ASAP7_75t_R s10330(
.D(net9278),
.CLK(clk),
.Q(net10367)
);

DLLx3_ASAP7_75t_R s10331(
.D(net9284),
.CLK(clk),
.Q(net10368)
);

DFFHQNx1_ASAP7_75t_R s10332(
.D(net9287),
.CLK(clk),
.QN(net10369)
);

DFFHQNx2_ASAP7_75t_R s10333(
.D(net9290),
.CLK(clk),
.QN(net10370)
);

DFFHQNx3_ASAP7_75t_R s10334(
.D(net9292),
.CLK(clk),
.QN(net10371)
);

DFFHQx4_ASAP7_75t_R s10335(
.D(net9294),
.CLK(clk),
.Q(net10372)
);

DFFLQNx1_ASAP7_75t_R s10336(
.D(net9295),
.CLK(clk),
.QN(net10373)
);

DFFLQNx2_ASAP7_75t_R s10337(
.D(net9299),
.CLK(clk),
.QN(net10374)
);

DFFLQNx3_ASAP7_75t_R s10338(
.D(net9300),
.CLK(clk),
.QN(net10375)
);

DFFLQx4_ASAP7_75t_R s10339(
.D(net9301),
.CLK(clk),
.Q(net10376)
);

DHLx1_ASAP7_75t_R s10340(
.D(net9302),
.CLK(clk),
.Q(net10377)
);

DHLx2_ASAP7_75t_R s10341(
.D(net9303),
.CLK(clk),
.Q(net10378)
);

DHLx3_ASAP7_75t_R s10342(
.D(net9304),
.CLK(clk),
.Q(net10379)
);

DLLx1_ASAP7_75t_R s10343(
.D(net9305),
.CLK(clk),
.Q(net10380)
);

DLLx2_ASAP7_75t_R s10344(
.D(net9306),
.CLK(clk),
.Q(net10381)
);

DLLx3_ASAP7_75t_R s10345(
.D(net9307),
.CLK(clk),
.Q(net10382)
);

DFFHQNx1_ASAP7_75t_R s10346(
.D(net9308),
.CLK(clk),
.QN(net10383)
);

DFFHQNx2_ASAP7_75t_R s10347(
.D(net9309),
.CLK(clk),
.QN(net10384)
);

DFFHQNx3_ASAP7_75t_R s10348(
.D(net9314),
.CLK(clk),
.QN(net10385)
);

DFFHQx4_ASAP7_75t_R s10349(
.D(net9320),
.CLK(clk),
.Q(net10386)
);

DFFLQNx1_ASAP7_75t_R s10350(
.D(net9322),
.CLK(clk),
.QN(net10387)
);

DFFLQNx2_ASAP7_75t_R s10351(
.D(net9328),
.CLK(clk),
.QN(net10388)
);

DFFLQNx3_ASAP7_75t_R s10352(
.D(net9331),
.CLK(clk),
.QN(net10389)
);

DFFLQx4_ASAP7_75t_R s10353(
.D(net9333),
.CLK(clk),
.Q(net10390)
);

DHLx1_ASAP7_75t_R s10354(
.D(net9335),
.CLK(clk),
.Q(net10391)
);

DHLx2_ASAP7_75t_R s10355(
.D(net9336),
.CLK(clk),
.Q(net10392)
);

DHLx3_ASAP7_75t_R s10356(
.D(net9338),
.CLK(clk),
.Q(net10393)
);

DLLx1_ASAP7_75t_R s10357(
.D(net9339),
.CLK(clk),
.Q(net10394)
);

DLLx2_ASAP7_75t_R s10358(
.D(net9340),
.CLK(clk),
.Q(net10395)
);

DLLx3_ASAP7_75t_R s10359(
.D(net9341),
.CLK(clk),
.Q(net10396)
);

DFFHQNx1_ASAP7_75t_R s10360(
.D(net9342),
.CLK(clk),
.QN(net10397)
);

DFFHQNx2_ASAP7_75t_R s10361(
.D(net9345),
.CLK(clk),
.QN(net10398)
);

DFFHQNx3_ASAP7_75t_R s10362(
.D(net9346),
.CLK(clk),
.QN(net10399)
);

DFFHQx4_ASAP7_75t_R s10363(
.D(net9347),
.CLK(clk),
.Q(net10400)
);

DFFLQNx1_ASAP7_75t_R s10364(
.D(net9348),
.CLK(clk),
.QN(net10401)
);

DFFLQNx2_ASAP7_75t_R s10365(
.D(net9349),
.CLK(clk),
.QN(net10402)
);

DFFLQNx3_ASAP7_75t_R s10366(
.D(net9350),
.CLK(clk),
.QN(net10403)
);

DFFLQx4_ASAP7_75t_R s10367(
.D(net9352),
.CLK(clk),
.Q(net10404)
);

DHLx1_ASAP7_75t_R s10368(
.D(net9355),
.CLK(clk),
.Q(net10405)
);

DHLx2_ASAP7_75t_R s10369(
.D(net9356),
.CLK(clk),
.Q(net10406)
);

DHLx3_ASAP7_75t_R s10370(
.D(net9357),
.CLK(clk),
.Q(net10407)
);

DLLx1_ASAP7_75t_R s10371(
.D(net9358),
.CLK(clk),
.Q(net10408)
);

DLLx2_ASAP7_75t_R s10372(
.D(net9359),
.CLK(clk),
.Q(net10409)
);

DLLx3_ASAP7_75t_R s10373(
.D(net9363),
.CLK(clk),
.Q(net10410)
);

DFFHQNx1_ASAP7_75t_R s10374(
.D(net9364),
.CLK(clk),
.QN(net10411)
);

DFFHQNx2_ASAP7_75t_R s10375(
.D(net9368),
.CLK(clk),
.QN(net10412)
);

DFFHQNx3_ASAP7_75t_R s10376(
.D(net9369),
.CLK(clk),
.QN(net10413)
);

DFFHQx4_ASAP7_75t_R s10377(
.D(net9371),
.CLK(clk),
.Q(net10414)
);

DFFLQNx1_ASAP7_75t_R s10378(
.D(net9375),
.CLK(clk),
.QN(net10415)
);

DFFLQNx2_ASAP7_75t_R s10379(
.D(net9377),
.CLK(clk),
.QN(net10416)
);

DFFLQNx3_ASAP7_75t_R s10380(
.D(net9378),
.CLK(clk),
.QN(net10417)
);

DFFLQx4_ASAP7_75t_R s10381(
.D(net9379),
.CLK(clk),
.Q(net10418)
);

DHLx1_ASAP7_75t_R s10382(
.D(net9381),
.CLK(clk),
.Q(net10419)
);

DHLx2_ASAP7_75t_R s10383(
.D(net9382),
.CLK(clk),
.Q(net10420)
);

DHLx3_ASAP7_75t_R s10384(
.D(net9383),
.CLK(clk),
.Q(net10421)
);

DLLx1_ASAP7_75t_R s10385(
.D(net9384),
.CLK(clk),
.Q(net10422)
);

DLLx2_ASAP7_75t_R s10386(
.D(net9386),
.CLK(clk),
.Q(net10423)
);

DLLx3_ASAP7_75t_R s10387(
.D(net9387),
.CLK(clk),
.Q(net10424)
);

DFFHQNx1_ASAP7_75t_R s10388(
.D(net9389),
.CLK(clk),
.QN(net10425)
);

DFFHQNx2_ASAP7_75t_R s10389(
.D(net9390),
.CLK(clk),
.QN(net10426)
);

DFFHQNx3_ASAP7_75t_R s10390(
.D(net9391),
.CLK(clk),
.QN(net10427)
);

DFFHQx4_ASAP7_75t_R s10391(
.D(net9393),
.CLK(clk),
.Q(net10428)
);

DFFLQNx1_ASAP7_75t_R s10392(
.D(net9395),
.CLK(clk),
.QN(net10429)
);

DFFLQNx2_ASAP7_75t_R s10393(
.D(net9396),
.CLK(clk),
.QN(net10430)
);

DFFLQNx3_ASAP7_75t_R s10394(
.D(net9398),
.CLK(clk),
.QN(net10431)
);

DFFLQx4_ASAP7_75t_R s10395(
.D(net9399),
.CLK(clk),
.Q(net10432)
);

DHLx1_ASAP7_75t_R s10396(
.D(net9400),
.CLK(clk),
.Q(net10433)
);

DHLx2_ASAP7_75t_R s10397(
.D(net9401),
.CLK(clk),
.Q(net10434)
);

DHLx3_ASAP7_75t_R s10398(
.D(net9402),
.CLK(clk),
.Q(net10435)
);

DLLx1_ASAP7_75t_R s10399(
.D(net9404),
.CLK(clk),
.Q(net10436)
);

DLLx2_ASAP7_75t_R s10400(
.D(net9406),
.CLK(clk),
.Q(net10437)
);

DLLx3_ASAP7_75t_R s10401(
.D(net9409),
.CLK(clk),
.Q(net10438)
);

DFFHQNx1_ASAP7_75t_R s10402(
.D(net9411),
.CLK(clk),
.QN(net10439)
);

DFFHQNx2_ASAP7_75t_R s10403(
.D(net9412),
.CLK(clk),
.QN(net10440)
);

DFFHQNx3_ASAP7_75t_R s10404(
.D(net9413),
.CLK(clk),
.QN(net10441)
);

DFFHQx4_ASAP7_75t_R s10405(
.D(net9414),
.CLK(clk),
.Q(net10442)
);

DFFLQNx1_ASAP7_75t_R s10406(
.D(net9416),
.CLK(clk),
.QN(net10443)
);

DFFLQNx2_ASAP7_75t_R s10407(
.D(net9417),
.CLK(clk),
.QN(net10444)
);

DFFLQNx3_ASAP7_75t_R s10408(
.D(net9418),
.CLK(clk),
.QN(net10445)
);

DFFLQx4_ASAP7_75t_R s10409(
.D(net9419),
.CLK(clk),
.Q(net10446)
);

DHLx1_ASAP7_75t_R s10410(
.D(net9420),
.CLK(clk),
.Q(net10447)
);

DHLx2_ASAP7_75t_R s10411(
.D(net9422),
.CLK(clk),
.Q(net10448)
);

DHLx3_ASAP7_75t_R s10412(
.D(net9424),
.CLK(clk),
.Q(net10449)
);

DLLx1_ASAP7_75t_R s10413(
.D(net9425),
.CLK(clk),
.Q(net10450)
);

DLLx2_ASAP7_75t_R s10414(
.D(net9427),
.CLK(clk),
.Q(net10451)
);

DLLx3_ASAP7_75t_R s10415(
.D(net9428),
.CLK(clk),
.Q(net10452)
);

DFFHQNx1_ASAP7_75t_R s10416(
.D(net9429),
.CLK(clk),
.QN(net10453)
);

DFFHQNx2_ASAP7_75t_R s10417(
.D(net9430),
.CLK(clk),
.QN(net10454)
);

DFFHQNx3_ASAP7_75t_R s10418(
.D(net9431),
.CLK(clk),
.QN(net10455)
);

DFFHQx4_ASAP7_75t_R s10419(
.D(net9434),
.CLK(clk),
.Q(net10456)
);

DFFLQNx1_ASAP7_75t_R s10420(
.D(net9435),
.CLK(clk),
.QN(net10457)
);

DFFLQNx2_ASAP7_75t_R s10421(
.D(net9436),
.CLK(clk),
.QN(net10458)
);

DFFLQNx3_ASAP7_75t_R s10422(
.D(net9439),
.CLK(clk),
.QN(net10459)
);

DFFLQx4_ASAP7_75t_R s10423(
.D(net9440),
.CLK(clk),
.Q(net10460)
);

DHLx1_ASAP7_75t_R s10424(
.D(net9441),
.CLK(clk),
.Q(net10461)
);

DHLx2_ASAP7_75t_R s10425(
.D(net9445),
.CLK(clk),
.Q(net10462)
);

DHLx3_ASAP7_75t_R s10426(
.D(net9447),
.CLK(clk),
.Q(net10463)
);

DLLx1_ASAP7_75t_R s10427(
.D(net9449),
.CLK(clk),
.Q(net10464)
);

DLLx2_ASAP7_75t_R s10428(
.D(net9450),
.CLK(clk),
.Q(net10465)
);

DLLx3_ASAP7_75t_R s10429(
.D(net9453),
.CLK(clk),
.Q(net10466)
);

DFFHQNx1_ASAP7_75t_R s10430(
.D(net9454),
.CLK(clk),
.QN(net10467)
);

DFFHQNx2_ASAP7_75t_R s10431(
.D(net9455),
.CLK(clk),
.QN(net10468)
);

DFFHQNx3_ASAP7_75t_R s10432(
.D(net9463),
.CLK(clk),
.QN(net10469)
);

DFFHQx4_ASAP7_75t_R s10433(
.D(net9464),
.CLK(clk),
.Q(net10470)
);

DFFLQNx1_ASAP7_75t_R s10434(
.D(net9465),
.CLK(clk),
.QN(net10471)
);

DFFLQNx2_ASAP7_75t_R s10435(
.D(net9472),
.CLK(clk),
.QN(net10472)
);

DFFLQNx3_ASAP7_75t_R s10436(
.D(net9474),
.CLK(clk),
.QN(net10473)
);

DFFLQx4_ASAP7_75t_R s10437(
.D(net9475),
.CLK(clk),
.Q(net10474)
);

DHLx1_ASAP7_75t_R s10438(
.D(net9476),
.CLK(clk),
.Q(net10475)
);

DHLx2_ASAP7_75t_R s10439(
.D(net9477),
.CLK(clk),
.Q(net10476)
);

DHLx3_ASAP7_75t_R s10440(
.D(net9478),
.CLK(clk),
.Q(net10477)
);

DLLx1_ASAP7_75t_R s10441(
.D(net9480),
.CLK(clk),
.Q(net10478)
);

DLLx2_ASAP7_75t_R s10442(
.D(net9482),
.CLK(clk),
.Q(net10479)
);

DLLx3_ASAP7_75t_R s10443(
.D(net9483),
.CLK(clk),
.Q(net10480)
);

DFFHQNx1_ASAP7_75t_R s10444(
.D(net9484),
.CLK(clk),
.QN(net10481)
);

DFFHQNx2_ASAP7_75t_R s10445(
.D(net9487),
.CLK(clk),
.QN(net10482)
);

DFFHQNx3_ASAP7_75t_R s10446(
.D(net9488),
.CLK(clk),
.QN(net10483)
);

DFFHQx4_ASAP7_75t_R s10447(
.D(net9490),
.CLK(clk),
.Q(net10484)
);

DFFLQNx1_ASAP7_75t_R s10448(
.D(net9491),
.CLK(clk),
.QN(net10485)
);

DFFLQNx2_ASAP7_75t_R s10449(
.D(net9493),
.CLK(clk),
.QN(net10486)
);

DFFLQNx3_ASAP7_75t_R s10450(
.D(net9494),
.CLK(clk),
.QN(net10487)
);

DFFLQx4_ASAP7_75t_R s10451(
.D(net9495),
.CLK(clk),
.Q(net10488)
);

DHLx1_ASAP7_75t_R s10452(
.D(net9496),
.CLK(clk),
.Q(net10489)
);

DHLx2_ASAP7_75t_R s10453(
.D(net9497),
.CLK(clk),
.Q(net10490)
);

DHLx3_ASAP7_75t_R s10454(
.D(net9499),
.CLK(clk),
.Q(net10491)
);

DLLx1_ASAP7_75t_R s10455(
.D(net9500),
.CLK(clk),
.Q(net10492)
);

DLLx2_ASAP7_75t_R s10456(
.D(net9501),
.CLK(clk),
.Q(net10493)
);

DLLx3_ASAP7_75t_R s10457(
.D(net9504),
.CLK(clk),
.Q(net10494)
);

DFFHQNx1_ASAP7_75t_R s10458(
.D(net9507),
.CLK(clk),
.QN(net10495)
);

DFFHQNx2_ASAP7_75t_R s10459(
.D(net9508),
.CLK(clk),
.QN(net10496)
);

DFFHQNx3_ASAP7_75t_R s10460(
.D(net9509),
.CLK(clk),
.QN(net10497)
);

DFFHQx4_ASAP7_75t_R s10461(
.D(net9510),
.CLK(clk),
.Q(net10498)
);

DFFLQNx1_ASAP7_75t_R s10462(
.D(net9512),
.CLK(clk),
.QN(net10499)
);

DFFLQNx2_ASAP7_75t_R s10463(
.D(net9513),
.CLK(clk),
.QN(net10500)
);

DFFLQNx3_ASAP7_75t_R s10464(
.D(net9514),
.CLK(clk),
.QN(net10501)
);

DFFLQx4_ASAP7_75t_R s10465(
.D(net9516),
.CLK(clk),
.Q(net10502)
);

DHLx1_ASAP7_75t_R s10466(
.D(net9517),
.CLK(clk),
.Q(net10503)
);

DHLx2_ASAP7_75t_R s10467(
.D(net9519),
.CLK(clk),
.Q(net10504)
);

DHLx3_ASAP7_75t_R s10468(
.D(net9520),
.CLK(clk),
.Q(net10505)
);

DLLx1_ASAP7_75t_R s10469(
.D(net9523),
.CLK(clk),
.Q(net10506)
);

DLLx2_ASAP7_75t_R s10470(
.D(net9524),
.CLK(clk),
.Q(net10507)
);

DLLx3_ASAP7_75t_R s10471(
.D(net9526),
.CLK(clk),
.Q(net10508)
);

DFFHQNx1_ASAP7_75t_R s10472(
.D(net9527),
.CLK(clk),
.QN(net10509)
);

DFFHQNx2_ASAP7_75t_R s10473(
.D(net9528),
.CLK(clk),
.QN(net10510)
);

DFFHQNx3_ASAP7_75t_R s10474(
.D(net9531),
.CLK(clk),
.QN(net10511)
);

DFFHQx4_ASAP7_75t_R s10475(
.D(net9533),
.CLK(clk),
.Q(net10512)
);

DFFLQNx1_ASAP7_75t_R s10476(
.D(net9536),
.CLK(clk),
.QN(net10513)
);

DFFLQNx2_ASAP7_75t_R s10477(
.D(net9537),
.CLK(clk),
.QN(net10514)
);

DFFLQNx3_ASAP7_75t_R s10478(
.D(net9539),
.CLK(clk),
.QN(net10515)
);

DFFLQx4_ASAP7_75t_R s10479(
.D(net9543),
.CLK(clk),
.Q(net10516)
);

DHLx1_ASAP7_75t_R s10480(
.D(net9546),
.CLK(clk),
.Q(net10517)
);

DHLx2_ASAP7_75t_R s10481(
.D(net9547),
.CLK(clk),
.Q(net10518)
);

DHLx3_ASAP7_75t_R s10482(
.D(net9548),
.CLK(clk),
.Q(net10519)
);

DLLx1_ASAP7_75t_R s10483(
.D(net9550),
.CLK(clk),
.Q(net10520)
);

DLLx2_ASAP7_75t_R s10484(
.D(net9552),
.CLK(clk),
.Q(net10521)
);

DLLx3_ASAP7_75t_R s10485(
.D(net9553),
.CLK(clk),
.Q(net10522)
);

DFFHQNx1_ASAP7_75t_R s10486(
.D(net9554),
.CLK(clk),
.QN(net10523)
);

DFFHQNx2_ASAP7_75t_R s10487(
.D(net9555),
.CLK(clk),
.QN(net10524)
);

DFFHQNx3_ASAP7_75t_R s10488(
.D(net9557),
.CLK(clk),
.QN(net10525)
);

DFFHQx4_ASAP7_75t_R s10489(
.D(net9559),
.CLK(clk),
.Q(net10526)
);

DFFLQNx1_ASAP7_75t_R s10490(
.D(net9560),
.CLK(clk),
.QN(net10527)
);

DFFLQNx2_ASAP7_75t_R s10491(
.D(net9561),
.CLK(clk),
.QN(net10528)
);

DFFLQNx3_ASAP7_75t_R s10492(
.D(net9562),
.CLK(clk),
.QN(net10529)
);

DFFLQx4_ASAP7_75t_R s10493(
.D(net9563),
.CLK(clk),
.Q(net10530)
);

DHLx1_ASAP7_75t_R s10494(
.D(net9564),
.CLK(clk),
.Q(net10531)
);

DHLx2_ASAP7_75t_R s10495(
.D(net9565),
.CLK(clk),
.Q(net10532)
);

DHLx3_ASAP7_75t_R s10496(
.D(net9566),
.CLK(clk),
.Q(net10533)
);

DLLx1_ASAP7_75t_R s10497(
.D(net9567),
.CLK(clk),
.Q(net10534)
);

DLLx2_ASAP7_75t_R s10498(
.D(net9568),
.CLK(clk),
.Q(net10535)
);

DLLx3_ASAP7_75t_R s10499(
.D(net9569),
.CLK(clk),
.Q(net10536)
);

DFFHQNx1_ASAP7_75t_R s10500(
.D(net9572),
.CLK(clk),
.QN(net10537)
);

DFFHQNx2_ASAP7_75t_R s10501(
.D(net9573),
.CLK(clk),
.QN(net10538)
);

DFFHQNx3_ASAP7_75t_R s10502(
.D(net9575),
.CLK(clk),
.QN(net10539)
);

DFFHQx4_ASAP7_75t_R s10503(
.D(net9576),
.CLK(clk),
.Q(net10540)
);

DFFLQNx1_ASAP7_75t_R s10504(
.D(net9578),
.CLK(clk),
.QN(net10541)
);

DFFLQNx2_ASAP7_75t_R s10505(
.D(net9579),
.CLK(clk),
.QN(net10542)
);

DFFLQNx3_ASAP7_75t_R s10506(
.D(net9580),
.CLK(clk),
.QN(net10543)
);

DFFLQx4_ASAP7_75t_R s10507(
.D(net9582),
.CLK(clk),
.Q(net10544)
);

DHLx1_ASAP7_75t_R s10508(
.D(net9583),
.CLK(clk),
.Q(net10545)
);

DHLx2_ASAP7_75t_R s10509(
.D(net9585),
.CLK(clk),
.Q(net10546)
);

DHLx3_ASAP7_75t_R s10510(
.D(net9586),
.CLK(clk),
.Q(net10547)
);

DLLx1_ASAP7_75t_R s10511(
.D(net9587),
.CLK(clk),
.Q(net10548)
);

DLLx2_ASAP7_75t_R s10512(
.D(net9588),
.CLK(clk),
.Q(net10549)
);

DLLx3_ASAP7_75t_R s10513(
.D(net9590),
.CLK(clk),
.Q(net10550)
);

DFFHQNx1_ASAP7_75t_R s10514(
.D(net9592),
.CLK(clk),
.QN(net10551)
);

DFFHQNx2_ASAP7_75t_R s10515(
.D(net9593),
.CLK(clk),
.QN(net10552)
);

DFFHQNx3_ASAP7_75t_R s10516(
.D(net9595),
.CLK(clk),
.QN(net10553)
);

DFFHQx4_ASAP7_75t_R s10517(
.D(net9596),
.CLK(clk),
.Q(net10554)
);

DFFLQNx1_ASAP7_75t_R s10518(
.D(net9597),
.CLK(clk),
.QN(net10555)
);

DFFLQNx2_ASAP7_75t_R s10519(
.D(net9600),
.CLK(clk),
.QN(net10556)
);

DFFLQNx3_ASAP7_75t_R s10520(
.D(net9603),
.CLK(clk),
.QN(net10557)
);

DFFLQx4_ASAP7_75t_R s10521(
.D(net9604),
.CLK(clk),
.Q(net10558)
);

DHLx1_ASAP7_75t_R s10522(
.D(net9607),
.CLK(clk),
.Q(net10559)
);

DHLx2_ASAP7_75t_R s10523(
.D(net9608),
.CLK(clk),
.Q(net10560)
);

DHLx3_ASAP7_75t_R s10524(
.D(net9609),
.CLK(clk),
.Q(net10561)
);

DLLx1_ASAP7_75t_R s10525(
.D(net9611),
.CLK(clk),
.Q(net10562)
);

DLLx2_ASAP7_75t_R s10526(
.D(net9612),
.CLK(clk),
.Q(net10563)
);

DLLx3_ASAP7_75t_R s10527(
.D(net9613),
.CLK(clk),
.Q(net10564)
);

DFFHQNx1_ASAP7_75t_R s10528(
.D(net9614),
.CLK(clk),
.QN(net10565)
);

DFFHQNx2_ASAP7_75t_R s10529(
.D(net9615),
.CLK(clk),
.QN(net10566)
);

DFFHQNx3_ASAP7_75t_R s10530(
.D(net9618),
.CLK(clk),
.QN(net10567)
);

DFFHQx4_ASAP7_75t_R s10531(
.D(net9620),
.CLK(clk),
.Q(net10568)
);

DFFLQNx1_ASAP7_75t_R s10532(
.D(net9623),
.CLK(clk),
.QN(net10569)
);

DFFLQNx2_ASAP7_75t_R s10533(
.D(net9624),
.CLK(clk),
.QN(net10570)
);

DFFLQNx3_ASAP7_75t_R s10534(
.D(net9625),
.CLK(clk),
.QN(net10571)
);

DFFLQx4_ASAP7_75t_R s10535(
.D(net9627),
.CLK(clk),
.Q(net10572)
);

DHLx1_ASAP7_75t_R s10536(
.D(net9629),
.CLK(clk),
.Q(net10573)
);

DHLx2_ASAP7_75t_R s10537(
.D(net9630),
.CLK(clk),
.Q(net10574)
);

DHLx3_ASAP7_75t_R s10538(
.D(net9631),
.CLK(clk),
.Q(net10575)
);

DLLx1_ASAP7_75t_R s10539(
.D(net9632),
.CLK(clk),
.Q(net10576)
);


endmodule
